* NGSPICE file created from tinyrv.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

.subckt tinyrv clk inst[0] inst[10] inst[11] inst[12] inst[13] inst[14] inst[15] inst[16]
+ inst[17] inst[18] inst[19] inst[1] inst[20] inst[21] inst[22] inst[23] inst[24]
+ inst[25] inst[26] inst[27] inst[28] inst[29] inst[2] inst[30] inst[31] inst[3] inst[4]
+ inst[5] inst[6] inst[7] inst[8] inst[9] mem_addr[0] mem_addr[10] mem_addr[11] mem_addr[12]
+ mem_addr[13] mem_addr[14] mem_addr[15] mem_addr[16] mem_addr[17] mem_addr[18] mem_addr[19]
+ mem_addr[1] mem_addr[20] mem_addr[21] mem_addr[22] mem_addr[23] mem_addr[24] mem_addr[25]
+ mem_addr[26] mem_addr[27] mem_addr[28] mem_addr[29] mem_addr[2] mem_addr[30] mem_addr[31]
+ mem_addr[3] mem_addr[4] mem_addr[5] mem_addr[6] mem_addr[7] mem_addr[8] mem_addr[9]
+ mem_ld_dat[0] mem_ld_dat[10] mem_ld_dat[11] mem_ld_dat[12] mem_ld_dat[13] mem_ld_dat[14]
+ mem_ld_dat[15] mem_ld_dat[16] mem_ld_dat[17] mem_ld_dat[18] mem_ld_dat[19] mem_ld_dat[1]
+ mem_ld_dat[20] mem_ld_dat[21] mem_ld_dat[22] mem_ld_dat[23] mem_ld_dat[24] mem_ld_dat[25]
+ mem_ld_dat[26] mem_ld_dat[27] mem_ld_dat[28] mem_ld_dat[29] mem_ld_dat[2] mem_ld_dat[30]
+ mem_ld_dat[31] mem_ld_dat[3] mem_ld_dat[4] mem_ld_dat[5] mem_ld_dat[6] mem_ld_dat[7]
+ mem_ld_dat[8] mem_ld_dat[9] mem_ld_en mem_ld_mask[0] mem_ld_mask[1] mem_ld_mask[2]
+ mem_ld_mask[3] mem_st_dat[0] mem_st_dat[10] mem_st_dat[11] mem_st_dat[12] mem_st_dat[13]
+ mem_st_dat[14] mem_st_dat[15] mem_st_dat[16] mem_st_dat[17] mem_st_dat[18] mem_st_dat[19]
+ mem_st_dat[1] mem_st_dat[20] mem_st_dat[21] mem_st_dat[22] mem_st_dat[23] mem_st_dat[24]
+ mem_st_dat[25] mem_st_dat[26] mem_st_dat[27] mem_st_dat[28] mem_st_dat[29] mem_st_dat[2]
+ mem_st_dat[30] mem_st_dat[31] mem_st_dat[3] mem_st_dat[4] mem_st_dat[5] mem_st_dat[6]
+ mem_st_dat[7] mem_st_dat[8] mem_st_dat[9] mem_st_en mem_st_mask[0] mem_st_mask[1]
+ mem_st_mask[2] mem_st_mask[3] pc[0] pc[10] pc[11] pc[12] pc[13] pc[14] pc[15] pc[16]
+ pc[17] pc[18] pc[19] pc[1] pc[20] pc[21] pc[22] pc[23] pc[24] pc[25] pc[26] pc[27]
+ pc[28] pc[29] pc[2] pc[30] pc[31] pc[3] pc[4] pc[5] pc[6] pc[7] pc[8] pc[9] pc_next[0]
+ pc_next[10] pc_next[11] pc_next[12] pc_next[13] pc_next[14] pc_next[15] pc_next[16]
+ pc_next[17] pc_next[18] pc_next[19] pc_next[1] pc_next[20] pc_next[21] pc_next[22]
+ pc_next[23] pc_next[24] pc_next[25] pc_next[26] pc_next[27] pc_next[28] pc_next[29]
+ pc_next[2] pc_next[30] pc_next[31] pc_next[3] pc_next[4] pc_next[5] pc_next[6] pc_next[7]
+ pc_next[8] pc_next[9] vdd vss
XANTENNA__5760__S0 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9002__S _4421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7963_ reg_file.reg_storage\[5\]\[31\] _3399_ _3752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6914_ _2798_ _2768_ _2805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8841__S _4315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7894_ _2967_ _3534_ _3036_ net48 _3691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6845_ _2583_ _2733_ _2738_ _2739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9633_ _0419_ clknet_leaf_126_clk reg_file.reg_storage\[4\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9564_ _0350_ clknet_leaf_102_clk reg_file.reg_storage\[10\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8640__I _3509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6776_ _2564_ _2672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8515_ reg_file.reg_storage\[13\]\[29\] _4109_ _4114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5727_ reg_file.reg_storage\[4\]\[19\] reg_file.reg_storage\[5\]\[19\] reg_file.reg_storage\[6\]\[19\]
+ reg_file.reg_storage\[7\]\[19\] _1590_ _1642_ _1643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_9495_ _0281_ clknet_leaf_108_clk reg_file.reg_storage\[8\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8446_ _4072_ _4073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6160__I _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ reg_file.reg_storage\[4\]\[22\] reg_file.reg_storage\[5\]\[22\] reg_file.reg_storage\[6\]\[22\]
+ reg_file.reg_storage\[7\]\[22\] _1463_ _1569_ _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_input73_I pc[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5589_ _1499_ _1502_ _1503_ _1504_ _1455_ _1395_ _1505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_115_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7893__A1 _3660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4609_ _0510_ _0527_ _0532_ _0487_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_8377_ _3933_ _4025_ _4032_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7328_ _3165_ _1692_ _3168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_13_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7259_ _3087_ _3090_ _3105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5504__I _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6335__I _2183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4631__A1 _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6070__I _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer7 net209 net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7636__B2 _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7636__A1 _2085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5742__S0 _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5111__A2 _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7939__A2 _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8661__S _4186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4960_ _0874_ _0875_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4891_ _0806_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6630_ _2531_ net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_58_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6561_ _2248_ _2178_ _2464_ _2465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_61_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5512_ _1359_ _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8300_ _3666_ _3973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8116__A2 _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6492_ _2157_ _2398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9280_ _0066_ clknet_leaf_132_clk reg_file.reg_storage\[2\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5443_ _1358_ _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8231_ _3921_ _3922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_76_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8162_ _3867_ _3879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5374_ _1289_ _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7113_ _1828_ _2989_ _2991_ net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7627__A1 _3428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8093_ reg_file.reg_storage\[2\]\[13\] _3598_ _3821_ _3836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5324__I _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7044_ _2926_ _2929_ _2930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6850__A2 _2439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4861__A1 _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8995_ reg_file.reg_storage\[1\]\[8\] _3530_ _4421_ _4423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6602__A2 _2224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7946_ _3360_ _3505_ _3737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7877_ _3660_ _3675_ _3676_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9616_ _0402_ clknet_leaf_70_clk reg_file.reg_storage\[1\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6828_ _1853_ _2721_ _2722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_77_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8355__A2 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4916__A2 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6759_ _1910_ _1909_ _2656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9547_ _0333_ clknet_leaf_1_clk reg_file.reg_storage\[10\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9478_ _0264_ clknet_leaf_32_clk reg_file.reg_storage\[8\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8429_ reg_file.reg_storage\[14\]\[27\] _4059_ _4062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5341__A2 _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7618__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6841__A2 _2304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5652__I0 _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6357__A1 _1938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__I _3442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5883__A3 _1797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5090_ reg_file.reg_storage\[8\]\[29\] reg_file.reg_storage\[9\]\[29\] reg_file.reg_storage\[10\]\[29\]
+ reg_file.reg_storage\[11\]\[29\] _0999_ _0903_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_71_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4983__I _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8034__A1 _3705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8585__A2 _4154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7800_ _3515_ _3605_ _3539_ _3606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8780_ reg_file.reg_storage\[11\]\[21\] _4286_ _4291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6596__A1 _2494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5399__A2 _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5992_ _0720_ _0726_ _0732_ _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__4932__B _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7731_ net128 _3432_ _3540_ _3541_ _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_4943_ reg_file.reg_storage\[1\]\[23\] _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_129_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8190__I _3873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7662_ _3477_ _3478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9401_ _0187_ clknet_leaf_96_clk reg_file.reg_storage\[14\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6613_ _1815_ _2487_ _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4874_ _0754_ _0789_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7545__B1 _3366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7593_ net33 net63 _3412_ _3413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_9332_ _0118_ clknet_leaf_24_clk reg_file.reg_storage\[6\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6544_ _1194_ _2446_ _2448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_6_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7848__A1 _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9263_ _0049_ clknet_leaf_58_clk reg_file.reg_storage\[3\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6475_ _1216_ _2363_ _1205_ _2381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_15_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8214_ _3740_ _3905_ _3908_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5426_ _1234_ _1341_ _0744_ _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9194_ reg_file.reg_storage\[15\]\[23\] _4511_ _4543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_7_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8145_ _3867_ _3868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5357_ reg_file.reg_storage\[2\]\[5\] reg_file.reg_storage\[3\]\[5\] _0637_ _1273_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5288_ _0890_ _1203_ _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8076_ _3826_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input36_I mem_ld_dat[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5087__A1 _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8365__I _4023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7027_ _2906_ _2912_ _2081_ _2913_ _2914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4893__I _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8576__A2 _4147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8978_ reg_file.reg_storage\[1\]\[1\] _4412_ _4413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7929_ _3399_ _3722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8328__A2 _3915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4988__I2 reg_file.reg_storage\[14\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5011__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8500__A2 _4101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7444__I net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8476__S _4078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6814__A2 _2707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5078__A1 _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8016__A1 _3638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__S1 _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4825__B2 _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8567__A2 _4147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8319__A2 _3922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4590_ reg_file.reg_storage\[8\]\[1\] reg_file.reg_storage\[9\]\[1\] reg_file.reg_storage\[10\]\[1\]
+ reg_file.reg_storage\[11\]\[1\] _0513_ _0514_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_142_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7354__I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6260_ _1768_ _2171_ _2172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5211_ reg_file.reg_storage\[12\]\[12\] reg_file.reg_storage\[13\]\[12\] reg_file.reg_storage\[14\]\[12\]
+ reg_file.reg_storage\[15\]\[12\] _0767_ _1047_ _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6191_ _1977_ _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ _0794_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5164__S1 _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_84_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5073_ _0954_ _0986_ _0987_ _0988_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8901_ reg_file.reg_storage\[9\]\[2\] _4185_ _4366_ _4367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8832_ reg_file.reg_storage\[10\]\[8\] _4200_ _4322_ _4324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_99_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8763_ _4261_ _4281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ net204 _0997_ _1890_ _1891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7714_ _3515_ _3523_ _3525_ _3526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4926_ _0635_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5792__A2 _1707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8694_ reg_file.reg_storage\[8\]\[23\] _4181_ _4235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7645_ net58 net35 net43 net52 _3407_ _3461_ _3462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_117_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4857_ _0772_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5049__I _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_22_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7576_ _3390_ _3395_ _3396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_62_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4888__I _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6527_ _1825_ _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9315_ _0101_ clknet_leaf_0_clk reg_file.reg_storage\[6\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4788_ _0703_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9246_ _0032_ clknet_leaf_116_clk reg_file.reg_storage\[3\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6458_ _2018_ _2298_ _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9177_ _4533_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5409_ reg_file.reg_storage\[4\]\[1\] reg_file.reg_storage\[5\]\[1\] reg_file.reg_storage\[6\]\[1\]
+ reg_file.reg_storage\[7\]\[1\] _0632_ _0641_ _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6389_ _1939_ _1940_ _2298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8128_ reg_file.reg_storage\[2\]\[28\] _3852_ _3856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output142_I net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8095__I _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5512__I _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8059_ _3421_ _3812_ _3814_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5091__S0 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6732__A1 _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4798__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5138__I2 _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7288__A2 _3123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7902__I _3417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7212__A2 _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5223__A1 _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5760_ reg_file.reg_storage\[12\]\[10\] reg_file.reg_storage\[13\]\[10\] reg_file.reg_storage\[14\]\[10\]
+ reg_file.reg_storage\[15\]\[10\] _0686_ _1657_ _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_69_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6971__A1 _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5774__A2 _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6253__I _2086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5691_ _1606_ _1607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4711_ net7 _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7430_ _3260_ _3261_ _3262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4642_ _0485_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_126_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7361_ _3157_ net102 _3158_ _3198_ _3199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4573_ _0498_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_24_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9100_ _4460_ _4486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7292_ _3122_ _3112_ _3134_ _3135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6312_ _2143_ _2222_ _2105_ _2223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_110_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9031_ _4404_ _4443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6243_ _2154_ _2155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5533__S _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8779__A2 _4288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6174_ _2086_ _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5137__S1 _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5125_ _1031_ _1040_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_137_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6872__B _2764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5056_ _0950_ _0951_ _0971_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_79_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4648__S0 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7203__A2 _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8815_ reg_file.reg_storage\[10\]\[1\] _4313_ _4314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6163__I _2076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5958_ _1495_ _1874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5765__A2 _1671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8746_ _4195_ _4262_ _4271_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4909_ _0824_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8677_ _4180_ _4223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5889_ _1804_ _1762_ _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_132_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6714__A1 _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7628_ _3431_ _3446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_51_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7559_ net89 _1381_ _3380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9539__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9229_ _0015_ clknet_leaf_13_clk reg_file.reg_storage\[5\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8818__I _4315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5540__I2 _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7442__A2 _3262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9195__A2 _4513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5205__A1 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8242__I1 _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8942__A2 _4386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6705__A1 _2573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_132_clk clknet_4_4_0_clk clknet_leaf_132_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_124_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer17 _1493_ net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer28 _0511_ net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6930_ _2246_ _2819_ _2820_ _2821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__9186__A2 _4536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6861_ _2038_ _2752_ _2753_ _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8600_ reg_file.reg_storage\[12\]\[29\] _4162_ _4167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9580_ _0366_ clknet_leaf_65_clk reg_file.reg_storage\[9\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8933__A2 _4381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6792_ _2684_ _2671_ _2574_ _2687_ _2688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5812_ _1723_ _1725_ _1726_ _1727_ _1595_ _1596_ _1728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ reg_file.reg_storage\[2\]\[11\] reg_file.reg_storage\[3\]\[11\] _1614_ _1659_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8531_ _4125_ _4126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6795__I1 _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5674_ _0566_ _1590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8462_ reg_file.reg_storage\[13\]\[6\] _4076_ _4084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_123_clk clknet_4_5_0_clk clknet_leaf_123_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8839__S _4322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8393_ _4041_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4625_ reg_file.reg_storage\[2\]\[4\] reg_file.reg_storage\[3\]\[4\] _0502_ _0547_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7413_ _3209_ net106 _3247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7344_ _2969_ _1704_ _1705_ _3183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_41_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4556_ net14 _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_130_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9110__A2 _4461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7121__A1 _1690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5263__S _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7275_ _3100_ net126 _3101_ _3119_ _3120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9014_ _3963_ _4430_ _4433_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6226_ _2059_ _2139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7672__A2 _3089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4730__I0 reg_file.reg_storage\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5683__A1 _1586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6157_ _2049_ _0677_ _2070_ _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5108_ reg_file.reg_storage\[8\]\[31\] reg_file.reg_storage\[9\]\[31\] reg_file.reg_storage\[10\]\[31\]
+ reg_file.reg_storage\[11\]\[31\] _0896_ _0961_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__8621__A1 reg_file.reg_storage\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6088_ _2001_ _2002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5039_ reg_file.reg_storage\[1\]\[19\] _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7975__A3 _3761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7188__A1 _3035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output105_I net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6935__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8729_ _4259_ _4260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_114_clk clknet_4_13_0_clk clknet_leaf_114_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_36_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5046__S0 _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__I reg_file.reg_storage\[1\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9101__A2 _4486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7112__A1 net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7663__A2 _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6068__I _1982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput97 net97 mem_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_37_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8612__A1 reg_file.reg_storage\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7179__A1 _1982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__I1 reg_file.reg_storage\[9\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5285__S0 _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5729__A2 _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6926__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_105_clk clknet_4_13_0_clk clknet_leaf_105_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5037__S0 _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5588__S1 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5147__I _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5390_ reg_file.reg_storage\[4\]\[2\] reg_file.reg_storage\[5\]\[2\] reg_file.reg_storage\[6\]\[2\]
+ reg_file.reg_storage\[7\]\[2\] _0809_ _1301_ _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_50_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4986__I _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7060_ _2139_ _2730_ _2946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8394__S _4028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6011_ _1269_ _1923_ _1925_ _1926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_118_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5417__A1 _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7962_ _3750_ _3751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6913_ _2725_ _2787_ _2795_ _2804_ net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_7893_ _3660_ _3689_ _3690_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8906__A2 _4362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9632_ _0418_ clknet_leaf_129_clk reg_file.reg_storage\[4\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6844_ _2256_ _2682_ _2737_ _2738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6917__A1 _2797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9563_ _0349_ clknet_leaf_99_clk reg_file.reg_storage\[10\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6775_ _2670_ _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6393__A2 _2301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7537__I _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8514_ _4004_ _4111_ _4113_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_99_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_9494_ _0280_ clknet_leaf_108_clk reg_file.reg_storage\[8\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5726_ _0567_ _1642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_73_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5440__I1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8445_ _3425_ _4021_ _4072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5657_ reg_file.reg_storage\[12\]\[22\] reg_file.reg_storage\[13\]\[22\] reg_file.reg_storage\[14\]\[22\]
+ reg_file.reg_storage\[15\]\[22\] _1387_ _1569_ _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_60_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7342__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5057__I _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5588_ reg_file.reg_storage\[8\]\[29\] reg_file.reg_storage\[9\]\[29\] reg_file.reg_storage\[10\]\[29\]
+ reg_file.reg_storage\[11\]\[29\] _1418_ _1489_ _1504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_41_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6597__B _1963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input66_I pc[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4608_ _0528_ _0531_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8376_ reg_file.reg_storage\[14\]\[4\] _4026_ _4032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7327_ _3165_ _3166_ _3167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7258_ _3103_ _3104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6209_ _2121_ _2122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7189_ _3040_ _3041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_5_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7447__I _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6351__I _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer8 net121 net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7884__A2 _3658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7636__A2 _3446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4890_ _0624_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__7572__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6560_ _2027_ _2187_ _2464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5511_ _1426_ _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_82_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6491_ _2316_ _2391_ _2396_ _2397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5442_ _1357_ _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8230_ _3920_ _3921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8161_ _3502_ _3869_ _3878_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5373_ _1284_ _1286_ _1287_ _1288_ _0964_ _0946_ _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_11_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6210__B _2122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7112_ net145 _2988_ _2991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8092_ _3835_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5638__A1 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7043_ _1874_ _2928_ _2929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8916__I _4360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8994_ _4422_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7945_ _3588_ _2977_ _3029_ _3713_ _3736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8651__I _3555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7876_ reg_file.reg_storage\[5\]\[20\] _3658_ _3676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9615_ _0401_ clknet_leaf_63_clk reg_file.reg_storage\[1\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6827_ _1848_ _2670_ _2674_ _2564_ _2721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_77_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7563__A1 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9546_ _0332_ clknet_leaf_2_clk reg_file.reg_storage\[10\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6758_ _2634_ _2429_ _2655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5709_ reg_file.reg_storage\[2\]\[17\] reg_file.reg_storage\[3\]\[17\] _0577_ _1625_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9477_ _0263_ clknet_leaf_41_clk reg_file.reg_storage\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6689_ _2585_ _2588_ _2326_ _2589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8428_ _4017_ _4061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8359_ _4016_ _4019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5877__B2 _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7079__B1 _2542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5515__I _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5451__S _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8043__A2 _3799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__A1 _1604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5652__I1 _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A2 _2231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7306__A1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8002__S _3775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7857__A2 _3658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8282__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8736__I _4265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5096__A2 _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6293__A1 _1765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6256__I _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _1902_ _1905_ _1906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_115_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ reg_file.reg_storage\[4\]\[23\] reg_file.reg_storage\[5\]\[23\] reg_file.reg_storage\[6\]\[23\]
+ reg_file.reg_storage\[7\]\[23\] _0855_ _0857_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_59_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7730_ _3048_ _3136_ _3497_ _1829_ _3472_ _3541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_86_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7661_ net123 _3432_ _3474_ _3476_ _3477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_46_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9400_ _0186_ clknet_leaf_90_clk reg_file.reg_storage\[14\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4873_ _0762_ _0777_ _0782_ _0783_ _0786_ _0788_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6612_ _2513_ _2514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7592_ _3411_ _3412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_61_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5536__S _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9331_ _0117_ clknet_leaf_74_clk reg_file.reg_storage\[6\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6543_ _1959_ _2416_ _2446_ _1194_ _2447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_9262_ _0048_ clknet_leaf_46_clk reg_file.reg_storage\[3\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6474_ _2110_ _2071_ _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_15_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8213_ reg_file.reg_storage\[6\]\[29\] _3903_ _3908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5403__S0 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5425_ _1241_ _1298_ _1340_ _1111_ _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_113_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9193_ _3983_ _4538_ _4542_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6520__A2 _2335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8144_ _3866_ _3867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5356_ reg_file.reg_storage\[4\]\[5\] reg_file.reg_storage\[5\]\[5\] reg_file.reg_storage\[6\]\[5\]
+ reg_file.reg_storage\[7\]\[5\] _0770_ _1271_ _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5287_ _1196_ _1200_ _1201_ _1202_ _0821_ _0787_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_8075_ reg_file.reg_storage\[2\]\[5\] _3491_ _3822_ _3826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_89_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7026_ _2906_ _2912_ _2076_ _2913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8025__A2 _3789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input29_I inst[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_94_clk clknet_4_15_0_clk clknet_leaf_94_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__A1 _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8977_ _4409_ _4412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7928_ _3400_ _3719_ _3721_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4598__A1 _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4988__I3 reg_file.reg_storage\[15\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7859_ _3427_ _3660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__S0 _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9529_ _0315_ clknet_leaf_101_clk reg_file.reg_storage\[11\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output97_I net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8757__S _4272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5078__A2 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5322__I0 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9213__A1 _4012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_85_clk clknet_4_14_0_clk clknet_leaf_85_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8016__A2 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6578__A2 _2450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8291__I _3648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7527__A1 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5002__A2 reg_file.reg_storage\[1\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5633__S0 _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_54_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5210_ reg_file.reg_storage\[1\]\[12\] _1125_ _1123_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6190_ _1028_ _2103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5141_ _1056_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4994__I _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _0957_ reg_file.reg_storage\[2\]\[28\] _0807_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8900_ _4365_ _4366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_leaf_76_clk clknet_4_9_0_clk clknet_leaf_76_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6018__A1 _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8831_ _4323_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_84_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8762_ _4280_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7713_ _0594_ _3524_ _3525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5974_ _1401_ _1519_ _1889_ _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_48_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4925_ reg_file.reg_storage\[1\]\[22\] _0840_ _0837_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8693_ _3695_ _4234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7644_ _3022_ _3461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_129_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4856_ _0771_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7575_ _3394_ _3395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6741__A2 _2638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6526_ _2002_ _2423_ _2430_ _2431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9314_ _0100_ clknet_leaf_18_clk reg_file.reg_storage\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4787_ _0702_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9245_ _0031_ clknet_leaf_114_clk reg_file.reg_storage\[5\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8494__A2 _4101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _1228_ _2363_ _1960_ _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9176_ reg_file.reg_storage\[15\]\[15\] _3623_ _4515_ _4533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5408_ net76 _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6388_ _2104_ _2297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8127_ _3726_ _3854_ _3855_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5339_ reg_file.reg_storage\[4\]\[6\] reg_file.reg_storage\[5\]\[6\] reg_file.reg_storage\[6\]\[6\]
+ reg_file.reg_storage\[7\]\[6\] _0860_ _0818_ _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__8246__A2 _3924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_126_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5014__B _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8058_ reg_file.reg_storage\[2\]\[0\] _3813_ _3814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output135_I net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_67_clk clknet_4_11_0_clk clknet_leaf_67_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7009_ _2333_ _2895_ _2896_ _2897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_98_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5949__B _1580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7757__A1 _2438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6980__A2 _2659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7509__A1 _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5091__S1 _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6732__A2 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8485__A2 _4088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5138__I3 _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_58_clk clknet_4_10_0_clk clknet_leaf_58_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_88_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6534__I _2438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4982__A1 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5690_ _1605_ _1606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_57_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4710_ net11 _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_62_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4641_ reg_file.reg_storage\[4\]\[5\] reg_file.reg_storage\[5\]\[5\] reg_file.reg_storage\[6\]\[5\]
+ reg_file.reg_storage\[7\]\[5\] _0556_ _0557_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__7920__A1 _3447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6723__A2 _2595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7360_ _3196_ _3197_ _3198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4572_ net14 _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7291_ net96 _3134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6311_ _1944_ _1936_ _2222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9030_ _3986_ _4412_ _4442_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6242_ _1109_ _1239_ _0883_ _0793_ _2154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_0_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_71_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6173_ _0733_ _2086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5124_ _0891_ _1039_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_49_clk clknet_4_10_0_clk clknet_leaf_49_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__9610__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5055_ _0969_ _0970_ _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7739__A1 _3447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6444__I _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8814_ _4309_ _4313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8400__A2 _4044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__S1 _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8745_ reg_file.reg_storage\[11\]\[6\] _4263_ _4271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5957_ _1478_ _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8676_ _3656_ _4222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_80_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6962__A2 _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4908_ _0823_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7627_ _3428_ _3443_ _3445_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input96_I pc[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5888_ net18 _1115_ _1479_ _1804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_117_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4839_ _0627_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6175__B1 _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ _3372_ _3375_ _3379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6509_ _1681_ net208 _2157_ _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7489_ net82 _1404_ _3316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_9228_ _0014_ clknet_leaf_61_clk reg_file.reg_storage\[5\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__S _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5540__I3 _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9159_ _4523_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_54_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8834__I _4310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_119_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_106_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_83_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8458__A2 _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_128_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_117_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6469__A1 _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_98_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4575__S0 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6641__A1 _2103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer18 _0564_ net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_137_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xrebuffer29 _2317_ net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_77_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6860_ _2122_ _2707_ _2753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6791_ _2685_ _2577_ _2686_ _2687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5811_ reg_file.reg_storage\[4\]\[15\] reg_file.reg_storage\[5\]\[15\] reg_file.reg_storage\[6\]\[15\]
+ reg_file.reg_storage\[7\]\[15\] _1615_ _1672_ _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_128_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5742_ reg_file.reg_storage\[8\]\[11\] reg_file.reg_storage\[9\]\[11\] reg_file.reg_storage\[10\]\[11\]
+ reg_file.reg_storage\[11\]\[11\] _1358_ _1657_ _1658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_91_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5809__S _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8530_ _4021_ _4124_ _4125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5673_ reg_file.reg_storage\[8\]\[16\] reg_file.reg_storage\[9\]\[16\] reg_file.reg_storage\[10\]\[16\]
+ reg_file.reg_storage\[11\]\[16\] _1587_ _1588_ _1589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_72_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6213__B _2125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8461_ _4083_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8392_ reg_file.reg_storage\[14\]\[11\] _3951_ _4035_ _4041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4624_ reg_file.reg_storage\[8\]\[4\] reg_file.reg_storage\[9\]\[4\] reg_file.reg_storage\[10\]\[4\]
+ reg_file.reg_storage\[11\]\[4\] _0496_ _0499_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7412_ _3238_ _3245_ _3246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_41_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7343_ _3180_ _3181_ _3182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4555_ _0480_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_130_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9013_ reg_file.reg_storage\[1\]\[16\] _4424_ _4433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_92_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7274_ _3113_ _3116_ _3118_ _3119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_110_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_109_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6225_ _2134_ _2137_ _2081_ _2138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4730__I1 reg_file.reg_storage\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5683__A2 _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6156_ _1311_ _1337_ _2018_ _2070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5107_ reg_file.reg_storage\[12\]\[31\] reg_file.reg_storage\[13\]\[31\] reg_file.reg_storage\[14\]\[31\]
+ reg_file.reg_storage\[15\]\[31\] _1021_ _1022_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__8654__I _3566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6087_ _1120_ _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5038_ _0774_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input11_I inst[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6174__I _2086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6989_ _2352_ _2863_ _2871_ _2877_ _2878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8728_ _3761_ _4178_ _4259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4946__A1 _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8688__A2 _4223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8659_ _4210_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5046__S1 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8829__I _4310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8860__A2 _4336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6349__I _2258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput98 net98 mem_addr[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_37_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6084__I _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5285__S1 _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__A1 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8679__A2 _4214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5037__S1 _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8851__A2 _4331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6259__I _2170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6862__A1 _2217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6010_ _1029_ _1183_ _1924_ _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input3_I inst[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5417__A2 _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7961_ net211 _3728_ _3729_ _3748_ _3749_ _3750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__4720__S0 _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7892_ reg_file.reg_storage\[5\]\[22\] _3458_ _3690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6912_ _1104_ _2796_ _2803_ _2804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6843_ _0848_ _1853_ _2345_ _2736_ _2737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_9631_ _0417_ clknet_leaf_18_clk reg_file.reg_storage\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7818__I _3622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9562_ _0348_ clknet_leaf_99_clk reg_file.reg_storage\[10\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8119__A1 _3705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6774_ _1116_ _1564_ _2669_ _2670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_57_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8513_ reg_file.reg_storage\[13\]\[28\] _4109_ _4113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5725_ reg_file.reg_storage\[12\]\[19\] reg_file.reg_storage\[13\]\[19\] reg_file.reg_storage\[14\]\[19\]
+ reg_file.reg_storage\[15\]\[19\] _0685_ _1623_ _1641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_9493_ _0279_ clknet_leaf_119_clk reg_file.reg_storage\[8\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8444_ _3912_ _4069_ _4071_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5028__S1 _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5656_ reg_file.reg_storage\[1\]\[22\] _1571_ _1569_ _1572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4607_ _0529_ _0530_ _0508_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7342__A2 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5587_ reg_file.reg_storage\[12\]\[29\] reg_file.reg_storage\[13\]\[29\] reg_file.reg_storage\[14\]\[29\]
+ reg_file.reg_storage\[15\]\[29\] _1418_ _1489_ _1503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_115_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8375_ _4031_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7326_ _3145_ _3154_ _3133_ _3166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input59_I mem_ld_dat[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7257_ net93 _3102_ _3103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6853__A1 _2742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6208_ _2097_ _2121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7188_ _3035_ _3039_ _3040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6605__A1 _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6139_ _2048_ _2051_ _2052_ _2053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_5_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6632__I _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7030__A1 _2036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5592__A1 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer9 _1742_ net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7333__A2 _3161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7463__I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6392__I0 _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5895__A2 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7097__A1 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8349__A1 reg_file.reg_storage\[7\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9010__A2 _4430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5510_ _1425_ _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8521__A1 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7324__A2 _3156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6490_ _2394_ _2395_ _2396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_140_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8469__I _4073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5441_ _0534_ _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_42_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8160_ reg_file.reg_storage\[6\]\[6\] _3870_ _3878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5372_ reg_file.reg_storage\[8\]\[4\] reg_file.reg_storage\[9\]\[4\] reg_file.reg_storage\[10\]\[4\]
+ reg_file.reg_storage\[11\]\[4\] _1020_ _0902_ _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_2_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7111_ net212 _2989_ _2990_ net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8091_ reg_file.reg_storage\[2\]\[12\] _3585_ _3821_ _3835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5822__S _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5638__A2 _1553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7042_ _2907_ _2927_ _2928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8824__A2 _4312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5621__I _1536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8993_ reg_file.reg_storage\[1\]\[7\] _3510_ _4421_ _4422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8052__A3 _3394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7944_ _3722_ _3734_ _3735_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6063__A2 _1902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7875_ _3674_ _3675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9001__A2 _4406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__S _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9614_ _0400_ clknet_leaf_62_clk reg_file.reg_storage\[1\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6826_ _2668_ _2677_ _2700_ _2718_ _2719_ _2720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_9545_ _0331_ clknet_leaf_52_clk reg_file.reg_storage\[10\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6757_ _2652_ _2653_ _2654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5708_ reg_file.reg_storage\[8\]\[17\] reg_file.reg_storage\[9\]\[17\] reg_file.reg_storage\[10\]\[17\]
+ reg_file.reg_storage\[11\]\[17\] _0658_ _1623_ _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5068__I _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6688_ _2469_ _2587_ _2120_ _2588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9476_ _0262_ clknet_leaf_120_clk reg_file.reg_storage\[8\]\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8427_ _3996_ _4018_ _4060_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5639_ _1400_ _1552_ _1554_ _1555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8358_ _4017_ _4018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output165_I net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7079__B2 _2682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7309_ _3149_ _3150_ _3151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8289_ reg_file.reg_storage\[7\]\[16\] _3947_ _3965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8815__A2 _4313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5404__I2 _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8503__A1 reg_file.reg_storage\[13\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7306__A2 _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9224__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4610__I _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6738__S _2335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7921__I _3047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5441__I _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8752__I _4260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _1795_ net227 _1904_ _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_86_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4941_ _0856_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7660_ net129 _3475_ _3476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4872_ _0787_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_24_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6611_ _2510_ _2512_ _2513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7591_ _3026_ _3411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9330_ _0116_ clknet_4_9_0_clk reg_file.reg_storage\[6\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6542_ _1667_ _2414_ _2446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_42_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9261_ _0047_ clknet_leaf_35_clk reg_file.reg_storage\[3\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6473_ _2379_ net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5616__I _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8212_ _3734_ _3905_ _3907_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9192_ reg_file.reg_storage\[15\]\[22\] _4511_ _4542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput200 net200 pc_next[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5403__S1 _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ _1299_ _1323_ _1339_ _1241_ _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_101_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8143_ _3424_ _3865_ _3866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8927__I _4361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5355_ _0640_ _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_7_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5286_ reg_file.reg_storage\[8\]\[10\] reg_file.reg_storage\[9\]\[10\] reg_file.reg_storage\[10\]\[10\]
+ reg_file.reg_storage\[11\]\[10\] _0839_ _0760_ _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8074_ _3478_ _3818_ _3825_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7025_ _1508_ _2912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8976_ _4410_ _4411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7927_ reg_file.reg_storage\[5\]\[26\] _3720_ _3721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7278__I net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7858_ _3600_ _3657_ _3659_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6809_ _2209_ _2704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7789_ _3587_ _3595_ _3596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5642__S1 _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9528_ _0314_ clknet_leaf_106_clk reg_file.reg_storage\[11\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9459_ _0245_ clknet_leaf_74_clk reg_file.reg_storage\[12\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_100_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5330__S0 _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5786__A1 _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8013__S _3768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5633__S1 _1483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4600__I3 reg_file.reg_storage\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5436__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5397__S0 _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5880__B _1795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8747__I _4260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5140_ _1046_ _0937_ _0835_ _1055_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_5071_ _0768_ reg_file.reg_storage\[3\]\[28\] _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5077__I0 _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8830_ reg_file.reg_storage\[10\]\[7\] _4197_ _4322_ _4323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7215__B2 _3064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5973_ _1401_ _1511_ _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8761_ reg_file.reg_storage\[11\]\[13\] _4211_ _4265_ _4280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7712_ _3506_ _3513_ _3524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4924_ reg_file.reg_storage\[2\]\[22\] reg_file.reg_storage\[3\]\[22\] _0839_ _0840_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8692_ _4232_ _4226_ _4233_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7518__A2 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8191__A2 _3893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7643_ _3416_ _3460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4855_ _0770_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7574_ _3392_ _3393_ net3 _3394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4786_ net6 _0701_ _0691_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_144_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6525_ _2424_ _2429_ _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9313_ _0099_ clknet_leaf_130_clk reg_file.reg_storage\[6\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9244_ _0030_ clknet_leaf_103_clk reg_file.reg_storage\[5\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _2106_ _2363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9175_ _3957_ _4531_ _4532_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6387_ _2056_ _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5407_ _1311_ _1322_ _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8657__I _3583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8126_ reg_file.reg_storage\[2\]\[27\] _3852_ _3855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5338_ net93 _0798_ _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input41_I mem_ld_dat[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8057_ _3810_ _3813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_126_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5269_ reg_file.reg_storage\[2\]\[11\] reg_file.reg_storage\[3\]\[11\] _0801_ _1185_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7008_ _2360_ _2790_ _2896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output128_I net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4626__S _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7757__A2 _3504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8959_ _4243_ _4398_ _4399_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7509__A2 _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9131__A1 _4012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6087__I _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8008__S _3768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5303__S0 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4640_ reg_file.reg_storage\[12\]\[5\] reg_file.reg_storage\[13\]\[5\] reg_file.reg_storage\[14\]\[5\]
+ reg_file.reg_storage\[15\]\[5\] _0556_ _0557_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_25_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6310_ _2210_ _2213_ _2220_ _2056_ _2221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4571_ _0496_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7290_ _3132_ _3133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6198__S _2097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7684__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6241_ _2152_ _2153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6172_ _2085_ net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
X_5123_ _1032_ _1036_ _1037_ _1038_ _0786_ _0788_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_5054_ _0830_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8813_ _4311_ _4312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5214__A3 _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5956_ _1029_ _1477_ _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8744_ _4270_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8675_ _4220_ _4214_ _4221_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5887_ _1279_ _1763_ _1803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4907_ net10 _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4838_ _0753_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7626_ reg_file.reg_storage\[5\]\[1\] _3444_ _3445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6175__A1 _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7911__A2 _3705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input89_I pc[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4769_ _0572_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7557_ _3368_ _1481_ _3378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6508_ net233 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_132_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7488_ _3144_ _3305_ _3306_ _3315_ net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_113_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8387__I _4023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9227_ _0013_ clknet_leaf_9_clk reg_file.reg_storage\[5\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6439_ _2345_ _2346_ _2347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7291__I net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9158_ reg_file.reg_storage\[15\]\[7\] _3510_ _4522_ _4523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8109_ _3667_ _3844_ _3845_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6836__S _2040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9089_ reg_file.reg_storage\[4\]\[13\] _3597_ _4465_ _4480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7466__I _1553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5913__A1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8297__I _3921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6469__A2 _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4575__S1 _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5772__S0 _1606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer19 _1618_ net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6790_ _2685_ _2578_ _2686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5810_ reg_file.reg_storage\[12\]\[15\] reg_file.reg_storage\[13\]\[15\] reg_file.reg_storage\[14\]\[15\]
+ reg_file.reg_storage\[15\]\[15\] _1611_ _1672_ _1726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_29_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5741_ _1627_ _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8460_ reg_file.reg_storage\[13\]\[5\] _3935_ _4079_ _4083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5672_ _1361_ _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_45_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7411_ _3240_ _3244_ _3245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8391_ _4040_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4623_ _0545_ net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_130_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7342_ net66 net67 _3165_ _3132_ _3181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_12_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4554_ net13 _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_114_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7273_ _3104_ _3109_ _3117_ _3118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7657__A1 _3081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9012_ _1167_ _4406_ _4432_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6224_ _2059_ _2137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4730__I2 reg_file.reg_storage\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6155_ _2061_ _2064_ _2068_ _2069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5106_ _0836_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6086_ _1999_ _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5037_ reg_file.reg_storage\[4\]\[19\] reg_file.reg_storage\[5\]\[19\] reg_file.reg_storage\[6\]\[19\]
+ reg_file.reg_storage\[7\]\[19\] _0921_ _0922_ _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6455__I _2022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8670__I _3637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8727_ _4170_ _4256_ _4258_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6988_ _2113_ _2796_ _2876_ _2877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5939_ _1846_ _1851_ _1854_ _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8658_ reg_file.reg_storage\[8\]\[12\] _4209_ _4186_ _4210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8589_ _3990_ _4121_ _4160_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_134_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7609_ _3427_ _3428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output195_I net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_105_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7648__A1 _3047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput99 net99 mem_addr[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8845__I _4311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6566__S _2052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8376__A2 _4026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9176__I1 _3623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6934__I0 _2269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5444__I _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5745__S0 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5665__A3 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7960_ _3702_ _3384_ _3496_ _1381_ _3749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__4720__S1 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6911_ _1983_ _2802_ _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7891_ _3688_ _3689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9630_ _0416_ clknet_leaf_112_clk reg_file.reg_storage\[4\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6842_ _2734_ _2576_ _2735_ _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9561_ _0347_ clknet_leaf_102_clk reg_file.reg_storage\[10\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8119__A2 _3812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6773_ _1378_ _1557_ _2669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5619__I _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8512_ _4000_ _4111_ _4112_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5724_ reg_file.reg_storage\[1\]\[19\] _1639_ _0878_ _1640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9492_ _0278_ clknet_leaf_117_clk reg_file.reg_storage\[8\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8443_ reg_file.reg_storage\[13\]\[0\] _4070_ _4071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5655_ reg_file.reg_storage\[2\]\[22\] reg_file.reg_storage\[3\]\[22\] _1369_ _1571_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7834__I _3637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4606_ reg_file.reg_storage\[8\]\[2\] reg_file.reg_storage\[9\]\[2\] reg_file.reg_storage\[10\]\[2\]
+ reg_file.reg_storage\[11\]\[2\] _0495_ net229 _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8374_ reg_file.reg_storage\[14\]\[3\] _3930_ _4029_ _4031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5586_ _1468_ _1001_ _1500_ _1501_ _1502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_115_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7325_ net68 _3165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_130_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7256_ _2229_ _1383_ _3102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_111_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7187_ _3038_ _3039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6207_ _2109_ _2120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6138_ _2021_ _2052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_5_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_82_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6069_ _1907_ _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7802__A1 _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output110_I net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5416__I0 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_97_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5529__I _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_62_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5592__A2 _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_20_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__S0 _1590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_35_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__A2 _2682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8046__A1 _3740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9149__I1 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_108_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _1353_ net19 _1355_ _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ reg_file.reg_storage\[12\]\[4\] reg_file.reg_storage\[13\]\[4\] reg_file.reg_storage\[14\]\[4\]
+ reg_file.reg_storage\[15\]\[4\] _1020_ _0902_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7110_ net134 _2988_ _2990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8090_ _3834_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7041_ _2912_ _2537_ _2927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8992_ _4414_ _4421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_2_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7943_ reg_file.reg_storage\[5\]\[28\] _3720_ _3735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7260__A2 _3090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5110__I2 _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7874_ net109 _3661_ _3670_ _3673_ _3674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_6825_ _0829_ _2699_ _2719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9613_ _0399_ clknet_leaf_35_clk reg_file.reg_storage\[1\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5349__I _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9544_ _0330_ clknet_leaf_53_clk reg_file.reg_storage\[10\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6756_ _2616_ _2629_ _2632_ _2653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5707_ _0570_ _1623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6687_ _2523_ _2586_ _2105_ _2587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9475_ _0261_ clknet_leaf_135_clk reg_file.reg_storage\[8\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8426_ reg_file.reg_storage\[14\]\[26\] _4059_ _4060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5638_ _1116_ _1553_ _1554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input71_I pc[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8357_ _4016_ _4017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5569_ _1419_ reg_file.reg_storage\[3\]\[30\] _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7308_ net66 _1671_ _3150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8288_ _3963_ _3964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output158_I net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8028__A1 _3682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7239_ _3077_ _3080_ _3086_ net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_129_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8579__A2 _4154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5637__I0 _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6817__A2 _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5253__A1 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4940_ _0641_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8990__A2 _4412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4871_ _0649_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7590_ _3023_ _3410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6610_ _2398_ _2511_ _2512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8742__A2 _4262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6541_ _2402_ _2415_ _2445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_28_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9260_ _0046_ clknet_leaf_46_clk reg_file.reg_storage\[3\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6472_ _2352_ _2357_ _2359_ _2259_ _2378_ _2379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_43_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8211_ reg_file.reg_storage\[6\]\[28\] _3903_ _3907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9191_ _3980_ _4538_ _4541_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput201 net201 pc_next[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5423_ _1337_ _1338_ _0973_ _1339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8142_ _3389_ _3807_ _3395_ _3865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_2_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5354_ net92 _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_140_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5285_ reg_file.reg_storage\[12\]\[10\] reg_file.reg_storage\[13\]\[10\] reg_file.reg_storage\[14\]\[10\]
+ reg_file.reg_storage\[15\]\[10\] _0839_ _0760_ _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_49_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8073_ reg_file.reg_storage\[2\]\[4\] _3819_ _3825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7024_ _2909_ _2910_ _2911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8975_ _4409_ _4410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5244__A1 _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7926_ _3398_ _3720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6992__A1 _2856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5634__I3 reg_file.reg_storage\[7\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7857_ reg_file.reg_storage\[5\]\[18\] _3658_ _3659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_136_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6808_ _2700_ _2702_ _2703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_34_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8733__A2 _4263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7788_ _3572_ _3182_ _3573_ _3593_ _3594_ _3595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_9527_ _0313_ clknet_leaf_108_clk reg_file.reg_storage\[11\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6739_ _2586_ _2636_ _2007_ _2637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9458_ _0244_ clknet_leaf_74_clk reg_file.reg_storage\[12\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4711__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8409_ _3970_ _4044_ _4050_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5743__S _1614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9389_ _0175_ clknet_leaf_12_clk reg_file.reg_storage\[14\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5235__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8972__A2 _4407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5330__S1 _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6983__A1 _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5786__A2 _1701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6735__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5397__S1 _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5452__I _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5070_ reg_file.reg_storage\[1\]\[28\] _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5849__I0 net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8763__I _4261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7215__A2 net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7600__C _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5972_ _1876_ _1886_ _1887_ _1888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8760_ _4279_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7711_ _3434_ _3516_ _3520_ _3522_ _3523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4923_ _0633_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_129_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8691_ reg_file.reg_storage\[8\]\[22\] _4181_ _4233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7642_ _3459_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4854_ _0627_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_117_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7573_ _0609_ _0600_ _0611_ _0664_ _3393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4785_ _0700_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_31_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9312_ _0098_ clknet_leaf_133_clk reg_file.reg_storage\[6\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6524_ _2300_ _2428_ _2198_ _2429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9243_ _0029_ clknet_leaf_103_clk reg_file.reg_storage\[5\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7151__A1 net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6455_ _2022_ _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9174_ reg_file.reg_storage\[15\]\[14\] _4525_ _4532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6386_ _2284_ _2287_ _2294_ _2295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5790__C _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5406_ _1312_ _1321_ _1282_ _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8125_ _3811_ _3854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__I _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5337_ _0831_ _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5268_ reg_file.reg_storage\[4\]\[11\] reg_file.reg_storage\[5\]\[11\] reg_file.reg_storage\[6\]\[11\]
+ reg_file.reg_storage\[7\]\[11\] _0779_ _0942_ _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8056_ _3811_ _3812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input34_I mem_ld_dat[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8673__I _3648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7007_ _2117_ _2842_ _2894_ _2362_ _2895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5199_ _0978_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5217__A1 _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7206__A2 _1982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8958_ reg_file.reg_storage\[9\]\[27\] _4396_ _4399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7909_ _3704_ _3705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8889_ _4354_ _4357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5076__S0 _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9131__A2 _4457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8890__A1 reg_file.reg_storage\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6317__B _2221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8945__A2 _4388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5303__S1 _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6831__I _2404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_135_clk clknet_4_4_0_clk clknet_leaf_135_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5447__I _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4570_ _0495_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_25_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9122__A2 _4496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7662__I _3477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7684__A2 _3138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6240_ _1903_ _0730_ _2152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_110_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6171_ _1984_ _1996_ _2084_ _2085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_21_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ reg_file.reg_storage\[8\]\[30\] reg_file.reg_storage\[9\]\[30\] reg_file.reg_storage\[10\]\[30\]
+ reg_file.reg_storage\[11\]\[30\] _0811_ _0761_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_20_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4727__S _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5053_ _0968_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__9189__A2 _4538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8812_ _4310_ _4311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ _1842_ _1869_ _1870_ _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8743_ reg_file.reg_storage\[11\]\[5\] _4193_ _4266_ _4270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8674_ reg_file.reg_storage\[8\]\[17\] _4203_ _4221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4906_ _0821_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_48_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_126_clk clknet_4_5_0_clk clknet_leaf_126_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5886_ _1778_ _1799_ _1801_ _1802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7625_ _3426_ _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4837_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6175__B3 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6175__A2 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9113__A2 _4463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7556_ _3144_ _3370_ _3371_ _3377_ net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4768_ _0683_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_132_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7124__A1 net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5293__S _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6507_ _2342_ _2386_ _2390_ _2412_ _2413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4699_ _0614_ _0602_ _0603_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_7487_ _3053_ _3314_ _3315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9226_ _0012_ clknet_leaf_7_clk reg_file.reg_storage\[5\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6438_ _2343_ _1827_ _2268_ _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_30_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9157_ _4510_ _4522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5686__A1 _1580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6188__I _2040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8108_ reg_file.reg_storage\[2\]\[19\] _3842_ _3845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6369_ _1809_ _2277_ _2278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_output140_I net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9088_ _4479_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8039_ _3719_ _3757_ _3800_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_106_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5297__S0 _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_117_clk clknet_4_1_0_clk clknet_leaf_117_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_65_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5267__I _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9104__A2 _4486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7115__A1 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5772__S1 _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8615__A1 _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5429__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9040__A1 _3999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8918__A2 _4362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6929__A1 _2217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_108_clk clknet_4_13_0_clk clknet_leaf_108_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5740_ _1380_ _1652_ _1655_ _1656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_9_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5671_ _1357_ _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_84_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7410_ _3243_ _3244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8390_ reg_file.reg_storage\[14\]\[10\] _3949_ _4035_ _4040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_96_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4622_ _0488_ _0544_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_80_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7341_ net69 _3180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7392__I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7272_ _3097_ _3102_ _3117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7657__A2 _3403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9011_ _3623_ _4405_ _4432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6223_ _2134_ _2135_ _2077_ _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__S0 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4730__I3 reg_file.reg_storage\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6154_ _2065_ _2067_ _2068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_57_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5105_ _1020_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6085_ _1998_ _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6736__I _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5036_ net75 _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__7680__I2 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8909__A2 _4363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6987_ _2174_ _2874_ _2875_ _2876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7567__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6396__A2 _2304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8726_ reg_file.reg_storage\[11\]\[0\] _4257_ _4258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5938_ _1852_ _1853_ _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ _1242_ _1253_ _1785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8657_ _3583_ _4209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8588_ reg_file.reg_storage\[12\]\[24\] _4122_ _4160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_134_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7608_ _3426_ _3427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8398__I _4024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output188_I net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7539_ _3345_ _3346_ _3362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_32_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7648__A2 _3068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9209_ _4006_ _4548_ _4551_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8073__A2 _3819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7281__B1 _3102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7678__S _3492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_9_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6934__I1 _2080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5745__S1 _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5122__I0 reg_file.reg_storage\[8\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6075__A1 _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9013__A1 reg_file.reg_storage\[1\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7890_ net111 _3661_ _3685_ _3687_ _3688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_6910_ _2797_ _2798_ _2266_ _2801_ _2802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XPHY_EDGE_ROW_59_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6841_ _2734_ _2304_ _2735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9560_ _0346_ clknet_leaf_106_clk reg_file.reg_storage\[10\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6622__I0 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8511_ reg_file.reg_storage\[13\]\[27\] _4109_ _4112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5681__S0 _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6772_ _2561_ _2663_ _2667_ _2668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_58_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5723_ reg_file.reg_storage\[2\]\[19\] reg_file.reg_storage\[3\]\[19\] _1357_ _1639_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9491_ _0277_ clknet_leaf_77_clk reg_file.reg_storage\[8\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8442_ _4067_ _4070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5654_ reg_file.reg_storage\[8\]\[22\] reg_file.reg_storage\[9\]\[22\] reg_file.reg_storage\[10\]\[22\]
+ reg_file.reg_storage\[11\]\[22\] _1463_ _1569_ _1570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4605_ reg_file.reg_storage\[12\]\[2\] reg_file.reg_storage\[13\]\[2\] reg_file.reg_storage\[14\]\[2\]
+ reg_file.reg_storage\[15\]\[2\] _0495_ net229 _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8373_ _4030_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5585_ _1431_ reg_file.reg_storage\[2\]\[29\] _1486_ _1501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_68_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7324_ _3121_ _3156_ _3164_ net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _3052_ _3101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6206_ _2117_ _1961_ _2118_ _2119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7186_ _0701_ _3037_ _1410_ _3038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__6466__I _2080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6137_ _2049_ _1206_ _2050_ _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_99_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6068_ _1982_ net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_77_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5813__A1 _1604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5019_ _0908_ _0910_ _0934_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8681__I _4187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output103_I net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6369__A2 _2277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_24_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9689_ _0475_ clknet_leaf_94_clk reg_file.reg_storage\[15\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8709_ _4243_ _4244_ _4245_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_86_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_133_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4942__I3 reg_file.reg_storage\[7\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8294__A2 _3959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__S1 _1642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_95_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9094__I1 _3623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6057__A1 _1795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5415__S0 _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5370_ reg_file.reg_storage\[1\]\[4\] _1285_ _1141_ _1286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7670__I _3484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7040_ _1041_ _2926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6048__A1 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5190__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8991_ _3937_ _4411_ _4420_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7942_ _3733_ _3734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_2_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9612_ _0398_ clknet_leaf_63_clk reg_file.reg_storage\[1\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6235__B _2147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7873_ _3671_ _3262_ _3634_ _3672_ _3673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6824_ _1849_ _2676_ _2699_ _0829_ _2718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__6220__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6755_ _0969_ _2651_ _2652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_9543_ _0329_ clknet_leaf_27_clk reg_file.reg_storage\[10\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5654__S0 _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9474_ _0260_ clknet_leaf_120_clk reg_file.reg_storage\[8\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5706_ _0488_ _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_9_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8425_ _4016_ _4059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_30_clk clknet_4_3_0_clk clknet_leaf_30_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6686_ _0934_ _1176_ _2586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_6_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5637_ _1438_ _1353_ _1412_ _1553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6523__A2 _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input64_I mem_ld_dat[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5568_ reg_file.reg_storage\[4\]\[30\] reg_file.reg_storage\[5\]\[30\] reg_file.reg_storage\[6\]\[30\]
+ reg_file.reg_storage\[7\]\[30\] _1482_ _1483_ _1484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8356_ _3809_ _4015_ _4016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8287_ _3637_ _3963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8676__I _3656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7307_ _3147_ _3141_ _3148_ _3149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7238_ _3059_ net123 _3061_ _3085_ _3086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5499_ net20 _1402_ _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6196__I _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_97_clk clknet_4_15_0_clk clknet_leaf_97_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_129_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7169_ _2969_ _2975_ _1900_ _3025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_95_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8028__A2 _3791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4709__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7787__A1 _3184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8200__A2 _3870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6211__A1 _2120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5645__S0 _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5476__S _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7490__I net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6817__A3 _2224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_88_clk clknet_4_14_0_clk clknet_leaf_88_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__9067__I1 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _0785_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_87_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6540_ _2443_ _2444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__7665__I net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_12_clk clknet_4_0_0_clk clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5159__I3 reg_file.reg_storage\[7\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6471_ _2342_ _2370_ _2377_ _2378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8210_ _3726_ _3905_ _3906_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_81_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9190_ reg_file.reg_storage\[15\]\[21\] _4536_ _4541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5422_ _0678_ _1030_ _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_140_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8141_ _3421_ _3862_ _3864_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput202 net202 pc_next[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5353_ _1268_ _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_96_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5284_ _0814_ _1197_ _1198_ _1199_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8072_ _3824_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9207__A1 _4003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_79_clk clknet_4_12_0_clk clknet_leaf_79_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7023_ _2885_ _2890_ _2883_ _2910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6441__A1 _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8974_ _3760_ _3387_ _3425_ _4409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5244__A2 _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7925_ _3718_ _3719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7856_ _3457_ _3658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_34_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6807_ _2701_ _2679_ _2702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7941__A1 net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ reg_file.reg_storage\[2\]\[16\] _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9526_ _0312_ clknet_leaf_109_clk reg_file.reg_storage\[11\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7575__I _3394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7787_ _3184_ _3438_ _3466_ _3594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_34_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6738_ _2616_ _2593_ _2335_ _2636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8497__A2 _4099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9457_ _0243_ clknet_leaf_31_clk reg_file.reg_storage\[12\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6669_ _2561_ _2567_ _2568_ _2569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9388_ _0174_ clknet_leaf_54_clk reg_file.reg_storage\[14\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_49_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8408_ reg_file.reg_storage\[14\]\[18\] _4049_ _4050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8339_ _3733_ _4003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_111_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_107_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5483__A2 _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6432__A1 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6983__A2 _2856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7932__B2 _3723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7932__A1 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4902__I _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8488__A2 _4094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_6_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5171__A1 _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5849__I1 _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_1_clk clknet_4_4_0_clk clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_88_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8412__A2 _4051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5971_ net205 _1522_ _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7710_ _3521_ _3522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4985__A1 _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4922_ reg_file.reg_storage\[4\]\[22\] reg_file.reg_storage\[5\]\[22\] reg_file.reg_storage\[6\]\[22\]
+ reg_file.reg_storage\[7\]\[22\] _0757_ _0837_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8690_ _3688_ _4232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_32_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7641_ reg_file.reg_storage\[5\]\[2\] _3456_ _3458_ _3459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4853_ _0768_ reg_file.reg_storage\[3\]\[20\] _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4784_ _0698_ _0699_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7572_ _0594_ _3034_ _3391_ _3392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_28_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6005__S _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9311_ _0097_ clknet_leaf_17_clk reg_file.reg_storage\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6523_ _2297_ _2364_ _2427_ _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9242_ _0028_ clknet_leaf_103_clk reg_file.reg_storage\[5\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6454_ _2360_ _1978_ _2361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7687__B1 _3495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5162__A1 _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5405_ _0800_ _1320_ _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_9173_ _4511_ _4531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6385_ _2289_ _2290_ _2293_ _2176_ _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_30_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8124_ _3719_ _3812_ _3853_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5336_ _1251_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8954__I _4354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8055_ _3810_ _3811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5267_ _1182_ _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7006_ _2117_ _2893_ _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_126_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5198_ _0672_ _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input27_I inst[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8403__A2 _4038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_50_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6414__A1 _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8957_ _4355_ _4398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7908_ net113 _3698_ _3699_ _3701_ _3703_ _3704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_8888_ _4355_ _4356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7839_ _3036_ _3642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_109_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7914__A1 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7914__B2 _3707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5818__I _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5076__S1 _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4722__I _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9509_ _0295_ clknet_leaf_40_clk reg_file.reg_storage\[11\]\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7390__A2 _3212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4900__A1 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6653__A1 _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6956__A2 _2638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8104__I _3816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5519__I0 reg_file.reg_storage\[12\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5144__A1 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6892__A1 _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6170_ _1997_ _2058_ _2072_ _2083_ _2084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5121_ reg_file.reg_storage\[12\]\[30\] reg_file.reg_storage\[13\]\[30\] reg_file.reg_storage\[14\]\[30\]
+ reg_file.reg_storage\[15\]\[30\] _0758_ _0761_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_110_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8633__A2 _4182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5052_ _0952_ _0913_ _0967_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_79_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8811_ _4309_ _4310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4958__A1 _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8742_ _4191_ _4262_ _4269_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5954_ _1524_ _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8673_ _3648_ _4220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4905_ _0648_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_75_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5885_ _1800_ _1119_ _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7058__C _2120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7624_ _3442_ _3443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4836_ _0747_ _0630_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_90_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7555_ _3372_ _3375_ _3376_ _3377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6175__A3 _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6506_ _2403_ _2406_ _2411_ _2412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4767_ _0654_ net215 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_16_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4698_ _0589_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7486_ _3309_ _3313_ _3314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9225_ _0011_ clknet_leaf_44_clk reg_file.reg_storage\[5\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6437_ _2073_ _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_132_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9156_ _3937_ _4512_ _4521_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6368_ _1771_ _2276_ _2277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_54_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8107_ _3822_ _3844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5319_ _0543_ _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6299_ _2209_ _2210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9087_ reg_file.reg_storage\[4\]\[12\] _3584_ _4465_ _4479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8038_ reg_file.reg_storage\[3\]\[26\] _3799_ _3800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4717__I _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5297__S1 _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4949__A1 _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5548__I _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8863__A2 _4338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6626__A1 _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_106_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5670_ _0792_ _1586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_127_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4621_ _0536_ _0538_ _0540_ _0541_ _0542_ _0543_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_127_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7340_ _3041_ _3179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7271_ _1769_ _1383_ _3116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_9010_ _3957_ _4430_ _4431_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_123_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6865__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _2060_ _2135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5212__S1 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_115_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6153_ _2066_ _2067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6617__A1 _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5104_ _0633_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6084_ _0745_ _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6953__S _2105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5035_ _0850_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7680__I3 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6986_ _1099_ _2856_ _2875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8725_ _4254_ _4257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5937_ _1577_ _1853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8656_ _4208_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7607_ _3424_ _3425_ _3426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input94_I pc[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5868_ _1344_ _1783_ _1784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_134_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5799_ reg_file.reg_storage\[4\]\[14\] reg_file.reg_storage\[5\]\[14\] reg_file.reg_storage\[6\]\[14\]
+ reg_file.reg_storage\[7\]\[14\] _1607_ _1362_ _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_clkbuf_4_14_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4819_ _0734_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8587_ _3987_ _4129_ _4159_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7583__I _3402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9098__A2 _4475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7538_ _3345_ _3346_ _3361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_16_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7469_ _3275_ _3278_ _3297_ _3298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9208_ reg_file.reg_storage\[15\]\[29\] _4546_ _4551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6856__A1 _2725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9139_ _4509_ _4510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7758__I _3566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9022__A2 _4437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7584__A2 _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7707__B net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8836__A2 _4312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5741__I _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4953__S0 _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__I1 reg_file.reg_storage\[9\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9013__A2 _4424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6840_ _0848_ _1853_ _2734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _2664_ _2630_ _2652_ _2665_ _2666_ _2667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_76_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6622__I1 _2523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8510_ _4068_ _4111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5722_ reg_file.reg_storage\[8\]\[19\] reg_file.reg_storage\[9\]\[19\] reg_file.reg_storage\[10\]\[19\]
+ reg_file.reg_storage\[11\]\[19\] _1614_ _0878_ _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5681__S1 _1596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9490_ _0276_ clknet_leaf_85_clk reg_file.reg_storage\[8\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8441_ _4068_ _4069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5653_ _1450_ _1569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5338__A1 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5584_ _1464_ reg_file.reg_storage\[3\]\[29\] _1500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4820__I _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8372_ reg_file.reg_storage\[14\]\[2\] _3926_ _4029_ _4030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4604_ _0521_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7323_ _3157_ net99 _3158_ _3163_ _3164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8827__A2 _4313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7254_ _3050_ _3100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7185_ _3036_ _1901_ _3037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_111_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6747__I _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6205_ _2012_ _1941_ _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ _2037_ _1150_ _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6067_ _1981_ _1982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5813__A2 _1728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5018_ _0933_ _0796_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7015__A1 _2180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5121__S0 _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5577__A1 _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_140_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6969_ _2836_ _2857_ _2858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9688_ _0474_ clknet_leaf_92_clk reg_file.reg_storage\[15\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8708_ reg_file.reg_storage\[8\]\[27\] _4241_ _4245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_62_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7318__A2 _1671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8639_ _4195_ _4182_ _4196_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6829__A1 _1852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_73_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5360__S0 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4905__I _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7006__A1 _2117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5017__B1 _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7557__A2 _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6765__B1 _2661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5032__A3 _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5415__S1 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__A1 _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5179__S0 _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5471__I _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I inst[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8990_ reg_file.reg_storage\[1\]\[6\] _4412_ _4420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7941_ net117 _3728_ _3729_ _3730_ _3732_ _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_77_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7872_ _3263_ _3645_ _3672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9611_ _0397_ clknet_leaf_11_clk reg_file.reg_storage\[1\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5559__A1 _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6823_ _2717_ net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9542_ _0328_ clknet_leaf_45_clk reg_file.reg_storage\[10\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6754_ _1647_ _2650_ _2651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_46_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5705_ _0950_ _1620_ _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6685_ _2139_ _2585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9473_ _0259_ clknet_leaf_126_clk reg_file.reg_storage\[8\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8424_ _3993_ _4018_ _4058_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5636_ _1462_ _1551_ _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8022__I _3769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5567_ _1450_ _1483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5731__A1 _1586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8355_ _1236_ _1106_ _4015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_41_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8286_ _3962_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7306_ net22 _1443_ _3134_ _3148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5498_ _1413_ _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input57_I mem_ld_dat[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7237_ _3078_ _3081_ _3084_ _3085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6287__A2 _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7168_ _3023_ _3024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_129_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_8_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7099_ net6 _2981_ _2982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6119_ _2005_ _2032_ _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4725__I _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7539__A2 _3346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4661__S _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__A2 _2184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8107__I _3822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4635__I _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_2_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6055__C _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__A1 _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5466__I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6470_ _2371_ _1830_ _2372_ _2376_ _2377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_54_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _1336_ _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8140_ reg_file.reg_storage\[6\]\[0\] _3863_ _3864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5352_ _1182_ _1268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_121_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6269__A2 _2180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8071_ reg_file.reg_storage\[2\]\[3\] _3470_ _3822_ _3824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5283_ _0772_ reg_file.reg_storage\[2\]\[10\] _0806_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7022_ _2906_ _2908_ _2909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8966__A1 reg_file.reg_storage\[9\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8973_ _3911_ _4406_ _4408_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7924_ net115 _3698_ _3699_ _3714_ _3717_ _3718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_78_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7855_ _3656_ _3657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8194__A2 _3895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6806_ _2684_ _2676_ _2701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7786_ _3537_ _3592_ _3579_ _3593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9525_ _0311_ clknet_leaf_119_clk reg_file.reg_storage\[11\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4998_ _0823_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_34_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6737_ _2634_ _2384_ _2635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7792__S _3569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9456_ _0242_ clknet_leaf_33_clk reg_file.reg_storage\[12\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6668_ _2561_ _2567_ _1983_ _2568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8407_ _4023_ _4049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5704__A1 _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5619_ _0563_ _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6599_ _2035_ _2500_ _2501_ _2502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9387_ _0173_ clknet_leaf_9_clk reg_file.reg_storage\[14\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8338_ _4000_ _4001_ _4002_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output163_I net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7457__A1 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8269_ _3950_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6432__A2 _2339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6156__B _2018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7766__I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8185__A2 _3882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5243__I0 _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5943__A1 _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7696__A1 _2309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5306__S0 _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5077__I3 _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6423__A2 _1797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5970_ _1877_ _1885_ _1442_ _1886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4921_ _0836_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4852_ _0767_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7640_ _3457_ _3458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_87_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6580__I _1707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6187__A1 _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9125__A1 _4003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4783_ _0614_ _0602_ _0603_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_16_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7571_ _0587_ _0605_ _0707_ _3391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_31_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9310_ _0096_ clknet_leaf_112_clk reg_file.reg_storage\[6\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6522_ _2011_ _2426_ _2427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5537__I1 reg_file.reg_storage\[13\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9241_ _0027_ clknet_leaf_103_clk reg_file.reg_storage\[5\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6453_ _2004_ _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7687__B2 _3500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7687__A1 net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8300__I _3666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9172_ _4530_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5404_ _1313_ _1317_ _1318_ _1319_ _0870_ _0871_ _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8123_ reg_file.reg_storage\[2\]\[26\] _3852_ _3853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6384_ _2248_ _2291_ _2292_ _2293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_2_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8100__A2 _3831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5335_ _1218_ _1249_ _1250_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__4984__B _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8054_ _3753_ _3809_ _3810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5266_ _0978_ _1180_ _1181_ _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_126_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7005_ _2879_ _2706_ _1100_ _2893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8239__I0 reg_file.reg_storage\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4673__A1 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5197_ _0720_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_39_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8956_ _4240_ _4356_ _4397_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8970__I _4405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7907_ _3702_ _3305_ _3497_ _1881_ _3703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_8887_ _4354_ _4355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7838_ _3534_ _3641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7769_ net36 _3411_ _3576_ _3404_ _3577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_53_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9508_ _0294_ clknet_leaf_121_clk reg_file.reg_storage\[11\]\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9439_ _0225_ clknet_leaf_131_clk reg_file.reg_storage\[12\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5770__S _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6169__A1 _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6169__B2 _1947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_95_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5519__I1 reg_file.reg_storage\[13\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5120_ _0765_ _1033_ _1034_ _1035_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6644__A2 _2542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5051_ _0754_ _0966_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_48_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8810_ _3865_ _4178_ _4309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_36_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8741_ reg_file.reg_storage\[11\]\[4\] _4263_ _4269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5953_ _1845_ _1856_ _1868_ _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_48_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8149__A2 _3869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8672_ _4218_ _4214_ _4219_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4904_ reg_file.reg_storage\[8\]\[21\] reg_file.reg_storage\[9\]\[21\] reg_file.reg_storage\[10\]\[21\]
+ reg_file.reg_storage\[11\]\[21\] _0817_ _0818_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_48_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5884_ _1777_ _1800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5907__A1 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7623_ _1981_ _3432_ _3441_ _3442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4835_ net77 _0750_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_106_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7554_ _3372_ _3375_ _3044_ _3376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4766_ _0681_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_133_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6505_ _2057_ _2410_ _2411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4697_ _0612_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7485_ _3292_ _3295_ _3289_ _3310_ _3312_ _3313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9224_ _0010_ clknet_4_10_0_clk reg_file.reg_storage\[5\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6436_ _2343_ _1827_ _2171_ _2344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9155_ reg_file.reg_storage\[15\]\[6\] _4513_ _4521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6367_ _2231_ _2154_ _2232_ _2152_ _2276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_8106_ _3657_ _3837_ _3843_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_54_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5318_ _1120_ _1233_ _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9086_ _4478_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6298_ _0745_ _2209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_4_10_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8037_ _3755_ _3799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5249_ net71 _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA_output126_I net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8388__A2 _4038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7060__A2 _2730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9626__CLK clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5071__A1 _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8939_ _4366_ _4388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4733__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8312__A2 _3975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5757__S0 _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6395__I _2170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6626__A2 _2510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4908__I _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5675__S _1590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9147__S _4516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4620_ _0485_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6562__A1 _2180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8303__A2 _3971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5474__I _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7270_ _3112_ _3114_ _3115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_13_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6314__A1 _2046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6865__A2 _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6221_ _1800_ _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_122_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6152_ _1789_ _0719_ _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5103_ _0954_ _1016_ _1017_ _1018_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5676__I0 reg_file.reg_storage\[1\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6083_ _1907_ _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4818__I _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7814__A1 _3205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5034_ _0949_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_79_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6985_ _2872_ _2373_ _2873_ _2874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6254__B _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8724_ _4255_ _4256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _0849_ _1852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8655_ reg_file.reg_storage\[8\]\[11\] _4207_ _4198_ _4208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7606_ _0880_ _3390_ _3394_ _3425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_63_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ net24 _0717_ _0703_ _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_134_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5798_ reg_file.reg_storage\[12\]\[14\] reg_file.reg_storage\[13\]\[14\] reg_file.reg_storage\[14\]\[14\]
+ reg_file.reg_storage\[15\]\[14\] _1607_ _1609_ _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5600__I0 reg_file.reg_storage\[12\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8586_ reg_file.reg_storage\[12\]\[23\] _4127_ _4159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4818_ _0668_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input87_I pc[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4749_ _0596_ _0598_ _0610_ _0664_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__5384__I net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7537_ _1498_ _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6305__A1 _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7468_ _3270_ _3287_ _3297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9207_ _4003_ _4548_ _4550_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_116_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6419_ _2261_ _0981_ _2326_ _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_116_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7399_ net72 _3211_ _3227_ _3234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9138_ _3761_ _4021_ _4509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4728__I _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9069_ reg_file.reg_storage\[4\]\[4\] _4463_ _4469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7281__A2 _3116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5044__A1 _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6164__B _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8781__A2 _4288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6792__A1 _2684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5347__A2 _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4953__S1 _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7272__A2 _3102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7949__I _3739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__A1 _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8221__A1 _3388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6770_ _2644_ _2651_ _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5721_ _0626_ _1582_ _1583_ _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_18_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8440_ _4067_ _4068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7878__A4 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5652_ _1437_ _1380_ _1412_ _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5583_ reg_file.reg_storage\[4\]\[29\] reg_file.reg_storage\[5\]\[29\] reg_file.reg_storage\[6\]\[29\]
+ reg_file.reg_storage\[7\]\[29\] _1482_ _1489_ _1499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8371_ _4028_ _4029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4603_ _0524_ _0526_ _0509_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_142_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7322_ _3160_ _3162_ _3163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4641__S0 _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6838__A2 _2525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7253_ _3097_ _3098_ _3099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_7184_ _2975_ _3036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_111_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ _2008_ _2117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _2034_ _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_99_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6066_ _0733_ _1906_ _1980_ _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5017_ _0911_ _0913_ _0835_ _0932_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8212__A1 _3734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5121__S1 _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8707_ _4173_ _4244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6968_ _2834_ _2484_ _2857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6774__A1 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7594__I _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9687_ _0473_ clknet_leaf_92_clk reg_file.reg_storage\[15\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6899_ _2362_ _2790_ _2791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5919_ _1667_ _1835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7869__A4 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8638_ reg_file.reg_storage\[8\]\[6\] _4183_ _4196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8569_ _4149_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_134_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6673__I _1580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5265__A1 _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5360__S1 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5017__A1 _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8754__A2 _4262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5017__B2 _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6765__A1 _2404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6517__A1 _2113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4921__I _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_143_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5179__S1 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9160__S _4522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6048__A3 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7245__A2 _3081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7940_ _3715_ _3357_ _3731_ _3732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_89_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7871_ _3485_ _3671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_77_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6822_ _1984_ _2703_ _2716_ _2717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9610_ _0396_ clknet_4_0_0_clk reg_file.reg_storage\[1\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8745__A2 _4263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5199__I _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9541_ _0327_ clknet_leaf_40_clk reg_file.reg_storage\[10\]\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6753_ _2565_ _2627_ _2649_ _2650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5927__I _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5704_ _0735_ _1603_ _1619_ _1620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6684_ _2261_ _2339_ _2584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9472_ _0258_ clknet_leaf_127_clk reg_file.reg_storage\[8\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8423_ reg_file.reg_storage\[14\]\[25\] _4019_ _4058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5635_ _1545_ _1548_ _1549_ _1550_ _1534_ _1537_ _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_61_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8354_ _4013_ _3916_ _4014_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5566_ _1369_ _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_115_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5731__A2 _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8285_ reg_file.reg_storage\[7\]\[15\] _3961_ _3927_ _3962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7305_ _3134_ net22 _3138_ _3147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_13_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5497_ _1352_ _1412_ _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_113_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7236_ _3082_ _3072_ _3083_ _3084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7167_ _3022_ _3023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_129_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_129_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7098_ _2969_ _2972_ _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6118_ _2029_ _1230_ _2031_ _2032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_142_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6049_ _1962_ _1963_ _1964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_1_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__S0 _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7475__A2 _3294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5238__A1 _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6986__A1 _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6109__S _2022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__A2 _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9152__A2 _4512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7163__A1 net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7163__B2 _1717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7962__I _3750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6910__A1 _2797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5420_ _1335_ _0831_ _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5351_ _1252_ _1253_ _1266_ _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5282_ _1061_ reg_file.reg_storage\[3\]\[10\] _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8070_ _3823_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7021_ _1508_ _2907_ _2908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8972_ reg_file.reg_storage\[1\]\[0\] _4407_ _4408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6977__A1 _2030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7923_ _3715_ _3328_ _3716_ _3717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7854_ net106 _3601_ _3653_ _3655_ _3656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_136_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7785_ _3588_ _3405_ _3407_ _3591_ _3592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_6805_ _2697_ _2699_ _2700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_19_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6736_ _2214_ _2634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9524_ _0310_ clknet_leaf_24_clk reg_file.reg_storage\[11\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _0912_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_34_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9143__A2 _4513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7154__A1 _1457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7154__B2 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9455_ _0241_ clknet_leaf_55_clk reg_file.reg_storage\[12\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6667_ _1580_ _2566_ _2567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9065__S _4466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8406_ _3967_ _4044_ _4048_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5618_ _1533_ _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5704__A2 _1603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6901__A1 _2137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6598_ _2018_ _2426_ _2501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9386_ _0172_ clknet_leaf_8_clk reg_file.reg_storage\[14\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8337_ reg_file.reg_storage\[7\]\[27\] _3997_ _4002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5549_ _1450_ _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7457__A2 _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5012__S0 _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8268_ reg_file.reg_storage\[7\]\[10\] _3949_ _3941_ _3950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_57_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output156_I net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8199_ reg_file.reg_storage\[6\]\[23\] _3868_ _3900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7219_ _3066_ _3067_ _3068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_70_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A1 _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6951__I _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5943__A2 _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7782__I net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7696__A2 _3504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5459__A1 _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4646__I _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8948__A2 _4361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5306__S1 _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6959__A1 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4920_ _0641_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4851_ _0756_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_136_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9125__A2 _4498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7570_ net30 _3390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4782_ _0597_ _0599_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_7_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6521_ _1962_ _2425_ _2426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_15_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8884__A1 reg_file.reg_storage\[10\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9240_ _0026_ clknet_leaf_104_clk reg_file.reg_storage\[5\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6302__S _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6452_ _1934_ _2328_ _2358_ _2284_ _2359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_43_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5242__S0 _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9171_ reg_file.reg_storage\[15\]\[13\] _3597_ _4515_ _4530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5403_ reg_file.reg_storage\[8\]\[3\] reg_file.reg_storage\[9\]\[3\] reg_file.reg_storage\[10\]\[3\]
+ reg_file.reg_storage\[11\]\[3\] _1122_ _0867_ _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8122_ _3810_ _3852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6383_ _2079_ _2129_ _2292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5334_ net94 _0748_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8053_ _3808_ _3809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6111__A2 _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5265_ _0490_ net218 _0715_ _0692_ _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7004_ _2061_ _2692_ _2892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5196_ _0981_ _1104_ _1111_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_126_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4673__A2 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8955_ reg_file.reg_storage\[9\]\[26\] _4396_ _4397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8886_ _3397_ _4171_ _4354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_129_clk clknet_4_5_0_clk clknet_leaf_129_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7906_ _3484_ _3702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7837_ _3631_ _3640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7375__A1 _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7768_ _3575_ _3406_ _3576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9116__A2 _4457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7127__A1 _1729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6719_ _2616_ _1858_ _2617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7699_ reg_file.reg_storage\[5\]\[7\] _3511_ _3492_ _3512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7816__B _3620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9507_ _0293_ clknet_leaf_135_clk reg_file.reg_storage\[11\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9438_ _0224_ clknet_leaf_87_clk reg_file.reg_storage\[12\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9369_ _0155_ clknet_leaf_97_clk reg_file.reg_storage\[7\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__S1 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__I _1765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__A1 _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7777__I _3584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_141_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9107__A2 _4488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7118__A1 _1664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5519__I2 reg_file.reg_storage\[14\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5050_ _0953_ _0960_ _0962_ _0963_ _0965_ _0929_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__9043__A1 _4003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7054__B1 _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5952_ _1857_ _1867_ _1579_ _1868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8740_ _4268_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4903_ reg_file.reg_storage\[12\]\[21\] reg_file.reg_storage\[13\]\[21\] reg_file.reg_storage\[14\]\[21\]
+ reg_file.reg_storage\[15\]\[21\] _0817_ _0818_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_62_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8671_ reg_file.reg_storage\[8\]\[16\] _4203_ _4219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5883_ _1796_ _1757_ _1797_ _1798_ _1799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_75_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7622_ _3436_ _3440_ _3441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4834_ _0749_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7553_ _3373_ _3363_ _3374_ _3375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4765_ _0663_ _0662_ _0593_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__4966__I0 _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6504_ _2015_ _2407_ _2408_ _2409_ _2410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_44_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9223_ _0009_ clknet_leaf_30_clk reg_file.reg_storage\[5\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4696_ _0609_ _0587_ _0601_ _0611_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7484_ _3311_ _3312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_113_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6435_ _1734_ _2343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_132_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9154_ _4520_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6366_ _2275_ net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_9085_ reg_file.reg_storage\[4\]\[11\] _3567_ _4472_ _4478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8105_ reg_file.reg_storage\[2\]\[18\] _3842_ _3843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8085__A2 _3831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5317_ _1179_ _1232_ _1103_ _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8036_ _3710_ _3757_ _3798_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6297_ _2205_ _2207_ _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5694__I1 reg_file.reg_storage\[9\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ _1162_ _1163_ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input32_I inst[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5438__A4 _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7832__A2 _3212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5179_ reg_file.reg_storage\[8\]\[27\] reg_file.reg_storage\[9\]\[27\] reg_file.reg_storage\[10\]\[27\]
+ reg_file.reg_storage\[11\]\[27\] _0855_ _0857_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__8981__I _4414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6399__A2 _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output119_I net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8938_ _4222_ _4381_ _4387_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8869_ _4236_ _4306_ _4344_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5454__S0 _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6571__A2 _2269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5757__S1 _1672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5781__S _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6676__I _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6625__B _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8000__A2 _3778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6562__A2 _2463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7511__A1 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6314__A2 _2224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ _2000_ _2115_ _2132_ _2057_ _2133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_40_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6151_ _0745_ _2065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5102_ _0957_ reg_file.reg_storage\[2\]\[31\] _0958_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6078__A1 _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6082_ _1991_ _1995_ _1996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_29_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5033_ _0936_ _0937_ _0948_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_79_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7578__A1 _3388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6984_ _2872_ _2077_ _2873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6250__A1 _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8723_ _4254_ _4255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5935_ _1847_ _1848_ _1543_ _1850_ _1851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8654_ _3566_ _4207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _1524_ _1651_ _1781_ _1782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8242__S _3928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_60_clk clknet_4_11_0_clk clknet_leaf_60_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7605_ _0975_ _1106_ _3424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_63_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6002__A1 _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _0720_ _0726_ _0732_ _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_35_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5797_ reg_file.reg_storage\[1\]\[14\] _1712_ _1362_ _1713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5600__I1 reg_file.reg_storage\[13\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8585_ _3984_ _4154_ _4158_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_134_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4748_ net26 _0589_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_7_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7536_ net86 _3359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6305__A2 _2215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4679_ net28 _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7467_ _3292_ _3295_ _3296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9206_ reg_file.reg_storage\[15\]\[28\] _4546_ _4550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6418_ _2209_ _2326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9137_ _3911_ _4506_ _4508_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_116_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8058__A2 _3813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7398_ net72 net73 _3211_ _3233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6349_ _2258_ _2259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_47_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5816__A1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9068_ _4468_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_94_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8019_ _3763_ _3789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8152__S _3873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_51_clk clknet_4_10_0_clk clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_32_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7790__I _3596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5122__I3 reg_file.reg_storage\[11\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_105_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8221__A2 _3754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9158__S _4522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5720_ _1632_ _1634_ _0908_ _1636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_58_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_42_clk clknet_4_8_0_clk clknet_leaf_42_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7186__B _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5651_ _0791_ _1566_ _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5485__I _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8370_ _4022_ _4028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4602_ reg_file.reg_storage\[1\]\[2\] _0525_ _0499_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5582_ _1497_ _1480_ _1413_ _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_131_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7321_ net67 _3161_ _3162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7252_ _1270_ _3088_ _3098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6203_ _2060_ _2116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7183_ _0663_ _3034_ _3035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_51_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _0935_ _1177_ _2047_ _2048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6065_ _1907_ _1970_ _1976_ _1979_ _1980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5016_ _0914_ _0925_ _0931_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5657__S0 _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6223__A1 _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6967_ _1441_ _2856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8706_ _3725_ _4243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6774__A2 _1564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5918_ _1683_ _1831_ _1833_ _1834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_24_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9686_ _0472_ clknet_leaf_86_clk reg_file.reg_storage\[15\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33_clk clknet_4_8_0_clk clknet_leaf_33_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6898_ _2029_ _2728_ _2789_ _2790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5409__S0 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8637_ _3501_ _4195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5849_ net160 _0741_ _0680_ _1765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_118_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8568_ reg_file.reg_storage\[12\]\[15\] _3961_ _4131_ _4149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output186_I net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7519_ _3226_ _3340_ _3342_ _3324_ _3343_ net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_32_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8499_ reg_file.reg_storage\[13\]\[22\] _4074_ _4105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_55_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6462__A1 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8451__A2 _4075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7986__S _3769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5017__A2 _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__A1 _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_24_clk clknet_4_1_0_clk clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_137_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__S0 _1605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7870_ _3640_ _3669_ _3652_ _3670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_54_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _2213_ _2571_ _2712_ _2641_ _2715_ _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_49_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7402__B1 _3235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6756__A2 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9540_ _0326_ clknet_leaf_121_clk reg_file.reg_storage\[10\]\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7953__A1 _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6752_ _1620_ _2439_ _2649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_15_clk clknet_4_0_0_clk clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6683_ _2582_ _2583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5703_ _1604_ _1586_ _1618_ _1619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_57_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9471_ _0257_ clknet_leaf_120_clk reg_file.reg_storage\[8\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8422_ _3990_ _4018_ _4057_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5634_ reg_file.reg_storage\[4\]\[23\] reg_file.reg_storage\[5\]\[23\] reg_file.reg_storage\[6\]\[23\]
+ reg_file.reg_storage\[7\]\[23\] _1471_ _1483_ _1550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_6_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8353_ reg_file.reg_storage\[7\]\[31\] _3914_ _4014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5811__S0 _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7304_ _3145_ _3133_ _3146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5565_ _0722_ _1480_ _1413_ _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_8284_ _3622_ _3961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5496_ _1411_ _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_113_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7235_ _3067_ _3069_ _3083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7166_ _3021_ _3022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_129_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6117_ _2030_ _1267_ _2031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7097_ net108 _2974_ _2980_ net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_142_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _1121_ _1130_ _0909_ _1963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_29_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output101_I net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7999_ _3763_ _3778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_138_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9669_ _0455_ clknet_leaf_39_clk reg_file.reg_storage\[15\]\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5853__I net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8121__A1 _3710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8672__A2 _4214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6986__A2 _2856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5797__I0 reg_file.reg_storage\[1\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8360__A1 reg_file.reg_storage\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xload_slew1 _2413_ net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_55_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6910__A2 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5350_ _1265_ _0910_ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5281_ reg_file.reg_storage\[1\]\[10\] _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7020_ _1521_ _2537_ _2881_ _2907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9171__S _4515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_4_clk clknet_4_4_0_clk clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8415__A2 _4049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8971_ _4404_ _4407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5229__A2 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7922_ _1356_ _3403_ _3716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5003__I _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7853_ _3607_ _3237_ _3634_ _3654_ _3655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_7784_ net37 _3411_ _3590_ _3404_ _3591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_6804_ _1848_ _2698_ _2699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4842__I _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4996_ _0620_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9523_ _0309_ clknet_leaf_76_clk reg_file.reg_storage\[11\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6735_ _1997_ _2632_ _2633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5401__A2 _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9454_ _0240_ clknet_leaf_57_clk reg_file.reg_storage\[12\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6666_ _2562_ _2565_ _2566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8405_ reg_file.reg_storage\[14\]\[17\] _4038_ _4048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9385_ _0171_ clknet_leaf_50_clk reg_file.reg_storage\[14\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6901__A2 _2588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5617_ _1532_ _1533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6597_ _2494_ _2142_ _1963_ _2500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_33_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8336_ _3914_ _4001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5548_ _1463_ _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4912__A1 _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input62_I mem_ld_dat[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8267_ _3555_ _3949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5012__S1 _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5479_ _1105_ _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6665__A1 _1707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7218_ net90 _3067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8198_ _3689_ _3895_ _3899_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output149_I net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8406__A2 _4044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7149_ net162 _2979_ _3015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7090__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8224__I _3913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8590__A1 reg_file.reg_storage\[12\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5243__I2 _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5156__A1 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8894__I _4360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6656__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5459__A2 _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7303__I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9070__A2 _4462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5631__A2 reg_file.reg_storage\[2\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7908__A1 net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__B _2272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4850_ reg_file.reg_storage\[1\]\[20\] _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7908__B2 _3701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7973__I _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6520_ _2387_ _2335_ _2425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _0677_ _0696_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_31_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8333__A1 _3996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5493__I _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6451_ _1967_ _1920_ _2137_ _2358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5242__S1 _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6382_ _2246_ _2119_ _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9170_ _4529_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5402_ reg_file.reg_storage\[12\]\[3\] reg_file.reg_storage\[13\]\[3\] reg_file.reg_storage\[14\]\[3\]
+ reg_file.reg_storage\[15\]\[3\] _1122_ _1123_ _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_140_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8121_ _3710_ _3812_ _3851_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5333_ _1248_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_100_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8052_ _3389_ _3807_ _3394_ _3808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_10_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5264_ _0882_ _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7003_ _2885_ _2890_ _2891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5195_ _1110_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_126_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9061__A2 _4463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8954_ _4354_ _4396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7905_ _2978_ _3519_ _3700_ _3701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_108_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8885_ _4252_ _4307_ _4353_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7836_ _3600_ _3638_ _3639_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4572__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7767_ net45 _3575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4979_ reg_file.reg_storage\[1\]\[17\] _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_108_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9076__S _4472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8324__A1 _3990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6718_ _0949_ _2616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7698_ _3510_ _3511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9506_ _0292_ clknet_leaf_121_clk reg_file.reg_storage\[11\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9437_ _0223_ clknet_leaf_88_clk reg_file.reg_storage\[13\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6649_ _2301_ _2549_ _2332_ _2550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9368_ _0154_ clknet_leaf_95_clk reg_file.reg_storage\[7\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9299_ _0085_ clknet_leaf_25_clk reg_file.reg_storage\[2\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8319_ reg_file.reg_storage\[7\]\[23\] _3922_ _3988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8219__I _3420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5310__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__A2 _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7063__A1 _2254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7366__A2 _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8889__I _4354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8866__A2 _4311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6877__A1 _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4657__I _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5951_ _1859_ _1866_ _1649_ _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5604__A2 _1519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8670_ _3637_ _4218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4902_ _0635_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7357__A2 _3184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5882_ _1310_ _0979_ _1798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_117_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4833_ _0748_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7621_ net76 _3401_ _1180_ _3439_ _3417_ _3440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_29_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7636__C _3453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7552_ _3359_ _3360_ _3374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4764_ _0679_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_132_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ _2027_ _2023_ _2065_ _2409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7483_ _3292_ _3295_ _3299_ _3284_ _3311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_9222_ _0008_ clknet_leaf_41_clk reg_file.reg_storage\[5\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6434_ _2192_ _2342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4695_ _0610_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7208__I net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9153_ reg_file.reg_storage\[15\]\[5\] _3490_ _4516_ _4520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6365_ _2087_ _2244_ _2274_ _2275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9084_ _4477_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8104_ _3816_ _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_54_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6296_ _2161_ _2206_ _2207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5316_ _1183_ _1206_ _1231_ _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8035_ reg_file.reg_storage\[3\]\[25\] _3758_ _3798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4567__I _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5247_ _0795_ _1163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5843__A2 _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5178_ reg_file.reg_storage\[12\]\[27\] reg_file.reg_storage\[13\]\[27\] reg_file.reg_storage\[14\]\[27\]
+ reg_file.reg_storage\[15\]\[27\] _0866_ _0857_ _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_input25_I inst[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8937_ reg_file.reg_storage\[9\]\[18\] _4386_ _4387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5151__S0 _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8868_ reg_file.reg_storage\[10\]\[24\] _4307_ _4344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8799_ _4248_ _4298_ _4301_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7819_ _3623_ _3624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_65_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5454__S1 _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7284__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9025__A2 _4435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_6_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5390__S0 _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5598__A1 _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7339__A2 _3167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4940__I _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4956__S0 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6150_ _2063_ _2064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5101_ _0892_ reg_file.reg_storage\[3\]\[31\] _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7275__B2 _3119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6081_ _1992_ _1993_ _1994_ _1995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__9016__A2 _4430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5032_ _0912_ _0938_ _0947_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5720__B _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7578__A2 _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _1099_ _2856_ _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8527__A1 reg_file.reg_storage\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8722_ _3754_ _4171_ _4254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5934_ _1849_ _1566_ _1850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6107__I _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8653_ _4206_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5865_ _1756_ _1780_ _1781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8322__I _3989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7604_ _3400_ _3421_ _3423_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4816_ _0704_ _0731_ _0724_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_113_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5796_ reg_file.reg_storage\[2\]\[14\] reg_file.reg_storage\[3\]\[14\] _1611_ _1712_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8584_ reg_file.reg_storage\[12\]\[22\] _4127_ _4158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5061__I0 _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7535_ _3045_ _3355_ _3357_ _3324_ _3358_ net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_4747_ _0607_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_4678_ _0595_ net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7466_ _1553_ _3295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9205_ _3999_ _4548_ _4549_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6417_ _2324_ _1233_ _2325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7397_ _3229_ _3231_ _3232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9136_ reg_file.reg_storage\[15\]\[0\] _4507_ _4508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_116_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6348_ _0704_ _0719_ _2258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8992__I _4414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6279_ _2176_ _2182_ _2190_ _2191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9067_ reg_file.reg_storage\[4\]\[3\] _3469_ _4466_ _4468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6313__I0 _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8018_ _3649_ _3784_ _3788_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_99_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5372__S0 _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9191__A1 _3980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8232__I _3922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8541__I1 _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7257__A1 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8407__I _4023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7009__A1 _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8509__A1 _3996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7980__A2 _3766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__A1 _1902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5650_ _1417_ _1557_ _1565_ _1566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_72_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__I net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4601_ reg_file.reg_storage\[2\]\[2\] reg_file.reg_storage\[3\]\[2\] _0502_ _0525_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5581_ net22 _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_142_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7914__C _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7320_ _1656_ _3161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_40_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4929__S0 _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7251_ net93 _3097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ _2102_ _2113_ _2114_ _2115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7182_ _0746_ _3034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5006__I _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6133_ _2006_ _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6064_ _1791_ _1978_ _1979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4845__I _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5015_ _0927_ _0930_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6471__A2 _2370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6966_ _2855_ net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__6223__A2 _2135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_140_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8705_ _4240_ _4174_ _4242_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5917_ _1669_ _1832_ _1833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_124_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9685_ _0471_ clknet_leaf_23_clk reg_file.reg_storage\[15\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6897_ _2012_ _2788_ _2789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5409__S1 _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input92_I pc[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8636_ _4194_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5848_ _1280_ _1763_ _1764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8567_ _3958_ _4147_ _4148_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_118_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5779_ _1588_ _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5734__A1 _1635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7518_ _3051_ net116 _3343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8498_ _3981_ _4101_ _4104_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_2_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output179_I net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7449_ _3279_ _3270_ _3280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9119_ reg_file.reg_storage\[4\]\[26\] _4496_ _4497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6462__A2 _2368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4755__I _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8227__I _3442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8163__S _3879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9164__A1 _3945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9058__I _4460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5820__S1 _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_140_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5027__S _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5697__S _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6820_ _2697_ _1542_ _2372_ _2714_ _2715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__9169__S _4515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7953__A2 _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6751_ _2644_ net240 _2574_ _2647_ _2648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__5964__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5702_ _1610_ _1613_ _1616_ _1617_ _1533_ _1536_ _1618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_9470_ _0256_ clknet_leaf_109_clk reg_file.reg_storage\[8\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6682_ _2066_ _2582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8421_ reg_file.reg_storage\[14\]\[24\] _4019_ _4057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5716__A1 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ reg_file.reg_storage\[12\]\[23\] reg_file.reg_storage\[13\]\[23\] reg_file.reg_storage\[14\]\[23\]
+ reg_file.reg_storage\[15\]\[23\] _1471_ _1483_ _1549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_45_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8352_ _4012_ _4013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5811__S1 _1672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5564_ _1479_ _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_115_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7303_ net66 _3145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8283_ _3958_ _3959_ _3960_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5495_ _0728_ _0682_ _0683_ _1410_ _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__5575__S0 _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7234_ net90 _3069_ _3082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7165_ _2970_ _1981_ _3021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5495__A3 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6116_ _2007_ _2030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7096_ _2979_ _2980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_129_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_31_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__S0 _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6047_ _1193_ _0909_ _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_29_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_46_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8197__A2 _3868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7944__A2 _3734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7998_ _3777_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_138_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6949_ _2833_ _2838_ _2839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_37_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9668_ _0454_ clknet_leaf_16_clk reg_file.reg_storage\[15\]\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8619_ _4181_ _4182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_134_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_104_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9599_ _0385_ clknet_4_7_0_clk reg_file.reg_storage\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8121__A2 _3812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_119_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8158__S _3873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7997__S _3775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8188__A2 _3893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6199__A1 _2110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7935__A2 _3726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5797__I1 _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9137__A1 _3911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6371__A1 _1938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8112__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5280_ reg_file.reg_storage\[4\]\[10\] reg_file.reg_storage\[5\]\[10\] reg_file.reg_storage\[6\]\[10\]
+ reg_file.reg_storage\[7\]\[10\] _0839_ _0902_ _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5557__S0 _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_74_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8970_ _4405_ _4406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7623__A1 _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7921_ _3047_ _3715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8179__A2 _3882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7852_ _3255_ _3645_ _3654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7783_ _3589_ _3406_ _3590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6803_ _2671_ _2674_ _2672_ _2698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4995_ net72 _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_19_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9522_ _0308_ clknet_leaf_67_clk reg_file.reg_storage\[11\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6734_ _2625_ _2630_ _2632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_34_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_9453_ _0239_ clknet_leaf_12_clk reg_file.reg_storage\[12\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8330__I _3995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8404_ _3964_ _4044_ _4047_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6665_ _1707_ _2486_ _2563_ _2564_ _2565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_45_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9384_ _0170_ clknet_leaf_48_clk reg_file.reg_storage\[14\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer28_I _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6596_ _2494_ _2483_ _2266_ _2498_ _2499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__6362__A1 _1938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5616_ _1531_ _1532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_42_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8335_ _3999_ _4000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5547_ _1390_ _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_112_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5478_ reg_file.reg_storage\[8\]\[25\] reg_file.reg_storage\[9\]\[25\] reg_file.reg_storage\[10\]\[25\]
+ reg_file.reg_storage\[11\]\[25\] _1387_ _1388_ _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_8266_ _3946_ _3923_ _3948_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input55_I mem_ld_dat[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6665__A2 _2486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7217_ _1300_ _3066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_111_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_92_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8197_ reg_file.reg_storage\[6\]\[22\] _3868_ _3899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7148_ _3006_ _1575_ _3014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6417__A2 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7079_ _2961_ _2169_ _2542_ _2682_ _2962_ _2963_ _2964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_68_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7917__A2 _3710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5243__I3 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__A2 _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5305__S _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5104__I _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7605__A1 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5092__A1 _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__C _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8581__A2 _4154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4780_ _0678_ _0695_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_129_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6592__A1 _2494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__A2 _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8333__A2 _3915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6344__A1 _2110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ _2355_ _2356_ _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_125_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6381_ _2128_ _2100_ _2003_ _2290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5401_ _1314_ _0775_ _1315_ _1316_ _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8097__A1 _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8120_ reg_file.reg_storage\[2\]\[25\] _3813_ _3851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5332_ _1243_ _1245_ _1246_ _1247_ _0648_ _0649_ _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_11_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8051_ net30 _3807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _1150_ _1177_ _1178_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7002_ _2832_ net235 _2887_ _2888_ _2889_ _2786_ _2890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5194_ _1109_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_126_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5702__S0 _1533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8953_ _4238_ _4356_ _4395_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7904_ _3631_ _3700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_108_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8884_ reg_file.reg_storage\[10\]\[31\] _4305_ _4353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5473__I3 reg_file.reg_storage\[7\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7835_ reg_file.reg_storage\[5\]\[16\] _3544_ _3639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8572__A2 _4141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7766_ net53 _3574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_4978_ reg_file.reg_storage\[4\]\[17\] reg_file.reg_storage\[5\]\[17\] reg_file.reg_storage\[6\]\[17\]
+ reg_file.reg_storage\[7\]\[17\] _0892_ _0893_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_47_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9505_ _0291_ clknet_leaf_127_clk reg_file.reg_storage\[11\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_137_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8324__A2 _3915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7697_ _3509_ _3510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6717_ _2025_ _2571_ _2615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9436_ _0222_ clknet_leaf_90_clk reg_file.reg_storage\[13\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6648_ _2428_ _2548_ _2185_ _2549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9367_ _0153_ clknet_leaf_91_clk reg_file.reg_storage\[7\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8318_ _3986_ _3987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6579_ _1820_ _2482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output161_I net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9298_ _0084_ clknet_leaf_67_clk reg_file.reg_storage\[2\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8249_ reg_file.reg_storage\[7\]\[5\] _3935_ _3928_ _3936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6810__A2 _2503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8012__A1 _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6574__A1 _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8315__A2 _3922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4938__I _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8145__I _3867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5950_ _1864_ _1865_ _1621_ _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4901_ _0801_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_87_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5881_ _0885_ _0677_ _1797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7620_ _3438_ _3439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4832_ _0747_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7551_ _3359_ _3360_ _3373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4763_ _0666_ _0667_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_126_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6502_ _2114_ _2053_ _2408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6317__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4694_ net12 net1 net23 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7482_ _3286_ _3296_ _3310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9221_ _0007_ clknet_leaf_38_clk reg_file.reg_storage\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6433_ _2289_ _2331_ _2340_ _2341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_132_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6364_ _2260_ _2273_ _2274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9152_ _3932_ _4512_ _4519_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8103_ _3649_ _3837_ _3841_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9083_ reg_file.reg_storage\[4\]\[10\] _3556_ _4472_ _4477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4848__I _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6295_ _2164_ _2206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5315_ _1183_ _1230_ _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8034_ _3705_ _3757_ _3797_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5246_ _1161_ _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5177_ _0899_ _1090_ _1091_ _1092_ _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5679__I _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5056__A1 _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8936_ _4360_ _4386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input18_I inst[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5151__S1 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4803__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8867_ _4234_ _4313_ _4343_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9087__S _4465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8798_ reg_file.reg_storage\[11\]\[29\] _4296_ _4301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7818_ _3622_ _3623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_65_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7749_ _3558_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6308__A1 _2217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9419_ _0205_ clknet_leaf_2_clk reg_file.reg_storage\[13\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7808__A1 net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4590__I0 reg_file.reg_storage\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7284__A2 _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8784__A2 _4261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8536__A2 _4128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4653__S0 _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4956__S1 _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4581__I0 reg_file.reg_storage\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4668__I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5100_ reg_file.reg_storage\[1\]\[31\] _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7275__A2 net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6080_ _1309_ _1989_ _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5031_ _0939_ _0943_ _0944_ _0945_ _0785_ _0946_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_73_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8721_ _4252_ _4175_ _4253_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _2421_ _2431_ _2870_ _2582_ _2871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_105_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5933_ _0791_ _1849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8652_ reg_file.reg_storage\[8\]\[10\] _4205_ _4198_ _4206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5864_ _1757_ _1775_ _1776_ _1779_ _1780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_8583_ _3981_ _4154_ _4157_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7603_ reg_file.reg_storage\[5\]\[0\] _3422_ _3423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4815_ _0730_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5795_ reg_file.reg_storage\[8\]\[14\] reg_file.reg_storage\[9\]\[14\] reg_file.reg_storage\[10\]\[14\]
+ reg_file.reg_storage\[11\]\[14\] _1607_ _1362_ _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_113_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7534_ _3051_ net117 _3358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6123__I _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4746_ _0588_ _0586_ _0601_ net230 _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_0_102_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4677_ _0594_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_43_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7465_ _3292_ _3293_ _3294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_32_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9204_ reg_file.reg_storage\[15\]\[27\] _4546_ _4549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6416_ _2139_ _2324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7396_ _3213_ _3223_ _3230_ _3231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9135_ _4504_ _4507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_116_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6347_ _1787_ _2257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7266__A2 _3099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _2177_ _2184_ _2188_ _2189_ _2190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_9066_ _4467_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8017_ reg_file.reg_storage\[3\]\[17\] _3778_ _3788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5229_ _0890_ _1144_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5372__S1 _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output124_I net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8919_ reg_file.reg_storage\[9\]\[10\] _4205_ _4372_ _4377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6529__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9191__A2 _4538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5201__A1 net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7257__A2 _3102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6208__I _2097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4951__I _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4600_ reg_file.reg_storage\[4\]\[2\] reg_file.reg_storage\[5\]\[2\] reg_file.reg_storage\[6\]\[2\]
+ reg_file.reg_storage\[7\]\[2\] _0513_ _0514_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_26_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5580_ _1495_ _1041_ _1496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7250_ _3077_ _3089_ _3096_ net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4929__S1 _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6201_ _2044_ _2114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_68_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7181_ _2984_ _3030_ _2971_ net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8445__A1 _3425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5259__A1 _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6132_ _2045_ _2046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7248__A2 _3090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6063_ _1977_ _1902_ _1946_ _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5014_ _0906_ _0928_ _0929_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6965_ _2839_ _2840_ _2848_ _2854_ _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__7658__B _3472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8704_ reg_file.reg_storage\[8\]\[26\] _4241_ _4242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9684_ _0470_ clknet_leaf_26_clk reg_file.reg_storage\[15\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5916_ _1682_ _1832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_119_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6896_ _2742_ _2706_ _1059_ _2788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8635_ reg_file.reg_storage\[8\]\[5\] _4193_ _4187_ _4194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_24_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5847_ _1382_ _0792_ _1354_ _1762_ _1763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_134_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8566_ reg_file.reg_storage\[12\]\[14\] _4141_ _4148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_118_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5734__A2 _1636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6931__A1 _2137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5778_ _1131_ _1693_ _1694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input85_I pc[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8497_ reg_file.reg_storage\[13\]\[21\] _4099_ _4104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4729_ _0634_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_17_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7517_ net84 _3341_ _3342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA_clkbuf_leaf_5_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110_clk clknet_4_13_0_clk clknet_leaf_110_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7448_ _3260_ _3263_ _3279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7379_ _3197_ _3206_ _3215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9118_ _4454_ _4496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7239__A2 _3080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9049_ _4012_ _4407_ _4453_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8987__A2 _4411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5345__S1 _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_103_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4771__I _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5422__A1 _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9164__A2 _4512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A2 _1511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7175__A1 _2972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_101_clk clknet_4_15_0_clk clknet_leaf_101_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7478__A2 net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_112_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8427__A1 _3996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8978__A2 _4412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6139__S _2052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5661__A1 _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ _2645_ _2577_ _2646_ _2647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4681__I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5701_ reg_file.reg_storage\[4\]\[18\] reg_file.reg_storage\[5\]\[18\] reg_file.reg_storage\[6\]\[18\]
+ reg_file.reg_storage\[7\]\[18\] _1615_ _1609_ _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__9155__A2 _4513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6681_ _2573_ _2562_ _2574_ _2580_ _2581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_46_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5716__A2 _1631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6913__A1 _2725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5632_ _1427_ _0859_ _1546_ _1547_ _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_rebuffer8_I net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8420_ _3987_ _4026_ _4056_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5272__S0 _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8351_ _3750_ _4012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ _1411_ _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_130_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6401__I _2309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7302_ _3075_ _3144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8282_ reg_file.reg_storage\[7\]\[14\] _3947_ _3960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5494_ _0608_ _0746_ _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5575__S1 _1483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7233_ _0741_ _3081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7164_ _1475_ _3002_ _3020_ _1729_ _2999_ net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5495__A4 _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6115_ _2028_ _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7095_ _2978_ _2979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5327__S1 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6046_ _1959_ _0951_ _1960_ _1961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_29_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7997_ reg_file.reg_storage\[3\]\[8\] _3531_ _3775_ _3777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8063__I _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6948_ _1085_ _2837_ _2838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_49_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5955__A2 _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7157__A1 _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7157__B2 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6879_ _2444_ _2450_ _2516_ _2771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9667_ _0453_ clknet_leaf_0_clk reg_file.reg_storage\[15\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9598_ _0384_ clknet_leaf_81_clk reg_file.reg_storage\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6904__A1 _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8618_ _4180_ _4181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8549_ _4126_ _4138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output191_I net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9082__A1 _3945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8238__I _3927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8174__S _3872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4749__A3 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6371__A2 _2234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5557__S1 _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4609__C _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7920_ _3447_ _3712_ _3029_ _3713_ _3714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_7851_ _3640_ _3651_ _3652_ _3653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _1847_ _2697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7782_ net46 _3589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4994_ _0909_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7139__A1 _3007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9521_ _0307_ clknet_leaf_66_clk reg_file.reg_storage\[11\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6733_ _2625_ _2630_ _2631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9452_ _0238_ clknet_leaf_54_clk reg_file.reg_storage\[12\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8611__I _4172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6664_ _2153_ _2564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8403_ reg_file.reg_storage\[14\]\[16\] _4038_ _4047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5615_ _0528_ _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_34_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9383_ _0169_ clknet_4_2_0_clk reg_file.reg_storage\[14\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6595_ _2495_ _2268_ _2497_ _2498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6362__A2 _2231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8334_ _3725_ _3999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5546_ _0492_ _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5477_ reg_file.reg_storage\[12\]\[25\] reg_file.reg_storage\[13\]\[25\] reg_file.reg_storage\[14\]\[25\]
+ reg_file.reg_storage\[15\]\[25\] _1387_ _1388_ _1393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8265_ reg_file.reg_storage\[7\]\[9\] _3947_ _3948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7216_ _3058_ _3042_ _3065_ net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input48_I mem_ld_dat[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__I2 reg_file.reg_storage\[14\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8196_ _3682_ _3895_ _3898_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5873__A1 _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7147_ _1539_ _3012_ _3013_ net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_70_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7078_ _2103_ _1477_ _2963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6029_ _1294_ _1282_ _1944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6050__A1 _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9119__A2 _4496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5236__S0 _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7853__A2 _3237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9055__A1 _3911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8802__A1 reg_file.reg_storage\[11\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7605__A2 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_92_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5092__A2 _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7369__A1 _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8030__A2 _3791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6041__A1 _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_30_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5227__S0 _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6380_ _2288_ _2289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_51_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5400_ reg_file.reg_storage\[2\]\[3\] _0813_ _0814_ _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ reg_file.reg_storage\[8\]\[7\] reg_file.reg_storage\[9\]\[7\] reg_file.reg_storage\[10\]\[7\]
+ reg_file.reg_storage\[11\]\[7\] _0644_ _0645_ _1247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_23_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_45_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8050_ _3751_ _3758_ _3806_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7001_ _2830_ _2886_ _2889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5262_ _0885_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7844__A2 _3235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5193_ _0545_ _1108_ _0679_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_126_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8606__I _3420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_103_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5702__S1 _1536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8952_ reg_file.reg_storage\[9\]\[25\] _4357_ _4395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8883_ _4250_ _4348_ _4352_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_108_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7903_ _3547_ _3699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_78_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_90_clk clknet_4_14_0_clk clknet_leaf_90_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7834_ _3637_ _3638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8021__A2 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__I _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7765_ _3525_ _3573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_118_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4977_ _0842_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6716_ _2614_ net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9504_ _0290_ clknet_leaf_128_clk reg_file.reg_storage\[11\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7780__A1 _2508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7696_ _2309_ _3504_ _3508_ _3509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_46_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9435_ _0221_ clknet_leaf_97_clk reg_file.reg_storage\[13\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6647_ _2297_ _2500_ _2547_ _2548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7532__A1 _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9366_ _0152_ clknet_leaf_96_clk reg_file.reg_storage\[7\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6578_ _2444_ _2450_ _2480_ _2481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_59_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5529_ _0491_ _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8317_ _3695_ _3986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9297_ _0083_ clknet_leaf_71_clk reg_file.reg_storage\[2\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7835__A2 _3544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8248_ _3489_ _3935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output154_I net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8179_ reg_file.reg_storage\[6\]\[14\] _3882_ _3889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7420__I _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8012__A2 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_81_clk clknet_4_12_0_clk clknet_leaf_81_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8251__I _3501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4954__I _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4900_ _0807_ _0808_ _0812_ _0815_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5880_ _0885_ _0676_ _1795_ _1796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_72_clk clknet_4_9_0_clk clknet_leaf_72_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_75_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4831_ _0663_ _0746_ _0710_ _0709_ _0661_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_16_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6565__A2 _2381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7550_ _3368_ _1481_ _3372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4762_ _0622_ _0651_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_126_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6501_ _1787_ _2001_ _2407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6317__A2 _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4693_ _0588_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7481_ _3307_ _3308_ _3309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6432_ _2333_ _2339_ _2340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9220_ _0006_ clknet_leaf_17_clk reg_file.reg_storage\[5\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9151_ reg_file.reg_storage\[15\]\[4\] _4513_ _4519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8102_ reg_file.reg_storage\[2\]\[17\] _3831_ _3841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6363_ _2068_ _2265_ _2272_ _1983_ _2273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_12_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9082_ _3945_ _4462_ _4476_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6294_ _1280_ _1805_ _2204_ _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5314_ _1217_ _1086_ _1229_ _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8490__A2 _4099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8033_ reg_file.reg_storage\[3\]\[24\] _3758_ _3797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5245_ _1151_ _1160_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4864__I _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5176_ _0863_ reg_file.reg_storage\[2\]\[27\] _0764_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8935_ _4220_ _4381_ _4385_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_63_clk clknet_4_11_0_clk clknet_leaf_63_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8866_ reg_file.reg_storage\[10\]\[23\] _4311_ _4343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8797_ _4246_ _4298_ _4300_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5695__I _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7817_ _3613_ _3621_ _3622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_65_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7748_ reg_file.reg_storage\[5\]\[10\] _3557_ _3492_ _3558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7679_ _3493_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9418_ _0204_ clknet_leaf_8_clk reg_file.reg_storage\[13\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9349_ _0135_ clknet_leaf_40_clk reg_file.reg_storage\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7659__I2 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7808__A2 _3472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8481__A2 _4088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5819__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5678__S0 _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6244__A1 _2153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_54_clk clknet_4_10_0_clk clknet_leaf_54_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7744__A1 _3547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6547__A2 _2450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4653__S1 _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__S0 _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7325__I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4581__I1 reg_file.reg_storage\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5030_ _0649_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4684__I net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6981_ _2704_ _2868_ _2869_ _2870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_49_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6235__A1 _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8720_ reg_file.reg_storage\[8\]\[31\] _4173_ _4253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5932_ _1541_ _1848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__4797__A1 _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_45_clk clknet_4_8_0_clk clknet_leaf_45_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8651_ _3555_ _4205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7735__A1 _3428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5863_ _1778_ _0697_ _1779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7602_ _3398_ _3422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8582_ reg_file.reg_storage\[12\]\[21\] _4152_ _4157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5794_ _1709_ _1582_ _1584_ _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_7_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4814_ _0713_ _0729_ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_133_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4745_ _0601_ _0590_ _0591_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7533_ _3345_ _3356_ _3357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_134_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4676_ _0587_ _0593_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7464_ _3284_ _3274_ _3293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9203_ _4505_ _4548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4859__I _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7395_ net72 _1585_ _3230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6415_ _2165_ _2321_ _2322_ _2323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_9134_ _4505_ _4506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_116_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6346_ _2135_ _2253_ _2255_ _2256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9065_ reg_file.reg_storage\[4\]\[2\] _3455_ _4466_ _4467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8016_ _3638_ _3784_ _3787_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5116__I3 reg_file.reg_storage\[7\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6277_ _1998_ _2189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8463__A2 _4075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6474__A1 _2110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5228_ _1136_ _1140_ _1142_ _1143_ _0964_ _0946_ _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA_input30_I inst[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5159_ reg_file.reg_storage\[4\]\[26\] reg_file.reg_storage\[5\]\[26\] reg_file.reg_storage\[6\]\[26\]
+ reg_file.reg_storage\[7\]\[26\] _0990_ _0984_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4580__S0 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_16_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_67_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output117_I net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8918_ _4202_ _4362_ _4376_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8849_ _4333_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5201__A2 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_25_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_133_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4960__A1 _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4769__I _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7965__A1 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_clk clknet_4_3_0_clk clknet_leaf_27_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7717__A1 _2350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5823__S0 _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4679__I net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7180_ _2971_ _3033_ net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6200_ _2041_ _2108_ _2112_ _2113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4703__A1 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6131_ _2044_ _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8087__S _3828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6062_ _1242_ _1977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5013_ _0787_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_144_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6964_ _2015_ _2849_ _2853_ _2854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_49_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_18_clk clknet_4_6_0_clk clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8614__I _3442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8703_ _4172_ _4241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9683_ _0469_ clknet_leaf_75_clk reg_file.reg_storage\[15\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6895_ _2769_ _2786_ _2787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5915_ _1228_ _1827_ _1754_ _1830_ _1216_ _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_91_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8550__S _4138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8634_ _3489_ _4193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5846_ _0489_ _0564_ _0673_ _0674_ _1762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_36_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4617__S1 _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8565_ _4127_ _4147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6931__A2 _2607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5777_ _1691_ _1692_ _0978_ _1693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8133__A1 _3746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8496_ _3978_ _4101_ _4103_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4728_ _0632_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_17_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7516_ net82 _3326_ _3322_ _3341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_31_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4659_ _0539_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input78_I pc[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7447_ _1525_ _3278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7378_ net71 _3205_ _3214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9117_ _3992_ _4456_ _4495_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6329_ _1805_ _2204_ _2239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9048_ reg_file.reg_storage\[1\]\[31\] _4449_ _4453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8524__I _4119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__A2 _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8460__S _4079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7175__A2 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8124__A1 _3719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7722__I1 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8675__A2 _4214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5489__A2 _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7635__B1 _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8635__S _4187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5661__A2 _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4962__I _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6610__A1 _2398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5700_ reg_file.reg_storage\[12\]\[18\] reg_file.reg_storage\[13\]\[18\] reg_file.reg_storage\[14\]\[18\]
+ reg_file.reg_storage\[15\]\[18\] _1615_ _0879_ _1616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_128_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6680_ _2575_ _2577_ _2579_ _2580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8363__A1 _3865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5177__A1 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5631_ _1432_ reg_file.reg_storage\[2\]\[23\] _1486_ _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_73_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8350_ _4010_ _4001_ _4011_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5272__S1 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5562_ _1029_ _1477_ _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8281_ _3922_ _3959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7301_ _3121_ _3136_ _3143_ net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8666__A2 _4214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5493_ _1098_ _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7232_ _3078_ _3079_ _3080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__7941__C _3732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_7_clk clknet_4_6_0_clk clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7163_ net220 _3002_ _3020_ _1717_ _2998_ net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_111_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8609__I _4172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8418__A2 _4051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7094_ _2977_ _2978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_95_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6114_ _1977_ _2028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5101__A1 _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6045_ _1217_ _0875_ _1960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8545__S _4132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8344__I _4006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4872__I _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7996_ _3776_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _2834_ _2836_ _2837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_49_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8354__A1 _4013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6878_ _1820_ _2488_ _2770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9666_ _0452_ clknet_leaf_5_clk reg_file.reg_storage\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9597_ _0383_ clknet_leaf_107_clk reg_file.reg_storage\[9\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8617_ _4179_ _4180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5168__A1 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5829_ _1734_ _1744_ _1745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_134_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8548_ _3938_ _4128_ _4137_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output184_I net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8479_ _4093_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8409__A2 _4044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4694__A3 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__A2 _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9082__A2 _4462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6840__A1 _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7148__A2 _1575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5882__A2 _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9073__A2 _4463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_128_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7850_ _3525_ _3652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_4_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6801_ _2696_ net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_81_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7781_ net54 _3588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_4993_ _0794_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9520_ _0306_ clknet_leaf_68_clk reg_file.reg_storage\[11\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6732_ _0950_ _2629_ _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_74_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6663_ _1719_ _1731_ _2563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9451_ _0237_ clknet_leaf_2_clk reg_file.reg_storage\[12\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_139_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ reg_file.reg_storage\[4\]\[21\] reg_file.reg_storage\[5\]\[21\] reg_file.reg_storage\[6\]\[21\]
+ reg_file.reg_storage\[7\]\[21\] _1368_ _1425_ _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8402_ _4046_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9382_ _0168_ clknet_leaf_44_clk reg_file.reg_storage\[14\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6594_ _2495_ _2496_ _2497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8333_ _3996_ _3915_ _3998_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5545_ _1442_ _1460_ _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8639__A2 _4182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5476_ reg_file.reg_storage\[1\]\[25\] _1391_ _1388_ _1392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8264_ _3921_ _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8339__I _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8195_ reg_file.reg_storage\[6\]\[21\] _3893_ _3898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_57_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7215_ _3059_ net119 _3061_ _3064_ _3065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7146_ net161 _3004_ _3013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5712__I3 reg_file.reg_storage\[15\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7077_ _2961_ _2171_ _2074_ _2962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5625__A2 _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6028_ _1299_ _1937_ _1939_ _1942_ _1943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5698__I _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4816__B _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7378__A2 _3205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7979_ _3762_ _3766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8327__A1 reg_file.reg_storage\[7\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9649_ _0435_ clknet_leaf_71_clk reg_file.reg_storage\[4\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5236__S1 _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8878__A2 _4346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7550__A2 _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5164__I1 reg_file.reg_storage\[13\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5313__A1 _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9055__A2 _4456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6813__A1 _2122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7369__A2 _3205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7756__C _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5227__S1 _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7541__A2 _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5330_ reg_file.reg_storage\[12\]\[7\] reg_file.reg_storage\[13\]\[7\] reg_file.reg_storage\[14\]\[7\]
+ reg_file.reg_storage\[15\]\[7\] _0644_ _0645_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_51_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5261_ _1164_ _1176_ _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7000_ _1409_ _2859_ _2888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5192_ _1105_ _1107_ _0739_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7057__A1 _2122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8951_ _4236_ _4356_ _4394_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7902_ _3417_ _3698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7012__B _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8882_ reg_file.reg_storage\[10\]\[30\] _4305_ _4352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4910__S0 _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7833_ net104 _3601_ _3633_ _3636_ _3637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_93_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7764_ _3484_ _3572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5091__I0 _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4976_ _0756_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6715_ _1984_ _2601_ _2613_ _2614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9503_ _0289_ clknet_leaf_123_clk reg_file.reg_storage\[11\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6142__I _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7695_ _3116_ _3505_ _3506_ _0595_ _3507_ _3508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_9434_ _0220_ clknet_leaf_97_clk reg_file.reg_storage\[13\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6646_ _2047_ _2546_ _2547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9365_ _0151_ clknet_leaf_23_clk reg_file.reg_storage\[7\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_59_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6577_ _1817_ _2442_ _2480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5543__A1 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8316_ _3984_ _3975_ _3985_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5528_ _0740_ _1443_ _1414_ _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input60_I mem_ld_dat[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9296_ _0082_ clknet_leaf_46_clk reg_file.reg_storage\[2\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5459_ _0672_ _1374_ _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8247_ _3933_ _3923_ _3934_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8178_ _3868_ _3888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5846__A2 _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output147_I net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7129_ _2978_ _3001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5457__S1 _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8532__I _4126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8720__A1 reg_file.reg_storage\[8\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7287__B2 _3130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9028__A2 _4437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5837__A2 _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6655__C _2555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4648__I0 reg_file.reg_storage\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5131__I _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8442__I _4067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4830_ _0662_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_16_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_103_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4761_ _0676_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6500_ _2404_ _2405_ _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _0607_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7480_ _1046_ _1881_ _3308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5525__A1 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6431_ _2197_ _2338_ _2183_ _2339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ _1938_ _2231_ _2266_ _2271_ _2272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9150_ _4518_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8101_ _3638_ _3837_ _3840_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5313_ _1228_ _1058_ _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9081_ reg_file.reg_storage\[4\]\[9\] _4475_ _4476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6293_ _1765_ _2155_ _2153_ _2204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__9019__A2 _4430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8032_ _3696_ _3766_ _3796_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_54_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5244_ _1014_ _1159_ _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5175_ _0861_ reg_file.reg_storage\[3\]\[27\] _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6846__B _2739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8617__I _4179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5136__S0 _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8934_ reg_file.reg_storage\[9\]\[17\] _4375_ _4385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5041__I _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8865_ _4232_ _4338_ _4342_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8352__I _4012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7816_ _3547_ _3618_ _3620_ _3621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_137_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8796_ reg_file.reg_storage\[11\]\[28\] _4296_ _4300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7747_ _3556_ _3557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5764__A1 _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _0830_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7678_ reg_file.reg_storage\[5\]\[5\] _3491_ _3492_ _3493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_91_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9417_ _0203_ clknet_leaf_51_clk reg_file.reg_storage\[13\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6629_ _1984_ _2519_ _2530_ _2531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7505__A2 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_89_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_9348_ _0134_ clknet_leaf_17_clk reg_file.reg_storage\[7\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7659__I3 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9279_ _0065_ clknet_leaf_121_clk reg_file.reg_storage\[2\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7431__I _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5678__S1 _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_98_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7992__A2 _3766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_44_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8262__I _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4558__A2 _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_102_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__S1 _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6180__A1 _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4581__I2 reg_file.reg_storage\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_117_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6483__A2 _1832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6980_ _2177_ _2659_ _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7432__A1 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _0829_ _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_105_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5994__A1 _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8650_ _4202_ _4182_ _4204_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5862_ _1777_ _1118_ _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4633__C _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8581_ _3978_ _4154_ _4156_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7601_ _3420_ _3421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5793_ _0712_ _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4813_ _0727_ _0708_ _0728_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_90_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7532_ _1088_ _3341_ _3356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8900__I _4365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4744_ _0652_ _0657_ _0659_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_126_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9202_ _3995_ _4506_ _4547_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8160__A2 _3870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4675_ _0592_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7463_ net80 _3292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7394_ _3227_ _3228_ _3229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_12_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6414_ _2316_ _2320_ _2322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_9133_ _4504_ _4505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_116_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6345_ _2179_ _2254_ _2255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8999__A1 _3945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6276_ _2114_ _2187_ _2188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9064_ _4465_ _4466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8347__I _3745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8015_ reg_file.reg_storage\[3\]\[16\] _3778_ _3787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6474__A2 _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5227_ reg_file.reg_storage\[8\]\[13\] reg_file.reg_storage\[9\]\[13\] reg_file.reg_storage\[10\]\[13\]
+ reg_file.reg_storage\[11\]\[13\] _1049_ _1141_ _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__7251__I net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__S1 _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input23_I inst[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5158_ net83 _0750_ _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5089_ reg_file.reg_storage\[12\]\[29\] reg_file.reg_storage\[13\]\[29\] reg_file.reg_storage\[14\]\[29\]
+ reg_file.reg_storage\[15\]\[29\] _0999_ _0903_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_79_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8917_ reg_file.reg_storage\[9\]\[9\] _4375_ _4376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_67_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8848_ reg_file.reg_storage\[10\]\[15\] _4216_ _4315_ _4333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6529__A3 _2080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8779_ _4228_ _4288_ _4290_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5596__S0 _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7965__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5520__S0 _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8921__S _4372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7717__A2 _3504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5823__S1 _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__S0 _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5900__A1 _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6130_ _1111_ _2044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4695__I _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8167__I _3867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6061_ _1335_ _1971_ _1347_ _1975_ _1976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5012_ reg_file.reg_storage\[12\]\[16\] reg_file.reg_storage\[13\]\[16\] reg_file.reg_storage\[14\]\[16\]
+ reg_file.reg_storage\[15\]\[16\] _0780_ _0781_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_144_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6963_ _2841_ _2834_ _2074_ _2852_ _2853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_49_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8702_ _3718_ _4240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9682_ _0468_ clknet_leaf_75_clk reg_file.reg_storage\[15\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6894_ _2777_ _2780_ _2785_ _2786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_76_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5914_ _1828_ _1829_ _1379_ _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5719__A1 _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8633_ _4191_ _4182_ _4192_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5845_ _1264_ _1760_ _1761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_24_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8381__A2 _4025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5776_ _0705_ _1581_ _1583_ _1692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_8_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8564_ _4146_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8495_ reg_file.reg_storage\[13\]\[20\] _4099_ _4103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4727_ reg_file.reg_storage\[1\]\[0\] _0639_ _0642_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7515_ _3337_ _3339_ _3340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6144__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7446_ _3274_ _3276_ _3277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4658_ _0481_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_32_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6695__A2 _2398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput90 pc[3] net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_101_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9116_ reg_file.reg_storage\[4\]\[25\] _4457_ _4495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7377_ _0911_ _1585_ _3213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4589_ _0482_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_101_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _2094_ _2149_ _2237_ _2150_ _2238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_9047_ _4009_ _4407_ _4452_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6259_ _2170_ _2171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_4_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7947__A2 _3366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8124__A2 _3812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7635__B2 _3402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7820__S _3569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5949__A1 _1635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8060__A1 _3753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5630_ _1429_ reg_file.reg_storage\[3\]\[23\] _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5561_ _1379_ _1475_ _1476_ _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_143_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8280_ _3957_ _3958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8115__A2 _3844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5492_ _1399_ _1407_ _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7300_ _3100_ net128 _3101_ _3142_ _3143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7874__A1 net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7231_ _3058_ _3067_ _3079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_113_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7874__B2 _3673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8098__S _3821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7162_ net223 _3002_ _3020_ _1702_ _2997_ net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_95_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7093_ _2976_ _2977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6113_ _2016_ _2027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6044_ _1669_ _1959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4860__A1 _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8625__I _4186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7995_ reg_file.reg_storage\[3\]\[7\] _3511_ _3775_ _3776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6946_ _2721_ _2743_ _2766_ _2835_ _2836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__6601__A2 _2503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_53_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8561__S _4131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _1057_ _2768_ _2769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9665_ _0451_ clknet_leaf_133_clk reg_file.reg_storage\[15\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5799__S0 _1607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9596_ _0382_ clknet_leaf_101_clk reg_file.reg_storage\[9\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8616_ _4124_ _4178_ _4179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5828_ _1735_ _1743_ _1744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_input90_I pc[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6365__A1 _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5759_ reg_file.reg_storage\[1\]\[10\] _1674_ _1672_ _1675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8547_ reg_file.reg_storage\[12\]\[6\] _4129_ _4137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6117__A1 _2030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7865__A1 net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8478_ reg_file.reg_storage\[13\]\[13\] _3955_ _4078_ _4093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_142_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7865__B2 _3665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7429_ _0952_ _3251_ _3261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7617__A1 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8042__A1 _3726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8270__I _3566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5714__S0 _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4973__I _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6800_ _2680_ _2683_ _2688_ _2695_ _2696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__8584__A2 _4127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4992_ net73 _0889_ _0891_ _0907_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_7780_ _2508_ _3460_ _3587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6731_ _1858_ _2628_ _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_46_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6662_ _1601_ _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_73_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9450_ _0236_ clknet_leaf_6_clk reg_file.reg_storage\[12\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_139_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ reg_file.reg_storage\[12\]\[21\] reg_file.reg_storage\[13\]\[21\] reg_file.reg_storage\[14\]\[21\]
+ reg_file.reg_storage\[15\]\[21\] _1368_ _1421_ _1529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_9381_ _0167_ clknet_leaf_39_clk reg_file.reg_storage\[14\]\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8401_ reg_file.reg_storage\[14\]\[15\] _3961_ _4028_ _4046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8332_ reg_file.reg_storage\[7\]\[26\] _3997_ _3998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6593_ _2170_ _2496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5309__I _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5544_ _1459_ _1056_ _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5475_ reg_file.reg_storage\[2\]\[25\] reg_file.reg_storage\[3\]\[25\] _1390_ _1391_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8263_ _3945_ _3946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8194_ _3675_ _3895_ _3897_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7214_ _3058_ _1238_ _3063_ _3064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7145_ _3001_ _3012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5086__A1 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7076_ _2103_ _1477_ _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6027_ _1299_ _1941_ _1942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_61_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8575__A2 _4152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7978_ _3764_ _3765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5633__I0 reg_file.reg_storage\[12\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6929_ _2217_ _2709_ _2820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_119_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9648_ _0434_ clknet_leaf_70_clk reg_file.reg_storage\[4\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7535__B1 _3357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5219__I _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_9579_ _0365_ clknet_leaf_1_clk reg_file.reg_storage\[9\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5561__A2 _1475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8566__A2 _4141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7774__B1 _3573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6329__A1 _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_109_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5001__A1 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__S _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6501__A1 _1787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5260_ _1175_ _1148_ _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_118_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5191_ _1106_ _0618_ _0616_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8950_ reg_file.reg_storage\[9\]\[24\] _4357_ _4394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7901_ _3444_ _3696_ _3697_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_39_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8881_ _4248_ _4348_ _4351_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_108_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4910__S1 _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7832_ _3607_ _3212_ _3634_ _3635_ _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_121_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4975_ _0890_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7763_ _2479_ _3460_ _3571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_127_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5240__A1 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9502_ _0288_ clknet_leaf_109_clk reg_file.reg_storage\[11\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6714_ _1935_ _2570_ _2609_ _2610_ _1636_ _2612_ _2613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_9433_ _0219_ clknet_leaf_97_clk reg_file.reg_storage\[13\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7694_ _3047_ _3115_ _3430_ _3507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_132_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6645_ _1955_ _2335_ _1952_ _2546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_143_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9364_ _0150_ clknet_leaf_22_clk reg_file.reg_storage\[7\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_59_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6576_ _2479_ net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__5543__A2 _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9295_ _0081_ clknet_leaf_58_clk reg_file.reg_storage\[2\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8315_ reg_file.reg_storage\[7\]\[22\] _3922_ _3985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5527_ _1412_ _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4878__I _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8246_ reg_file.reg_storage\[7\]\[4\] _3924_ _3934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7296__A2 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input53_I mem_ld_dat[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_136_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5458_ _0492_ _1373_ _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_30_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8177_ _3887_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5389_ reg_file.reg_storage\[12\]\[2\] reg_file.reg_storage\[13\]\[2\] reg_file.reg_storage\[14\]\[2\]
+ reg_file.reg_storage\[15\]\[2\] _0919_ _1301_ _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7128_ _2979_ _3000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5449__I3 reg_file.reg_storage\[7\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7059_ _2941_ _2944_ _2945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5502__I _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8548__A2 _4128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7756__B1 _3546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8813__I _4311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4665__S0 _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6731__A1 _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5090__S0 _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4788__I _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7287__A2 net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5298__A1 _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6508__I net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5222__A1 _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6970__A1 _2856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4760_ _0622_ _0651_ _0660_ _0672_ net216 _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4691_ net26 _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_136_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8711__A2 _4241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5525__A2 _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6430_ _2334_ _2337_ _2338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6361_ _2267_ _2268_ _2270_ _2271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8100_ reg_file.reg_storage\[2\]\[16\] _3831_ _3840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5312_ _1227_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_140_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9080_ _4460_ _4475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5289__A1 _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6292_ _2203_ net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5243_ _1152_ _1156_ _1157_ _1158_ _0965_ _1025_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_87_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8031_ reg_file.reg_storage\[3\]\[23\] _3764_ _3796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5174_ reg_file.reg_storage\[1\]\[27\] _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8778__A2 _4286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5136__S1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6789__A1 _2684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8933_ _4218_ _4381_ _4384_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8864_ reg_file.reg_storage\[10\]\[22\] _4311_ _4342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6354__S _2022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7815_ _3572_ _3202_ _3486_ _3619_ _3620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_8795_ _4243_ _4298_ _4299_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6153__I _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7746_ _3555_ _3556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5764__A2 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4958_ _0853_ _0873_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_47_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4889_ reg_file.reg_storage\[4\]\[21\] reg_file.reg_storage\[5\]\[21\] reg_file.reg_storage\[6\]\[21\]
+ reg_file.reg_storage\[7\]\[21\] _0802_ _0804_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7677_ _3427_ _3492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_46_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9416_ _0202_ clknet_leaf_52_clk reg_file.reg_storage\[13\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6713__A1 _1635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6628_ _2296_ _2522_ _2526_ _2342_ _2529_ _2530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4602__S _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4575__I0 reg_file.reg_storage\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_9347_ _0133_ clknet_leaf_136_clk reg_file.reg_storage\[7\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ _2407_ _2463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_42_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9278_ _0064_ clknet_leaf_116_clk reg_file.reg_storage\[2\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8229_ _3424_ _3761_ _3920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8218__A1 _3751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8769__A2 _4281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7441__A2 net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9194__A2 _4511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8941__A2 _4388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6952__A1 _2841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6704__A1 _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_131_clk clknet_4_4_0_clk clknet_leaf_131_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8919__S _4372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4581__I3 reg_file.reg_storage\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5140__B1 _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4981__I _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5930_ _1578_ _1846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_49_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8453__I _4078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8932__A2 _4375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5861_ _1312_ _1321_ _1777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7600_ net65 _3401_ _0689_ _3403_ _3419_ _3420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_118_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8580_ reg_file.reg_storage\[12\]\[20\] _4152_ _4156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5792_ _1146_ _1707_ _1708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4812_ _0700_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4743_ _0658_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7531_ _3345_ _3346_ _3354_ _3355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7462_ _3076_ _3285_ _3290_ _3046_ _3291_ net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_9201_ reg_file.reg_storage\[15\]\[26\] _4546_ _4547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4674_ _0588_ _0589_ _0590_ _0591_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6413_ _2316_ _2320_ _2321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_102_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6171__A2 _1996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7393_ _1705_ _1633_ _3228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_3_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9132_ _3754_ _4015_ _4504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6344_ _2110_ _2029_ _1044_ _2254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7120__A1 net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8999__A2 _4411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9063_ _4459_ _4465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6275_ _2063_ _1179_ _2186_ _2187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__8628__I _3468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8014_ _3786_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5226_ reg_file.reg_storage\[12\]\[13\] reg_file.reg_storage\[13\]\[13\] reg_file.reg_storage\[14\]\[13\]
+ reg_file.reg_storage\[15\]\[13\] _1049_ _1141_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_110_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ _1059_ _1072_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5088_ _0765_ _1001_ _1002_ _1003_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7423__A2 _3255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8916_ _4360_ _4375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_67_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4891__I _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7974__A3 _3394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I inst[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8847_ _4213_ _4331_ _4332_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8778_ reg_file.reg_storage\[11\]\[20\] _4286_ _4290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7729_ _3515_ _3538_ _3539_ _3540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_105_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_113_clk clknet_4_13_0_clk clknet_leaf_113_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5596__S1 _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8739__S _4266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8439__A1 _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7111__A1 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8538__I _4131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8474__S _4085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4720__I0 reg_file.reg_storage\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7414__A2 _3237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8273__I _3583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5520__S1 _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6925__A1 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_104_clk clknet_4_13_0_clk clknet_leaf_104_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_100_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5587__S1 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4976__I _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8448__I _4074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5339__S1 _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input8_I inst[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6060_ _1972_ _1348_ _1974_ _1975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5011_ net9 _0926_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_90_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6962_ _2850_ _2168_ _2851_ _2852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5967__A2 _1881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7169__A1 _2969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8701_ _4238_ _4174_ _4239_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9681_ _0467_ clknet_leaf_31_clk reg_file.reg_storage\[15\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6893_ _2781_ _2782_ _2783_ _2784_ _2779_ _2667_ _2785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_76_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5913_ net22 _1411_ _1829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__7955__C _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8911__I _4360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8632_ reg_file.reg_storage\[8\]\[4\] _4183_ _4192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8905__A2 _4363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5844_ _1758_ _1759_ _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_118_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_62_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8563_ reg_file.reg_storage\[12\]\[13\] _3955_ _4131_ _4146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5775_ _1690_ _1691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7514_ _3330_ _3331_ _3338_ _3339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_118_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8494_ _3974_ _4101_ _4102_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4726_ _0641_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_142_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4657_ _0576_ net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8559__S _4138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7445_ _3260_ _3261_ _3275_ _3276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_141_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7892__A2 _3458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput91 pc[4] net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput80 pc[23] net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7376_ _0911_ _3211_ _3212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_13_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4886__I _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9115_ _3989_ _4456_ _4494_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6327_ _2161_ _2162_ _2205_ _2237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4588_ _0495_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_43_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9046_ reg_file.reg_storage\[1\]\[30\] _4449_ _4452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6258_ _0731_ _1345_ _2170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5209_ reg_file.reg_storage\[2\]\[12\] reg_file.reg_storage\[3\]\[12\] _0920_ _1125_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6189_ _2098_ _2100_ _2101_ _2102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output122_I net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_58_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6606__I _2508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_101_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6080__A1 _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6907__A1 _2797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_116_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9383__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6341__I _1787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4796__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6843__B1 _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5949__A2 _1636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8060__A2 _3808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__A1 _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8731__I _4261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__S0 _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5560_ _1353_ _1400_ _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5491_ _1401_ _1404_ _1405_ _1406_ _1407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_14_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7230_ net91 _3078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7874__A2 _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7161_ net234 _3018_ _3020_ _1690_ _2996_ net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_TAPCELL_ROW_113_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8178__I _3868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7092_ _1709_ _0714_ _2975_ _2976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6112_ _1998_ _2026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7015__C _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7626__A2 _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6043_ _1954_ _1957_ _1268_ _1958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_1_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7994_ _3763_ _3775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6870__B _2762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6945_ _2807_ _2797_ _2672_ _2835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_124_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8641__I _4180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _1459_ _2767_ _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9664_ _0450_ clknet_leaf_133_clk reg_file.reg_storage\[15\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5799__S1 _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9595_ _0381_ clknet_leaf_100_clk reg_file.reg_storage\[9\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8615_ _1236_ _3387_ _4178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_63_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5827_ _0669_ _1742_ _1743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_29_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5758_ reg_file.reg_storage\[2\]\[10\] reg_file.reg_storage\[3\]\[10\] _1614_ _1674_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8546_ _4136_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input83_I pc[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4709_ net9 _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_8477_ _4092_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_75_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5689_ _0534_ _1605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7428_ net77 _3260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7865__A2 _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__I _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7359_ _3192_ _1710_ _3197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_9_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9029_ reg_file.reg_storage\[1\]\[23\] _4410_ _4442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8290__A2 _3959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6336__I _2120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__A1 _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6272__S _2183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__I1 reg_file.reg_storage\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5867__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5714__S1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5478__S0 _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4991_ _0894_ _0901_ _0904_ _0905_ _0906_ _0788_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_105_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _2565_ _2627_ _2628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6661_ _2560_ _2561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_34_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8400_ _3958_ _4044_ _4045_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5612_ reg_file.reg_storage\[1\]\[21\] _1527_ _1425_ _1528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6592_ _2494_ _2483_ _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9380_ _0166_ clknet_leaf_15_clk reg_file.reg_storage\[14\]\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_139_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8331_ _3913_ _3997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5543_ _1114_ _1444_ _1458_ _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_6_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7805__I _3610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7847__A2 _3544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5474_ _0659_ _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8262_ _3542_ _3945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5858__A1 _1767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8837__S _4322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9049__A1 _4012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8193_ reg_file.reg_storage\[6\]\[20\] _3893_ _3897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7026__B _2076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7213_ _3054_ _3055_ _3062_ _3063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5325__I _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5402__S0 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__I3 reg_file.reg_storage\[7\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7144_ _0555_ _3010_ _3011_ net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_100_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7075_ _2257_ _2958_ _2959_ _2960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6026_ _1734_ _1282_ _1940_ _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8024__A2 _3791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7977_ _3763_ _3764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8371__I _4028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6928_ _2036_ _2817_ _2818_ _2819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9647_ _0433_ clknet_leaf_62_clk reg_file.reg_storage\[4\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6859_ _2751_ _1917_ _2752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9578_ _0364_ clknet_leaf_3_clk reg_file.reg_storage\[9\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8529_ _3395_ _4117_ _4124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_60_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6649__I0 _2301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8015__A2 _3778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_84_clk clknet_4_14_0_clk clknet_leaf_84_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6026__A1 _1734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8281__I _3922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7774__B2 _3580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6329__A2 _2204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7625__I _3426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4760__B2 _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5145__I _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5190_ net2 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__8254__A2 _3923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8392__S _4035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7900_ reg_file.reg_storage\[5\]\[23\] _3458_ _3697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8880_ reg_file.reg_storage\[10\]\[29\] _4346_ _4351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_75_clk clknet_4_9_0_clk clknet_leaf_75_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_108_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6568__A2 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7831_ _1585_ _3439_ _3635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7762_ _3570_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4974_ _0753_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7693_ net62 net48 net39 net57 _3021_ _3025_ _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_129_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9501_ _0287_ clknet_leaf_107_clk reg_file.reg_storage\[8\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6713_ _1635_ _2169_ _2611_ _2174_ _2612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_59_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7517__A1 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9432_ _0218_ clknet_leaf_89_clk reg_file.reg_storage\[13\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6644_ _2251_ _2542_ _2544_ _2545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9363_ _0149_ clknet_leaf_79_clk reg_file.reg_storage\[7\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6575_ _2451_ _2462_ _2466_ _2296_ _2478_ _2479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_143_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9294_ _0080_ clknet_4_11_0_clk reg_file.reg_storage\[2\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8314_ _3983_ _3984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5526_ _1409_ _1441_ _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5483__C _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5457_ _1365_ _1367_ _1370_ _1371_ _1372_ _1105_ _1373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA_rebuffer19_I _1618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8245_ _3932_ _3933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8493__A2 _4099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7296__A3 _3138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input46_I mem_ld_dat[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8176_ reg_file.reg_storage\[6\]\[13\] _3598_ _3872_ _3887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5388_ reg_file.reg_storage\[1\]\[2\] _1303_ _1301_ _1304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7127_ _1729_ _2995_ _2999_ net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4894__I _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8366__I _4024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7058_ _1043_ _2942_ _2943_ _2120_ _2944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6009_ _1042_ _1924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_66_clk clknet_4_11_0_clk clknet_leaf_66_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_83_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7756__B2 _3563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7756__A1 _3161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4665__S1 _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7508__A1 _3035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5090__S1 _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6495__A1 _2398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8276__I _3596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6247__A1 _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6798__A2 _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_57_clk clknet_4_10_0_clk clknet_leaf_57_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4690_ net65 _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_136_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4979__I reg_file.reg_storage\[1\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6722__A2 _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6360_ _2267_ _2269_ _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ _1218_ _1225_ _1226_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8030_ _3689_ _3791_ _3795_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_load_slew1_I _2413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5289__A2 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6291_ _2164_ _2166_ _2202_ _2203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5242_ reg_file.reg_storage\[8\]\[14\] reg_file.reg_storage\[9\]\[14\] reg_file.reg_storage\[10\]\[14\]
+ reg_file.reg_storage\[11\]\[14\] _1021_ _1022_ _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_121_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5173_ reg_file.reg_storage\[4\]\[27\] reg_file.reg_storage\[5\]\[27\] reg_file.reg_storage\[6\]\[27\]
+ reg_file.reg_storage\[7\]\[27\] _1061_ _1063_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xinput1 inst[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8932_ reg_file.reg_storage\[9\]\[16\] _4375_ _4384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_48_clk clknet_4_10_0_clk clknet_leaf_48_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8863_ _4230_ _4338_ _4341_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5461__A2 _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6434__I _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7814_ _3205_ _3438_ _3619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8794_ reg_file.reg_storage\[11\]\[27\] _4296_ _4299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7745_ net233 _3504_ _3554_ _3555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_93_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4957_ _0800_ _0872_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4888_ _0803_ _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_62_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7676_ _3490_ _3491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9415_ _0201_ clknet_leaf_35_clk reg_file.reg_storage\[13\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6627_ _2509_ _2510_ _2372_ _2528_ _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_132_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4575__I1 reg_file.reg_storage\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _2443_ _2461_ _2351_ _2462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_9346_ _0132_ clknet_leaf_6_clk reg_file.reg_storage\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9277_ _0063_ clknet_leaf_78_clk reg_file.reg_storage\[3\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5509_ _1421_ _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6489_ _1217_ _2392_ _2393_ _2319_ _1734_ _2395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_140_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7674__B1 _3483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8228_ _3918_ _3919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output152_I net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8159_ _3877_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5513__I _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_39_clk clknet_4_2_0_clk clknet_leaf_39_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5835__S0 _1532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6952__A2 _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7901__A1 _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7903__I _3547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6468__A1 _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_9_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5140__A1 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5140__B2 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ _1335_ _1178_ _1776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4811_ net5 _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_132_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5791_ _1703_ _1706_ _1707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_127_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7530_ _3313_ _3348_ _3353_ _3354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4742_ _0556_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_114_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4673_ net26 net23 _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
X_7461_ _3272_ net111 _3291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9200_ _4504_ _4546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4706__A1 _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6412_ _1228_ _2319_ _2320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7392_ net73 _3227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_116_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9131_ _4012_ _4457_ _4503_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6343_ _2019_ _2009_ _2010_ _2253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__9006__S _4414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9062_ _3918_ _4462_ _4464_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6274_ _2185_ _0974_ _2186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8013_ reg_file.reg_storage\[3\]\[15\] _3624_ _3768_ _3786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5225_ _0642_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5682__A2 _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__I _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5156_ _1071_ _0796_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5087_ _0773_ reg_file.reg_storage\[2\]\[29\] _0899_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8644__I _3529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8915_ _4374_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_2_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8846_ reg_file.reg_storage\[10\]\[14\] _4325_ _4332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8777_ _4225_ _4288_ _4289_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5709__S _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5989_ _1903_ _0730_ _0695_ _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5737__A3 _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7728_ _3525_ _3539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8136__A1 _3388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7659_ net59 net36 net45 net53 _3028_ _3410_ _3475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_133_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9329_ _0115_ clknet_leaf_70_clk reg_file.reg_storage\[6\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8439__A2 _4015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8755__S _4272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput190 net190 pc_next[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_27_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4720__I1 reg_file.reg_storage\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8554__I _4126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8127__A1 _3726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6802__I _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_133_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8678__A2 _4223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8729__I _4259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8850__A2 _4325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5010_ reg_file.reg_storage\[8\]\[16\] reg_file.reg_storage\[9\]\[16\] reg_file.reg_storage\[10\]\[16\]
+ reg_file.reg_storage\[11\]\[16\] _0780_ _0781_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6861__A1 _2038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8464__I _4073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6185__S _2097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5102__B _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8700_ reg_file.reg_storage\[8\]\[25\] _4175_ _4239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6961_ _2850_ _2496_ _2851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9680_ _0466_ clknet_leaf_33_clk reg_file.reg_storage\[15\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6892_ _1843_ _2745_ _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5912_ _0493_ _1751_ _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_49_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8631_ _3477_ _4191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ _0489_ _0575_ _0691_ _0674_ _1759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_124_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5719__A3 _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8562_ _4145_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5774_ _1622_ _1689_ _1690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7513_ _3326_ _1356_ _3338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8493_ reg_file.reg_storage\[13\]\[19\] _4099_ _4102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4725_ _0640_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_126_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4656_ _0494_ _0575_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7444_ net78 _3275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4587_ _0512_ net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7375_ _1165_ _3201_ _3211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput70 pc[14] net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput81 pc[24] net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_130_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9114_ reg_file.reg_storage\[4\]\[24\] _4457_ _4494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput92 pc[5] net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6326_ _2235_ _2236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9045_ _4006_ _4407_ _4451_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6257_ _2168_ _2169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6188_ _2040_ _2101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5208_ reg_file.reg_storage\[4\]\[12\] reg_file.reg_storage\[5\]\[12\] reg_file.reg_storage\[6\]\[12\]
+ reg_file.reg_storage\[7\]\[12\] _1122_ _1123_ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5139_ _1054_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_4_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output115_I net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8829_ _4310_ _4322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_67_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7718__I _3529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6907__A2 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7654__S _3458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8549__I _4126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6069__I _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6843__A1 _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8284__I _3622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8596__A1 reg_file.reg_storage\[12\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5257__S1 _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7628__I _3431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5490_ _1060_ _1070_ _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8520__A1 _4013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4987__I _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7323__A2 net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5334__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7160_ _2973_ _3020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_112_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6111_ _2002_ _2015_ _2024_ _2025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_21_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7091_ _0705_ _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8823__A2 _4313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6834__A1 _1852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6042_ _1955_ _1030_ _1956_ _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7993_ _3502_ _3765_ _3774_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_1_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6944_ _1376_ _2834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_124_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9000__A2 _4405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9663_ _0449_ clknet_leaf_5_clk reg_file.reg_storage\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6875_ _2721_ _2743_ _2766_ _2767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_48_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8614_ _3442_ _4177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9594_ _0380_ clknet_leaf_100_clk reg_file.reg_storage\[9\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5826_ _1741_ _0690_ _1742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_91_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7562__A2 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5757_ reg_file.reg_storage\[8\]\[10\] reg_file.reg_storage\[9\]\[10\] reg_file.reg_storage\[10\]\[10\]
+ reg_file.reg_storage\[11\]\[10\] _1358_ _1672_ _1673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_72_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8545_ reg_file.reg_storage\[12\]\[5\] _3935_ _4132_ _4136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4708_ _0623_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8476_ reg_file.reg_storage\[13\]\[12\] _3953_ _4078_ _4092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8511__A1 reg_file.reg_storage\[13\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5688_ _0690_ _1604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_60_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input76_I pc[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7427_ _3249_ _3259_ net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4639_ reg_file.reg_storage\[1\]\[5\] _0559_ _0557_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7358_ _3195_ _3189_ _3185_ _3196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_9_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ _2216_ _2219_ _1999_ _2220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7078__A1 _2103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7289_ net95 net96 _3112_ _3132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6825__A1 _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9028_ _3983_ _4437_ _4441_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8279__I _3610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7305__A2 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5867__A2 _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7069__A1 _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6816__A1 _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6955__C _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4922__S0 _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5478__S1 _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7241__A1 _3058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4990_ _0784_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_81_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6262__I _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_42_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6660_ _2536_ _2558_ _2559_ _2560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7544__A2 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4989__S0 _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5611_ reg_file.reg_storage\[2\]\[21\] reg_file.reg_storage\[3\]\[21\] _0659_ _1527_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6591_ _1820_ _2494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_27_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_139_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8330_ _3995_ _3996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_121_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5542_ _1386_ _1457_ _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_57_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_100_clk_I clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8261_ _3944_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5473_ reg_file.reg_storage\[4\]\[25\] reg_file.reg_storage\[5\]\[25\] reg_file.reg_storage\[6\]\[25\]
+ reg_file.reg_storage\[7\]\[25\] _1387_ _1388_ _1389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__9049__A2 _4407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8192_ _3667_ _3895_ _3896_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7212_ net76 _1180_ _3062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5402__S1 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5858__A2 _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7143_ _3006_ _1563_ _3010_ _3011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7074_ _2257_ _2550_ _2959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5166__S0 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_115_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7480__A1 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6437__I _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6025_ _1252_ _1086_ _1940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_138_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7976_ _3762_ _3763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6172__I _2085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6927_ _2038_ _2752_ _2818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5794__A1 _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7268__I net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9646_ _0432_ clknet_leaf_61_clk reg_file.reg_storage\[4\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6858_ _1843_ _2706_ _2751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9577_ _0363_ clknet_leaf_52_clk reg_file.reg_storage\[9\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ reg_file.reg_storage\[1\]\[15\] _1724_ _0879_ _1725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8528_ _3912_ _4121_ _4123_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6789_ _2684_ _2671_ _2685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5516__I _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8459_ _3933_ _4075_ _4082_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6649__I1 _2549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4904__S0 _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6347__I _1787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7887__B _3573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7774__A2 _3167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7906__I _3484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5148__S0 _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6257__I _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7797__B net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7214__A1 _3058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7830_ _3431_ _3634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_108_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7088__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7761_ reg_file.reg_storage\[5\]\[11\] _3568_ _3569_ _3570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5776__A1 _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4973_ _0888_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5091__I3 _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9500_ _0286_ clknet_leaf_101_clk reg_file.reg_storage\[8\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6712_ _1635_ _2171_ _2611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7692_ _3392_ _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_9431_ _0217_ clknet_leaf_89_clk reg_file.reg_storage\[13\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6643_ _2251_ _2543_ _2544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5528__A1 _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9362_ _0148_ clknet_leaf_79_clk reg_file.reg_storage\[7\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6574_ _2473_ _2477_ _2478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9293_ _0079_ clknet_leaf_15_clk reg_file.reg_storage\[2\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8313_ _3688_ _3983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8848__S _4315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5525_ _1114_ _1416_ _1440_ _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5336__I _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5456_ _0509_ _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8244_ _3477_ _3932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8647__I _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8175_ _3886_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5387_ reg_file.reg_storage\[2\]\[2\] reg_file.reg_storage\[3\]\[2\] _0628_ _1303_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7126_ net163 _2987_ _2999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input39_I mem_ld_dat[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__I _2080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7057_ _2122_ _2893_ _2943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7453__A1 _3144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6008_ _1921_ _1922_ _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8382__I _4023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7756__A2 _3402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7959_ _3614_ _2977_ _3028_ _3713_ _3748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_83_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9629_ _0415_ clknet_leaf_82_clk reg_file.reg_storage\[1\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7508__A2 _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5298__A3 _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6247__A2 _2157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6798__A3 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9197__A1 _3989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__S0 _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_5_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5357__S _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8668__S _4186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6290_ _1767_ _2175_ _2191_ _2057_ _2193_ _2201_ _2202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_51_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5310_ net95 _0749_ _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5241_ reg_file.reg_storage\[12\]\[14\] reg_file.reg_storage\[13\]\[14\] reg_file.reg_storage\[14\]\[14\]
+ reg_file.reg_storage\[15\]\[14\] _1021_ _1022_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_5172_ net84 _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_8931_ _4383_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 inst[10] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8862_ reg_file.reg_storage\[10\]\[21\] _4336_ _4341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_69_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7813_ _3515_ _3617_ _3618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8793_ _4255_ _4298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5749__A1 _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7744_ _3547_ _3551_ _3553_ _3554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _0858_ _0865_ _0868_ _0869_ _0870_ _0871_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_52_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4887_ _0640_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7546__I net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7675_ _3489_ _3490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9414_ _0200_ clknet_leaf_44_clk reg_file.reg_storage\[13\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6626_ _2509_ _2510_ _2081_ _2527_ _2528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_62_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6557_ _2458_ _2459_ _2460_ _2461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_6_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9345_ _0131_ clknet_leaf_130_clk reg_file.reg_storage\[7\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5508_ reg_file.reg_storage\[4\]\[27\] reg_file.reg_storage\[5\]\[27\] reg_file.reg_storage\[6\]\[27\]
+ reg_file.reg_storage\[7\]\[27\] _1419_ _1423_ _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4575__I2 reg_file.reg_storage\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9276_ _0062_ clknet_leaf_85_clk reg_file.reg_storage\[3\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6488_ _2392_ _2393_ _2371_ _2394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_58_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8227_ _3442_ _3918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5439_ _1354_ _1355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6477__A2 _2381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8158_ reg_file.reg_storage\[6\]\[5\] _3491_ _3873_ _3877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_output145_I net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ _2988_ _2989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8089_ reg_file.reg_storage\[2\]\[11\] _3568_ _3828_ _3834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5532__S0 _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5988__A1 _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5835__S1 _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_67_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5912__A1 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_76_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8287__I _3637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6468__A2 _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5771__S0 _1606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__S0 _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6535__I _2153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_85_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4810_ _0721_ _0718_ _0725_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_56_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5790_ _0727_ _1704_ _1705_ _1115_ _1706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_8_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_64_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _0654_ _0656_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4672_ net12 net1 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7460_ _3286_ _3289_ _3290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4706__A2 _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6411_ _1744_ _2318_ _2319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9130_ reg_file.reg_storage\[4\]\[31\] _4455_ _4503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7391_ _3044_ _3226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6342_ _2116_ _2250_ _2251_ _2252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_116_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9061_ reg_file.reg_storage\[4\]\[1\] _4463_ _4464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ _2021_ _2185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6459__A2 _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8012_ _3611_ _3784_ _3785_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5224_ _0764_ _1137_ _1138_ _1139_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5762__S0 _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5155_ _1060_ _1070_ _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5086_ _0897_ reg_file.reg_storage\[3\]\[29\] _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8914_ reg_file.reg_storage\[9\]\[8\] _4200_ _4372_ _4374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6445__I _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8845_ _4311_ _4331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_67_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8660__I _3596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8776_ reg_file.reg_storage\[11\]\[19\] _4286_ _4289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5988_ _0702_ _0724_ _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7727_ _3024_ _3533_ _3536_ _3537_ _3538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_75_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4939_ _0854_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_47_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8136__A2 _3809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7658_ _3048_ _3080_ _3472_ _3473_ _3474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_133_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6698__A2 _2595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6609_ _2483_ _2486_ _2511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7589_ _3405_ _3408_ _3409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_62_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9328_ _0114_ clknet_leaf_32_clk reg_file.reg_storage\[6\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9259_ _0045_ clknet_leaf_11_clk reg_file.reg_storage\[3\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput191 net191 pc_next[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput180 net180 pc_next[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4720__I2 reg_file.reg_storage\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6870__A2 _2682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4881__A1 _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7895__B _3573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6689__A2 _2588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5370__S _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6265__I _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6960_ _2841_ _2834_ _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5911_ _1744_ _1827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7169__A3 _1900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6891_ _1843_ _2745_ _2741_ _2783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__8480__I _4074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8630_ _4190_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5842_ net19 _1116_ _1480_ _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_33_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5773_ _1684_ _1686_ _1687_ _1688_ _1532_ _1535_ _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_8561_ reg_file.reg_storage\[12\]\[12\] _3953_ _4131_ _4145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8118__A2 _3813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4724_ net8 _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7512_ _3334_ _3336_ _3337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8492_ _4079_ _4101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7877__A1 _3660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4655_ _0568_ _0571_ _0573_ _0574_ _0542_ _0563_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_7443_ net77 net78 _3261_ _3274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xinput60 mem_ld_dat[5] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4586_ _0494_ net231 _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_77_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7374_ _3200_ _3202_ _3207_ _3046_ _3210_ net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_4_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput71 pc[15] net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput82 pc[25] net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9113_ _3986_ _4463_ _4493_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput93 pc[6] net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6325_ _1264_ _2234_ _2235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9044_ reg_file.reg_storage\[1\]\[29\] _4449_ _4451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6256_ _2167_ _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5207_ _0983_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6187_ _2034_ _1910_ _1911_ _2099_ _2100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__8054__A1 _3753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5138_ _1048_ _1051_ _1052_ _1053_ _0822_ _0871_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_input21_I inst[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5069_ reg_file.reg_storage\[4\]\[28\] reg_file.reg_storage\[5\]\[28\] reg_file.reg_storage\[6\]\[28\]
+ reg_file.reg_storage\[7\]\[28\] _0780_ _0984_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_clkbuf_4_13_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output108_I net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8828_ _4195_ _4312_ _4321_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5415__I0 reg_file.reg_storage\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8759_ reg_file.reg_storage\[11\]\[12\] _4209_ _4265_ _4279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8109__A2 _3844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5040__A1 _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5591__A2 _1506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7868__A1 _3660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5343__A2 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8766__S _4265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8565__I _4127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7909__I _3704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8006__S _3768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7020__A2 _2537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_1_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6110_ _2017_ _2023_ _2024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7090_ net97 _2973_ _2974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_119_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _1147_ _1042_ _1956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8036__A1 _3710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8587__A2 _4129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7992_ reg_file.reg_storage\[3\]\[6\] _3766_ _3774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6598__A1 _2018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6943_ _2786_ _2830_ _2832_ _2833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7819__I _3623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9662_ _0448_ clknet_leaf_84_clk reg_file.reg_storage\[15\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6874_ _1555_ _2672_ _2766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5825_ _1736_ _1738_ _1739_ _1740_ _1531_ _1235_ _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_8613_ _4170_ _4174_ _4176_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9593_ _0379_ clknet_leaf_101_clk reg_file.reg_storage\[9\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5756_ _1627_ _1672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_97_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8544_ _3933_ _4128_ _4135_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8475_ _4091_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4707_ net8 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5687_ _0914_ _1380_ _1581_ _1603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_142_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7426_ _3250_ _3252_ _3258_ _3053_ _3259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4638_ reg_file.reg_storage\[2\]\[5\] reg_file.reg_storage\[3\]\[5\] _0503_ _0559_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_142_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input69_I pc[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5074__I _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4569_ net13 _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_9_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7357_ _3180_ _3184_ _3195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_9_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5708__S0 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6308_ _2217_ _1966_ _2218_ _2045_ _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_7288_ _3121_ _3123_ _3131_ net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_31_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_9027_ reg_file.reg_storage\[1\]\[22\] _4410_ _4441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6239_ _2094_ _2149_ _2150_ _2151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8578__A2 _4152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7250__A2 _3089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5403__I3 reg_file.reg_storage\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8502__A2 _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7305__A3 _3138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5316__A2 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5867__A3 _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8295__I _3656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__A1 _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4922__S1 _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7241__A2 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7639__I _3426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5610_ reg_file.reg_storage\[8\]\[21\] reg_file.reg_storage\[9\]\[21\] reg_file.reg_storage\[10\]\[21\]
+ reg_file.reg_storage\[11\]\[21\] _1368_ _1425_ _1526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6590_ _2212_ _2328_ _2491_ _2492_ _2493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_73_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8741__A2 _4263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_140_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_139_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5541_ _1445_ _1456_ _1457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_6_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4998__I _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8260_ reg_file.reg_storage\[7\]\[8\] _3943_ _3941_ _3944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_81_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5472_ _1363_ _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_112_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6504__A1 _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7211_ _3060_ _3061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8191_ reg_file.reg_storage\[6\]\[19\] _3893_ _3896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7142_ _2985_ _3010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6718__I _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7073_ _2002_ _2756_ _2957_ _2958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5166__S1 _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _1938_ _1295_ _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7480__A2 _1881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7975_ _3760_ _3387_ _3761_ _3762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_85_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _2798_ _2107_ _2816_ _2817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_92_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _2634_ _2549_ _2750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9645_ _0431_ clknet_leaf_13_clk reg_file.reg_storage\[4\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9576_ _0362_ clknet_leaf_53_clk reg_file.reg_storage\[9\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6788_ _1849_ _2684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5808_ reg_file.reg_storage\[2\]\[15\] reg_file.reg_storage\[3\]\[15\] _1587_ _1724_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_33_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8527_ reg_file.reg_storage\[12\]\[0\] _4122_ _4123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5739_ net30 _0716_ _1653_ _1654_ _1652_ _1655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_17_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8458_ reg_file.reg_storage\[13\]\[4\] _4076_ _4082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8389_ _3946_ _4025_ _4039_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output175_I net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7409_ _3230_ _3241_ _3242_ _3243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4809__A1 _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4904__S1 _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5482__A1 _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5609__I0 _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7931__B1 _3496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5707__I _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__S _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_1_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5442__I _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5148__S1 _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7462__A2 _3285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7214__A2 _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7760_ _3457_ _3569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_47_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4972_ _0748_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_121_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6711_ _2067_ _2610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_59_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7691_ _3466_ _3504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_144_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9430_ _0216_ clknet_leaf_87_clk reg_file.reg_storage\[13\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8714__A2 _4241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6642_ _2290_ _2285_ _2059_ _2543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5528__A2 _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5084__S0 _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9361_ _0147_ clknet_leaf_70_clk reg_file.reg_storage\[7\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_80_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8312_ _3981_ _3975_ _3982_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5617__I _1532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _1132_ _1818_ _2266_ _2476_ _2477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_54_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9292_ _0078_ clknet_leaf_58_clk reg_file.reg_storage\[2\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5524_ _0493_ _1417_ _1439_ _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_42_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7150__A1 _3014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5455_ reg_file.reg_storage\[8\]\[26\] reg_file.reg_storage\[9\]\[26\] reg_file.reg_storage\[10\]\[26\]
+ reg_file.reg_storage\[11\]\[26\] _1360_ _1364_ _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8243_ _3931_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8174_ reg_file.reg_storage\[6\]\[12\] _3585_ _3872_ _3886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7125_ _1717_ _2995_ _2998_ net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_112_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5386_ reg_file.reg_storage\[8\]\[2\] reg_file.reg_storage\[9\]\[2\] reg_file.reg_storage\[10\]\[2\]
+ reg_file.reg_storage\[11\]\[2\] _0809_ _1301_ _1302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5352__I _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_105_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7056_ _2905_ _2107_ _2030_ _2942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8663__I _3610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6007_ _1010_ _0831_ _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7958_ _3722_ _3746_ _3747_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6964__A1 _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6909_ _2799_ _2168_ _2800_ _2801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7889_ _3671_ _3285_ _3499_ _3686_ _3687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_119_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9628_ _0414_ clknet_leaf_83_clk reg_file.reg_storage\[1\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5075__S0 _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9559_ _0345_ clknet_leaf_105_clk reg_file.reg_storage\[10\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7141__A1 _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_41_clk_I clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6358__I _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4889__S0 _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__S1 _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_56_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6093__I _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8944__A2 _4386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_134_clk clknet_4_4_0_clk clknet_leaf_134_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6707__A1 _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_114_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5240_ _0899_ _1153_ _1154_ _1155_ _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7652__I _3468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_129_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5171_ _1085_ _1086_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5172__I net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7435__A2 _3253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8930_ reg_file.reg_storage\[9\]\[15\] _4216_ _4365_ _4383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__9188__A2 _4536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 inst[11] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8861_ _4228_ _4338_ _4340_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_69_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7812_ _3522_ _3615_ _3616_ _3617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8935__A2 _4381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8792_ _4240_ _4256_ _4297_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5749__A2 _1664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7743_ _3485_ _3146_ _3552_ _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4955_ _0824_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4886_ _0801_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7674_ _3480_ _3460_ _3483_ _3488_ _3489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_9413_ _0199_ clknet_leaf_39_clk reg_file.reg_storage\[13\]\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6625_ _2509_ _2510_ _2374_ _2527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6556_ _2396_ _2445_ _2447_ _2448_ _2460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_9344_ _0130_ clknet_leaf_134_clk reg_file.reg_storage\[7\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9275_ _0061_ clknet_leaf_84_clk reg_file.reg_storage\[3\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5507_ _1422_ _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4575__I3 reg_file.reg_storage\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9112__A2 _4461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8226_ _3912_ _3915_ _3917_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7123__A1 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6487_ _2318_ _2353_ _1753_ _2393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input51_I mem_ld_dat[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5438_ _0593_ _0746_ _0706_ _0657_ _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8157_ _3478_ _3869_ _3876_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5369_ reg_file.reg_storage\[2\]\[4\] reg_file.reg_storage\[3\]\[4\] _0809_ _1285_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7108_ _2987_ _2988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8088_ _3833_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7426__A2 _3252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5780__S1 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6906__I _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7039_ _2925_ net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4627__S _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output138_I net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9179__A2 _4531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5532__S1 _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5988__A2 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6937__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5296__S0 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7737__I _3546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_116_clk clknet_4_12_0_clk clknet_leaf_116_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5912__A2 _1751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5220__S0 _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5771__S1 _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__S1 _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8917__A2 _4375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6928__A1 _2036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5287__S0 _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_107_clk clknet_4_13_0_clk clknet_leaf_107_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4740_ _0614_ _0602_ _0603_ _0655_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_113_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4671_ net29 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7390_ _3179_ _3212_ _3225_ net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6410_ _2155_ _2232_ net217 _2152_ _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_98_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6341_ _1787_ _2251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7105__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_116_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9060_ _4459_ _4463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6272_ _1232_ _1298_ _2183_ _2184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8011_ reg_file.reg_storage\[3\]\[14\] _3778_ _3785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5223_ _0772_ reg_file.reg_storage\[2\]\[13\] _0806_ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5211__S0 _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8605__A1 _4013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5762__S1 _1596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5831__S _1605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5154_ _0937_ _0938_ _1069_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7408__A2 _3228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8456__I1 _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5085_ reg_file.reg_storage\[1\]\[29\] _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8913_ _4373_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6919__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8844_ _4330_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5987_ _0696_ _1902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8775_ _4266_ _4288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7726_ _3521_ _3537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4938_ _0638_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4869_ _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_62_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7344__A1 _2969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7657_ _3081_ _3403_ _3473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6608_ _1720_ _2510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7588_ net40 net49 _3407_ _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9327_ _0113_ clknet_leaf_57_clk reg_file.reg_storage\[6\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6539_ _1132_ _2442_ _2443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_31_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9258_ _0044_ clknet_leaf_14_clk reg_file.reg_storage\[3\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput170 net170 mem_st_mask[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8209_ reg_file.reg_storage\[6\]\[27\] _3903_ _3906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9189_ _3977_ _4538_ _4540_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput192 net192 pc_next[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput181 net181 pc_next[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4720__I3 reg_file.reg_storage\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6636__I _2398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5188__S _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_133_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6320__B _1759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5649__A1 _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6074__A1 _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5910_ _1825_ _1667_ _1826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6890_ _2778_ _2746_ _2782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_76_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5841_ _1309_ _1240_ _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_124_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8560_ _4144_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6281__I _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5772_ reg_file.reg_storage\[4\]\[12\] reg_file.reg_storage\[5\]\[12\] reg_file.reg_storage\[6\]\[12\]
+ reg_file.reg_storage\[7\]\[12\] _1606_ _1608_ _1688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_8_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8491_ _3970_ _4094_ _4100_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4723_ reg_file.reg_storage\[2\]\[0\] reg_file.reg_storage\[3\]\[0\] _0638_ _0639_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7511_ net84 _3335_ _3336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7442_ _3200_ _3262_ _3269_ _3271_ _3273_ net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_17_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4654_ reg_file.reg_storage\[4\]\[6\] reg_file.reg_storage\[5\]\[6\] reg_file.reg_storage\[6\]\[6\]
+ reg_file.reg_storage\[7\]\[6\] _0572_ _0570_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_4_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5888__A1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput61 mem_ld_dat[6] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput50 mem_ld_dat[25] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4585_ _0501_ _0505_ _0506_ _0507_ _0509_ _0510_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_52_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7373_ _3209_ net103 _3210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput72 pc[16] net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9112_ reg_file.reg_storage\[4\]\[23\] _4461_ _4493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput94 pc[7] net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput83 pc[26] net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4560__A1 _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6324_ _2231_ _2233_ _2234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_9043_ _4003_ _4445_ _4450_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8936__I _4360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6255_ _1784_ _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5206_ _0854_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6186_ _2097_ _1918_ _2099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8054__A2 _3809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5137_ reg_file.reg_storage\[8\]\[24\] reg_file.reg_storage\[9\]\[24\] reg_file.reg_storage\[10\]\[24\]
+ reg_file.reg_storage\[11\]\[24\] _0767_ _1047_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_4_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5068_ _0983_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_4_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6065__A1 _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input14_I inst[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8827_ reg_file.reg_storage\[10\]\[6\] _4313_ _4321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8758_ _4278_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7709_ _2976_ _2981_ _3521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8689_ _4230_ _4226_ _4231_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__A1 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5879__B2 _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8293__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8045__A2 _3799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7556__A1 _3144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7197__I _3047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_61_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7308__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5445__I _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__S0 _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8808__A1 reg_file.reg_storage\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6531__A2 _2431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6040_ _1162_ _1955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_0_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I inst[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7991_ _3773_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _2810_ _2831_ _2832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_124_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9661_ _0447_ clknet_leaf_115_clk reg_file.reg_storage\[4\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6873_ _2765_ net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_48_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5824_ reg_file.reg_storage\[4\]\[8\] reg_file.reg_storage\[5\]\[8\] reg_file.reg_storage\[6\]\[8\]
+ reg_file.reg_storage\[7\]\[8\] _1605_ _0578_ _1740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8612_ reg_file.reg_storage\[8\]\[0\] _4175_ _4176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9592_ _0378_ clknet_leaf_107_clk reg_file.reg_storage\[9\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6770__A2 _2651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7562__A4 _3356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8543_ reg_file.reg_storage\[12\]\[4\] _4129_ _4135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5755_ _0722_ _1355_ _1671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_127_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8474_ reg_file.reg_storage\[13\]\[11\] _3951_ _4085_ _4091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5686_ _1580_ _1601_ _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4706_ _0606_ _0621_ _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_115_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7056__B _2030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5355__I _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7425_ _3254_ _3257_ _3258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4637_ reg_file.reg_storage\[8\]\[5\] reg_file.reg_storage\[9\]\[5\] reg_file.reg_storage\[10\]\[5\]
+ reg_file.reg_storage\[11\]\[5\] _0556_ _0557_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_130_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4568_ _0493_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7356_ _3192_ _3193_ _3194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5708__S1 _1623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7570__I net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7287_ _3100_ net127 _3101_ _3130_ _3131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6307_ _2052_ _1943_ _2218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9026_ _3980_ _4437_ _4440_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6238_ _1777_ _2089_ _2150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8027__A2 _3789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6169_ _2075_ _2078_ _2082_ _2064_ _1947_ _2083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
Xclkbuf_leaf_96_clk clknet_4_15_0_clk clknet_leaf_96_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6038__A1 _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output120_I net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6761__A2 _2604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20_clk clknet_4_7_0_clk clknet_leaf_20_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_133_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6513__A2 _2405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8266__A2 _3923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8018__A2 _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4827__A2 _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_87_clk clknet_4_14_0_clk clknet_leaf_87_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_128_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7616__I2 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7241__A3 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5635__S0 _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6752__A2 _2439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_139_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5540_ _1448_ _1452_ _1453_ _1454_ _1455_ _1395_ _1456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_54_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_clk clknet_4_0_0_clk clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ _1359_ _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7701__A1 _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7210_ _3052_ _3060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8190_ _3873_ _3895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7141_ _1645_ _3000_ _3009_ net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_10_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7072_ _2360_ _2955_ _2956_ _2027_ _2957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6268__A1 _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6023_ _1265_ _1938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_78_clk clknet_4_12_0_clk clknet_leaf_78_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5491__A2 _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7974_ _3389_ _3390_ _3394_ _3761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_6925_ _1071_ _2363_ _2816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9644_ _0430_ clknet_leaf_62_clk reg_file.reg_storage\[4\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6856_ _2725_ _2748_ _2749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6787_ _2182_ _2682_ _2683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_9575_ _0361_ clknet_leaf_26_clk reg_file.reg_storage\[9\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5807_ reg_file.reg_storage\[8\]\[15\] reg_file.reg_storage\[9\]\[15\] reg_file.reg_storage\[10\]\[15\]
+ reg_file.reg_storage\[11\]\[15\] _1615_ _0879_ _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_17_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8526_ _4119_ _4122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5738_ _1431_ _0716_ _1654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input81_I pc[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8496__A2 _4101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5669_ _0806_ _1582_ _1584_ _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_44_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8457_ _4081_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8388_ reg_file.reg_storage\[14\]\[9\] _4038_ _4039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7408_ _3227_ _3228_ _3242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7339_ _3121_ _3167_ _3178_ net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9009_ reg_file.reg_storage\[1\]\[14\] _4424_ _4431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4809__A2 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5482__A2 _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9020__I _4415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8420__A2 _4026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6982__A2 _2431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_0_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8184__A1 _3638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5196__S _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7931__B2 _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8487__A2 _4088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7695__B1 _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_0_clk clknet_4_4_0_clk clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8411__A2 _4049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _0833_ _0877_ _0886_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_121_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4984__A1 _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6710_ _2407_ _2361_ _2602_ _2608_ _2609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_58_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7690_ _3428_ _3502_ _3503_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6641_ _2103_ _2158_ _2542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_144_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5084__S1 _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9360_ _0146_ clknet_leaf_33_clk reg_file.reg_storage\[7\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7922__A1 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__I _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5119__B _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8311_ reg_file.reg_storage\[7\]\[21\] _3971_ _3982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6572_ _2474_ _2268_ _2475_ _2476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5523_ _1424_ _1434_ _1435_ _1436_ _1437_ _1438_ _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_81_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9291_ _0077_ clknet_leaf_11_clk reg_file.reg_storage\[2\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5454_ reg_file.reg_storage\[12\]\[26\] reg_file.reg_storage\[13\]\[26\] reg_file.reg_storage\[14\]\[26\]
+ reg_file.reg_storage\[15\]\[26\] _1369_ _1364_ _1370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_112_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8242_ reg_file.reg_storage\[7\]\[3\] _3930_ _3928_ _3931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6489__B2 _1734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8173_ _3885_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5161__A1 _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5385_ _0759_ _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7124_ net162 _2987_ _2998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8650__A2 _4182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7055_ _2010_ _2843_ _2941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6006_ _1041_ _0910_ _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6413__A1 _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7957_ reg_file.reg_storage\[5\]\[30\] _3399_ _3747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6908_ _2799_ _2496_ _2800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7888_ _3299_ _3464_ _3686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9627_ _0413_ clknet_leaf_83_clk reg_file.reg_storage\[1\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6839_ _2000_ _2265_ _2731_ _2732_ _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_134_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5075__S1 _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7295__I _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7913__B2 _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9558_ _0344_ clknet_leaf_113_clk reg_file.reg_storage\[10\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8509_ _3996_ _4069_ _4110_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9489_ _0275_ clknet_leaf_67_clk reg_file.reg_storage\[8\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8854__I _4310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4889__S1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6707__A2 _2604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5915__B1 _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7380__A2 _3184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7933__I _3725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__A1 _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8880__A2 _4346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6891__A1 _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5170_ _0795_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput4 inst[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_36_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8860_ reg_file.reg_storage\[10\]\[20\] _4336_ _4340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_69_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7811_ net39 _3517_ _3481_ _3616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_8791_ reg_file.reg_storage\[11\]\[26\] _4296_ _4297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4954_ _0821_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_86_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4957__A1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7742_ _1671_ _3402_ _3416_ _3552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_144_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _0638_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_9412_ _0198_ clknet_leaf_16_clk reg_file.reg_storage\[13\]\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5628__I _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7673_ _3090_ _3403_ _3487_ _3488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_35_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6624_ _2264_ _2525_ _2001_ _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8939__I _4366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9343_ _0129_ clknet_leaf_6_clk reg_file.reg_storage\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6555_ _2391_ _2445_ _2459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9274_ _0060_ clknet_leaf_86_clk reg_file.reg_storage\[3\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5506_ _1421_ _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8225_ reg_file.reg_storage\[7\]\[0\] _3916_ _3917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_rebuffer17_I _1493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6486_ _1753_ _2318_ _2353_ _2392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_112_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5437_ _1352_ _1353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input44_I mem_ld_dat[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8156_ reg_file.reg_storage\[6\]\[4\] _3870_ _3876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5368_ reg_file.reg_storage\[4\]\[4\] reg_file.reg_storage\[5\]\[4\] reg_file.reg_storage\[6\]\[4\]
+ reg_file.reg_storage\[7\]\[4\] _1020_ _1141_ _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7107_ _2986_ _2987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8087_ reg_file.reg_storage\[2\]\[10\] _3557_ _3828_ _3833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5299_ _1207_ _1214_ _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7038_ _2352_ _2911_ _2916_ _2924_ _2925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4707__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6937__A2 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6398__B1 _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8989_ _4419_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5296__S1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4948__A1 _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7898__B1 _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7362__A2 _3194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8862__A2 _4336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5220__S1 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6625__A1 _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4731__S0 _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9330__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5287__S1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4670_ net28 _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7353__A2 _3182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6340_ _2048_ _2020_ _2063_ _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8853__A2 _4331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5183__I _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6271_ _2040_ _2183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8010_ _3764_ _3784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5222_ _1061_ reg_file.reg_storage\[3\]\[13\] _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5211__S1 _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5667__A2 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _1064_ _1066_ _1067_ _1068_ _0870_ _1025_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_5084_ reg_file.reg_storage\[4\]\[29\] reg_file.reg_storage\[5\]\[29\] reg_file.reg_storage\[6\]\[29\]
+ reg_file.reg_storage\[7\]\[29\] _0999_ _0903_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_142_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8912_ reg_file.reg_storage\[9\]\[7\] _4197_ _4372_ _4373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__9030__A2 _4412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8843_ reg_file.reg_storage\[10\]\[13\] _4211_ _4315_ _4330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5986_ _1901_ net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8774_ _4222_ _4281_ _4287_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7725_ _3410_ _3535_ _3536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4937_ net80 _0852_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_40_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4868_ _0625_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7656_ _3430_ _3472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_144_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6607_ _1955_ _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7587_ _3406_ _3407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_9326_ _0112_ clknet_leaf_57_clk reg_file.reg_storage\[6\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5294__S _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4799_ _0673_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_132_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9097__A2 _4481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_55_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6538_ _1818_ _2441_ _2442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9257_ _0043_ clknet_leaf_44_clk reg_file.reg_storage\[3\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6469_ _2371_ _1830_ _2373_ _2375_ _2376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xoutput160 net160 mem_st_dat[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_112_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8208_ _3861_ _3905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9188_ reg_file.reg_storage\[15\]\[20\] _4536_ _4540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output150_I net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8139_ _3860_ _3863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput171 net171 pc_next[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput182 net182 pc_next[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput193 net193 pc_next[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4638__S _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_113_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9021__A2 _4435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_128_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5594__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__A2 _1812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7099__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8835__A2 _4325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5649__A2 _1564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4952__S0 _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5121__I1 reg_file.reg_storage\[13\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6074__A2 _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9012__A2 _4406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5840_ _1668_ _1683_ _1733_ _1755_ _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_9_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5585__A1 _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5771_ reg_file.reg_storage\[12\]\[12\] reg_file.reg_storage\[13\]\[12\] reg_file.reg_storage\[14\]\[12\]
+ reg_file.reg_storage\[15\]\[12\] _1606_ _0878_ _1687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8490_ reg_file.reg_storage\[13\]\[18\] _4099_ _4100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7510_ _1414_ _1415_ _3335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4722_ _0637_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_118_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8523__A1 _4015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8489__I _4073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6129__A3 _2042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7441_ _3272_ net109 _3273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8374__I1 _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput40 mem_ld_dat[16] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4653_ reg_file.reg_storage\[12\]\[6\] reg_file.reg_storage\[13\]\[6\] reg_file.reg_storage\[14\]\[6\]
+ reg_file.reg_storage\[15\]\[6\] _0572_ _0570_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_4_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput62 mem_ld_dat[7] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput51 mem_ld_dat[26] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7372_ _3208_ _3209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput73 pc[17] net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4584_ net16 _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5888__A2 _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9111_ _3983_ _4488_ _4492_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput95 pc[8] net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput84 pc[27] net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4560__A2 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6323_ _2155_ _2232_ _2152_ _2233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9042_ reg_file.reg_storage\[1\]\[28\] _4449_ _4450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6254_ _2151_ _2163_ _2165_ _2166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_90_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5205_ net68 _0852_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6185_ _1915_ _1928_ _2097_ _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5136_ reg_file.reg_storage\[12\]\[24\] reg_file.reg_storage\[13\]\[24\] reg_file.reg_storage\[14\]\[24\]
+ reg_file.reg_storage\[15\]\[24\] _0802_ _0804_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5067_ _0759_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_4_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7565__A2 net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8826_ _4320_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8757_ reg_file.reg_storage\[11\]\[11\] _4207_ _4272_ _4278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5969_ _1880_ _1884_ _1377_ _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_23_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7708_ _3517_ _3519_ _3520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8688_ reg_file.reg_storage\[8\]\[21\] _4223_ _4231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7639_ _3426_ _3457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9309_ _0095_ clknet_4_12_0_clk reg_file.reg_storage\[2\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5803__A2 _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7556__A2 _3370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8505__A1 reg_file.reg_storage\[13\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7308__A2 _1671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5726__I _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__S1 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5178__S0 _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8772__I _4260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6047__A2 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7990_ reg_file.reg_storage\[3\]\[5\] _3491_ _3769_ _3773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6941_ _2805_ _2811_ _2831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9660_ _0446_ clknet_leaf_94_clk reg_file.reg_storage\[4\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6872_ _2747_ _2749_ _2764_ _2765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4805__I _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8611_ _4172_ _4175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5823_ reg_file.reg_storage\[12\]\[8\] reg_file.reg_storage\[13\]\[8\] reg_file.reg_storage\[14\]\[8\]
+ reg_file.reg_storage\[15\]\[8\] _0577_ _0578_ _1739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_9591_ _0377_ clknet_leaf_107_clk reg_file.reg_storage\[9\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7547__A2 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8542_ _4134_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5754_ _0734_ _1670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8473_ _4090_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5685_ _1600_ _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4705_ _0620_ _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_115_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7424_ _3238_ _3245_ _3256_ _3257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4636_ _0483_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_130_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5730__A1 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7355_ _1134_ _3181_ _3193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4567_ _0492_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6306_ _2062_ _2217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_9_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7286_ _3127_ _3129_ _3130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9025_ reg_file.reg_storage\[1\]\[21\] _4435_ _4440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6467__I _2076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6237_ _2093_ _2091_ _2149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6168_ _1947_ _2079_ _2081_ _2082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5119_ _0773_ reg_file.reg_storage\[2\]\[30\] _0775_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_99_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6099_ _2012_ _1044_ _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output113_I net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8809_ _4170_ _4306_ _4308_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7538__A2 _3346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4651__S _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5546__I _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5721__A1 _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8857__I _4316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8592__I _4119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7616__I3 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8974__A1 _3760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5332__S0 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8726__A1 reg_file.reg_storage\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7936__I _3417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6588__I0 _2215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5635__S1 _1537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5456__I _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5960__A1 _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5470_ _1385_ _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7701__A2 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7140_ net159 _3004_ _3009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7071_ _2217_ _2866_ _2956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6022_ _1936_ _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7973_ _0975_ _3760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_55_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6924_ _2404_ _2814_ _2815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8717__A1 reg_file.reg_storage\[8\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9643_ _0429_ clknet_leaf_9_clk reg_file.reg_storage\[4\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7846__I _3648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8193__A2 _3893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6855_ _2741_ _2726_ _2746_ _2748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9574_ _0360_ clknet_leaf_45_clk reg_file.reg_storage\[9\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6786_ _2681_ _2682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5806_ _0863_ _1704_ _1584_ _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_45_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8525_ _4120_ _4121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_135_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7067__B _2537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7940__A2 _3357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5737_ _0747_ _0684_ _1410_ _1653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_134_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8456_ reg_file.reg_storage\[13\]\[3\] _3930_ _4079_ _4081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5668_ _1583_ _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input74_I pc[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7407_ _3227_ _3228_ _3241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5599_ _1468_ _0986_ _1513_ _1514_ _1515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8677__I _4180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8387_ _4023_ _4038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5703__A1 _1604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4619_ _0521_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_103_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7338_ _3157_ net100 _3158_ _3177_ _3178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7269_ _3097_ _3098_ _3113_ _3114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7456__A1 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9008_ _4410_ _4430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_67_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8184__A2 _3888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6195__A1 _2103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4745__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7695__B2 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7695__A1 _3116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6670__A2 _2258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4970_ _0885_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_129_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5387__S _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6640_ _2532_ _2536_ _2540_ _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6186__A1 _2097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6571_ _2474_ _2269_ _2475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7922__A2 _3403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8310_ _3980_ _3981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_80_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5522_ _1105_ _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_143_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9290_ _0076_ clknet_leaf_15_clk reg_file.reg_storage\[2\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5453_ _1368_ _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_42_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8241_ _3468_ _3930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8172_ reg_file.reg_storage\[6\]\[11\] _3568_ _3879_ _3885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5384_ net87 _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7123_ _1702_ _2995_ _2997_ net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7989__A2 _3765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7054_ _2926_ _1874_ _2075_ _2939_ _2940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6005_ _1913_ _1919_ _1240_ _1920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7956_ _3745_ _3746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7887_ _3632_ _3684_ _3573_ _3685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6907_ _2797_ _2798_ _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9626_ _0412_ clknet_4_14_0_clk reg_file.reg_storage\[1\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6838_ _2634_ _2525_ _2210_ _2732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9557_ _0343_ clknet_leaf_119_clk reg_file.reg_storage\[10\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8508_ reg_file.reg_storage\[13\]\[26\] _4109_ _4110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9115__A1 _3989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _0949_ _2629_ _2651_ _2644_ _2665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_9488_ _0274_ clknet_leaf_68_clk reg_file.reg_storage\[8\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8401__S _4028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_28_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8439_ _3397_ _4015_ _4067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output180_I net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7429__A1 _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_37_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6404__A2 _2277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6604__B _2499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6168__A1 _1947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8157__A2 _3869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_46_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5915__B2 _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5915__A1 _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 inst[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7810_ _3614_ _3433_ _3461_ _3615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_69_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8790_ _4254_ _4296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7741_ _3514_ _3550_ _3551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_82_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4953_ reg_file.reg_storage\[8\]\[23\] reg_file.reg_storage\[9\]\[23\] reg_file.reg_storage\[10\]\[23\]
+ reg_file.reg_storage\[11\]\[23\] _0866_ _0867_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_143_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8148__A2 _3870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7672_ _3485_ _3089_ _3486_ _3487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4884_ _0753_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6623_ _2383_ _2524_ _2052_ _2525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9411_ _0197_ clknet_leaf_135_clk reg_file.reg_storage\[13\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9342_ _0128_ clknet_leaf_88_clk reg_file.reg_storage\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _2454_ _2455_ _2456_ _2457_ _2458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_113_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9273_ _0059_ clknet_leaf_85_clk reg_file.reg_storage\[3\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5505_ _1420_ _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6485_ _2320_ _2355_ _2391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8224_ _3913_ _3916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8320__A2 _3924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5436_ net25 _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8155_ _3875_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5367_ _1281_ _1282_ _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7106_ _2985_ _2982_ _2986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8086_ _3543_ _3818_ _3832_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5298_ _0621_ _0938_ _1213_ _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input37_I mem_ld_dat[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7037_ _2421_ _2505_ _2923_ _2610_ _2924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7831__A1 _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4924__S _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__A1 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8988_ reg_file.reg_storage\[1\]\[5\] _3490_ _4415_ _4419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4948__A2 reg_file.reg_storage\[2\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7939_ _3346_ _3505_ _3731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9609_ _0395_ clknet_leaf_50_clk reg_file.reg_storage\[1\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7898__A1 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7898__B2 _3694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6570__A1 _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8311__A2 _3971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6322__A1 _1765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5508__S0 _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7822__A1 _3010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6625__A2 _2510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4731__S1 _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7105__A3 _2972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5464__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5747__S0 _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6270_ _2177_ _2178_ _2181_ _2182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_11_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5221_ reg_file.reg_storage\[1\]\[13\] _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4875__A1 _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8775__I _4266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5667__A3 _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5152_ reg_file.reg_storage\[8\]\[25\] reg_file.reg_storage\[9\]\[25\] reg_file.reg_storage\[10\]\[25\]
+ reg_file.reg_storage\[11\]\[25\] _0855_ _1063_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__6616__A2 _2461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6509__B _2157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5083_ _0817_ _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8911_ _4360_ _4372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_2_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8369__A2 _4025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8842_ _4329_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8773_ reg_file.reg_storage\[11\]\[18\] _4286_ _4287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7041__A2 _2537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7724_ _3534_ _3032_ net50 _3535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5985_ _1900_ _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5052__A1 _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9169__I1 _3584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4936_ _0749_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4867_ reg_file.reg_storage\[8\]\[20\] reg_file.reg_storage\[9\]\[20\] reg_file.reg_storage\[10\]\[20\]
+ reg_file.reg_storage\[11\]\[20\] _0758_ _0781_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_7_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7655_ _3471_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7586_ _3026_ _3406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6606_ _2508_ net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_28_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9325_ _0111_ clknet_leaf_13_clk reg_file.reg_storage\[6\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6537_ _2439_ _2440_ _2441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4798_ net5 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5374__I _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9256_ _0042_ clknet_leaf_45_clk reg_file.reg_storage\[3\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6468_ _2371_ _1830_ _2374_ _2375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput161 net161 mem_st_dat[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput150 net150 mem_st_dat[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_140_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8207_ _3719_ _3862_ _3904_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9187_ _3973_ _4538_ _4539_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6399_ _2068_ _2302_ _2307_ _2308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5419_ _1334_ _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7803__B _3446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8138_ _3861_ _3862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput194 net194 pc_next[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput172 net172 pc_next[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput183 net183 pc_next[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_output143_I net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7804__A1 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4718__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7804__B2 _3609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8069_ reg_file.reg_storage\[2\]\[2\] _3456_ _3822_ _3823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7280__A2 _3116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5291__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5043__A1 _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8780__A2 _4286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7764__I _3484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6543__A1 _1959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7886__A4 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8048__A1 _3746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4952__S1 _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4609__A1 _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5282__A1 _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8771__A2 _4281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5770_ reg_file.reg_storage\[1\]\[12\] _1685_ _1608_ _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4721_ _0627_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8523__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4652_ _0503_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7440_ _3208_ _3272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7731__B1 _3540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput30 inst[7] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_25_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput63 mem_ld_dat[8] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 mem_ld_dat[17] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput52 mem_ld_dat[27] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9110_ reg_file.reg_storage\[4\]\[22\] _4461_ _4492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4583_ _0508_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7371_ _3049_ _3208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4640__S0 _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5194__I _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput96 pc[9] net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput74 pc[18] net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput85 pc[28] net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4560__A3 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6322_ _1765_ _1763_ _2232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
X_9041_ _4404_ _4449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6837__A2 _2730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6253_ _2086_ _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8039__A1 _3719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5922__I _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5204_ _1119_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6184_ _1971_ _2097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5135_ reg_file.reg_storage\[1\]\[24\] _1050_ _1047_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5066_ net85 _0750_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8825_ reg_file.reg_storage\[10\]\[5\] _4193_ _4316_ _4320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8756_ _4277_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5968_ _1399_ _1407_ _1883_ _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7707_ _3518_ _3032_ net49 _3519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_81_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4919_ _0834_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_23_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8687_ _3681_ _4230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5899_ _1703_ _1706_ _1815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7638_ _3455_ _3456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7569_ net31 _3389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_62_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9308_ _0094_ clknet_leaf_85_clk reg_file.reg_storage\[2\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9239_ _0025_ clknet_leaf_114_clk reg_file.reg_storage\[5\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4649__S _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8202__A1 _3705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5016__A1 _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8753__A2 _4275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6764__A1 _2463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6819__A2 _1542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5178__S1 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7244__A2 _3081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _2769_ _2810_ _2811_ _2830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6452__B1 _2358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_54_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6871_ _2583_ _2758_ _2763_ _2764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5189__I _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8610_ _4173_ _4174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5822_ reg_file.reg_storage\[1\]\[8\] _1737_ _1361_ _1738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9590_ _0376_ clknet_leaf_110_clk reg_file.reg_storage\[9\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6755__A1 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7547__A3 _3356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5753_ _1195_ _1204_ _1669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8541_ reg_file.reg_storage\[12\]\[3\] _3930_ _4132_ _4134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4704_ _0619_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4821__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8472_ reg_file.reg_storage\[13\]\[10\] _3949_ _4085_ _4090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5684_ _0670_ _1585_ _1599_ _1600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7180__A1 _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_112_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7423_ net74 _3255_ _3256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4635_ _0496_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_115_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _0491_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_53_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7354_ net70 _3192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4613__S0 _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5730__A2 _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6305_ _2214_ _2215_ _2216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9024_ _3977_ _4437_ _4439_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7285_ _3122_ _3128_ _3129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_clkbuf_leaf_127_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6236_ _2148_ net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__5494__A1 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6167_ _2080_ _2081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5118_ _0897_ reg_file.reg_storage\[3\]\[30\] _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6098_ _2011_ _2012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5049_ _0964_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_95_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output106_I net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8808_ reg_file.reg_storage\[10\]\[0\] _4307_ _4308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8739_ reg_file.reg_storage\[11\]\[3\] _4189_ _4266_ _4268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9034__I _4405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7474__A2 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8423__A1 reg_file.reg_storage\[14\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7226__A2 _3068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4906__I _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5332__S1 _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6588__I1 _2211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9151__A2 _4513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7162__B2 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8984__S _4415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7070_ _2036_ _2918_ _2954_ _2955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6021_ _1281_ _1295_ _1936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7972_ _3421_ _3757_ _3759_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _2805_ _2806_ _2812_ _2814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_85_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9642_ _0428_ clknet_leaf_11_clk reg_file.reg_storage\[4\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6854_ _2741_ _2726_ _2746_ _2747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9573_ _0359_ clknet_4_2_0_clk reg_file.reg_storage\[9\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6785_ _1998_ _1113_ _2681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5805_ _1161_ _1720_ _1721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_9_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8524_ _4119_ _4120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5736_ _0682_ _0684_ _1652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8455_ _4080_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5667_ _0706_ _0652_ _0657_ net25 _1583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_115_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7406_ _3220_ _3222_ _3239_ _3240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_5_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4618_ reg_file.reg_storage\[4\]\[3\] reg_file.reg_storage\[5\]\[3\] reg_file.reg_storage\[6\]\[3\]
+ reg_file.reg_storage\[7\]\[3\] _0481_ _0535_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_130_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5598_ _1431_ reg_file.reg_storage\[2\]\[28\] _1486_ _1514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8386_ _4037_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5703__A2 _1586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input67_I pc[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7337_ _3168_ _3176_ _3177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_130_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7268_ net94 _3113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7456__A2 _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6219_ _2116_ _2126_ _2131_ _2026_ _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_9007_ _4429_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8405__A1 reg_file.reg_storage\[14\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7199_ _3049_ _3050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7102__I _1982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__I _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8708__A2 _4241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5758__S _1614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4662__S _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6195__A2 _2105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7144__A1 _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5250__S0 _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8892__A1 _3425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7695__A2 _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6388__I _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5458__A1 _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6655__B1 _2550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8947__A2 _4388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__I _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5630__A1 _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5069__S0 _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6570_ _1132_ _1818_ _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9124__A2 _4496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5521_ _1372_ _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_82_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8240_ _3929_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5241__S0 _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5452_ _0659_ _1368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7686__A2 _3099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8171_ _3884_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6298__I _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5383_ _1178_ _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7122_ net161 _2992_ _2997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_100_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7053_ _2937_ _2576_ _2938_ _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6004_ _1915_ _1918_ _1268_ _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8938__A2 _4381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7955_ net120 _3728_ _3729_ _3742_ _3744_ _3745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_82_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7886_ _2967_ _3534_ _3036_ net47 _3684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6906_ _1057_ _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_128_clk clknet_4_5_0_clk clknet_leaf_128_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_119_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9625_ _0411_ clknet_leaf_83_clk reg_file.reg_storage\[1\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6837_ _2116_ _2730_ _2731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5377__I _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9556_ _0342_ clknet_leaf_118_clk reg_file.reg_storage\[10\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8507_ _4067_ _4109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_135_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9115__A2 _4456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6768_ _2599_ _2621_ _2597_ _2664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9487_ _0273_ clknet_leaf_64_clk reg_file.reg_storage\[8\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7126__A1 net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6699_ _2596_ _2597_ _2598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5719_ _0908_ _1632_ _1634_ _1635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_61_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8438_ _4013_ _4019_ _4066_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8369_ _3919_ _4025_ _4027_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5783__S1 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6652__A3 _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8929__A2 _4381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7767__I net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_119_clk clknet_4_7_0_clk clknet_leaf_119_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9106__A2 _4486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7117__A1 net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6628__B1 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5151__I0 reg_file.reg_storage\[12\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 inst[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_69_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5454__I1 reg_file.reg_storage\[13\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5603__A1 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6581__I _2439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7740_ _3434_ _3548_ _3549_ _3522_ _3550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_87_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4952_ reg_file.reg_storage\[12\]\[23\] reg_file.reg_storage\[13\]\[23\] reg_file.reg_storage\[14\]\[23\]
+ reg_file.reg_storage\[15\]\[23\] _0866_ _0867_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_86_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7671_ _3429_ _3486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4883_ net78 _0798_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _2467_ _2523_ _2047_ _2524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9410_ _0196_ clknet_leaf_4_clk reg_file.reg_storage\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9341_ _0127_ clknet_leaf_115_clk reg_file.reg_storage\[6\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6553_ _2311_ _2312_ _2314_ _2457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_144_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9272_ _0058_ clknet_leaf_81_clk reg_file.reg_storage\[3\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5504_ _0539_ _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6484_ _2387_ _1832_ _2372_ _2389_ _2390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_14_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8223_ _3914_ _3915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5435_ _0736_ _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8608__A1 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8154_ reg_file.reg_storage\[6\]\[3\] _3470_ _3873_ _3875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5366_ _1058_ _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7105_ net6 _2970_ _2972_ _2985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5297_ _1208_ _1210_ _1211_ _1212_ _0784_ _0824_ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_8085_ reg_file.reg_storage\[2\]\[9\] _3831_ _3832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7036_ _2704_ _2921_ _2922_ _2923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__9033__A1 _3989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5842__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6398__A2 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8987_ _3932_ _4411_ _4418_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7938_ _3574_ _3712_ _3029_ _3713_ _3730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_78_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6642__I0 _2290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7869_ _2968_ _3641_ _3642_ net45 _3669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_9608_ _0394_ clknet_leaf_46_clk reg_file.reg_storage\[1\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7898__A2 _3446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9539_ _0325_ clknet_4_4_0_clk reg_file.reg_storage\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6322__A2 _1763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5508__S1 _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7822__A2 _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7889__A2 _3285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6010__A1 _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5747__S1 _1596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5220_ reg_file.reg_storage\[4\]\[13\] reg_file.reg_storage\[5\]\[13\] reg_file.reg_storage\[6\]\[13\]
+ reg_file.reg_storage\[7\]\[13\] _1049_ _1135_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_11_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9153__S _4516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7181__B _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ reg_file.reg_storage\[12\]\[25\] reg_file.reg_storage\[13\]\[25\] reg_file.reg_storage\[14\]\[25\]
+ reg_file.reg_storage\[15\]\[25\] _0855_ _0857_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6576__I _2479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8066__A2 _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5082_ net86 _0889_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9015__A1 reg_file.reg_storage\[1\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8910_ _4195_ _4362_ _4371_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8841_ reg_file.reg_storage\[10\]\[12\] _4209_ _4315_ _4329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8772_ _4260_ _4286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6624__I0 _2264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6017__S _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4824__I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7723_ _3518_ _3534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_59_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5052__A2 _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5984_ _0697_ _0733_ _1794_ _1899_ _1900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_75_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4935_ _0850_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4866_ reg_file.reg_storage\[12\]\[20\] reg_file.reg_storage\[13\]\[20\] reg_file.reg_storage\[14\]\[20\]
+ reg_file.reg_storage\[15\]\[20\] _0780_ _0781_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_75_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6001__A1 _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7654_ reg_file.reg_storage\[5\]\[3\] _3470_ _3458_ _3471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7585_ _3404_ _3405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6605_ _2165_ _2490_ _2507_ _2508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_43_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4797_ _0705_ _0706_ _0708_ _0711_ _0712_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_9324_ _0110_ clknet_leaf_55_clk reg_file.reg_storage\[6\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_rebuffer22_I _1631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6536_ _1666_ _1682_ net206 _2440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9255_ _0041_ clknet_leaf_35_clk reg_file.reg_storage\[3\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6467_ _2076_ _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6687__S _2105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput140 net140 mem_st_dat[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput151 net151 mem_st_dat[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8206_ reg_file.reg_storage\[6\]\[26\] _3903_ _3904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9186_ reg_file.reg_storage\[15\]\[19\] _4536_ _4539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6398_ _1252_ _1772_ _2075_ _2306_ _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_2_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5418_ _1324_ _0913_ _1333_ _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput162 net162 mem_st_dat[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8137_ _3860_ _3861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput195 net195 pc_next[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput173 net173 pc_next[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput184 net184 pc_next[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5349_ _1264_ _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7804__A2 _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8068_ _3821_ _3822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output136_I net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7019_ _2905_ _2906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_98_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7568__A1 _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50_clk clknet_4_10_0_clk clknet_leaf_50_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_80_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4909__I _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__A1 _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7559__A1 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5676__S _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_41_clk clknet_4_8_0_clk clknet_leaf_41_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4720_ reg_file.reg_storage\[4\]\[0\] reg_file.reg_storage\[5\]\[0\] reg_file.reg_storage\[6\]\[0\]
+ reg_file.reg_storage\[7\]\[0\] _0633_ _0635_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_83_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7176__B _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ reg_file.reg_storage\[1\]\[6\] _0569_ _0570_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7731__B2 _3541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7731__A1 net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput31 inst[8] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput20 inst[27] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput64 mem_ld_dat[9] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput42 mem_ld_dat[18] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 mem_ld_dat[28] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4582_ net15 _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7370_ _3204_ _3206_ _3207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput75 pc[19] net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput86 pc[29] net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6321_ _2230_ _2231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_122_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9040_ _3999_ _4445_ _4448_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5345__I0 reg_file.reg_storage\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6252_ _2151_ _2163_ _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_90_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4819__I _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6183_ _2092_ _2095_ _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5203_ _1118_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5134_ reg_file.reg_storage\[2\]\[24\] reg_file.reg_storage\[3\]\[24\] _1049_ _1050_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__9087__I1 _3584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _0887_ _0974_ _0980_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6470__A1 _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_64_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8824_ _4191_ _4312_ _4319_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4554__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8755_ reg_file.reg_storage\[11\]\[10\] _4205_ _4272_ _4277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6773__A2 _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5967_ _1401_ _1881_ _1882_ _1056_ _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_48_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7706_ _0714_ _3518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8686_ _4228_ _4226_ _4229_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_32_clk clknet_4_8_0_clk clknet_leaf_32_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4918_ _0619_ _0631_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_8_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5898_ _1732_ _1814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_7_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7637_ _3454_ _3455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4849_ _0764_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6525__A2 _2429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5385__I _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_73_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7568_ _1236_ _3387_ _3388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_15_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9307_ _0093_ clknet_leaf_85_clk reg_file.reg_storage\[2\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8696__I _3704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6519_ _2332_ _2424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7499_ _3226_ _3321_ _3323_ _3324_ _3325_ net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9238_ _0024_ clknet_leaf_112_clk reg_file.reg_storage\[5\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6289__A1 _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4729__I _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_99_clk clknet_4_15_0_clk clknet_leaf_99_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_9169_ reg_file.reg_storage\[15\]\[12\] _3584_ _4515_ _4529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_110_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6944__I _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8450__A2 _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_82_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5647__S0 _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5016__A2 _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7961__A1 net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7961__B2 _3748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_23_clk clknet_4_1_0_clk clknet_leaf_23_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_108_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7713__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_91_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5575__I0 reg_file.reg_storage\[8\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7724__B net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6452__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _2287_ _2682_ _2762_ _2763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5821_ reg_file.reg_storage\[2\]\[8\] reg_file.reg_storage\[3\]\[8\] _0572_ _1737_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6755__A2 _2651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5752_ _1193_ _1667_ _1668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8540_ _4133_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_14_clk clknet_4_0_0_clk clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_44_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4703_ _0608_ _0613_ _0616_ _0618_ _0605_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_8471_ _3946_ _4075_ _4089_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5683_ _1586_ _1598_ _1599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6507__A2 _2386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4634_ _0555_ net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_7422_ _0914_ _1704_ _1705_ _3255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_5_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5933__I _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5810__S0 _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4565_ _0490_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7353_ _3179_ _3182_ _3191_ net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5191__A1 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6304_ _1958_ _1913_ _2062_ _2215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9023_ reg_file.reg_storage\[1\]\[20\] _4435_ _4439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7284_ net21 _1443_ _3128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_139_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9209__A1 _4006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6235_ _2087_ _2096_ _2147_ _2148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6166_ _1973_ _2080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5117_ reg_file.reg_storage\[1\]\[30\] _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6097_ _2006_ _2011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9140__I _4510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5048_ _0784_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_79_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input12_I inst[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8196__A1 _3682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8807_ _4304_ _4307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5629__S0 _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6999_ _1409_ _2859_ _2861_ _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_48_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8738_ _4267_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_36_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8499__A2 _4074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8669_ _4217_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5557__I0 reg_file.reg_storage\[8\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5182__A1 _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8671__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6674__I _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8974__A3 _3425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6737__A2 _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4748__A1 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5239__B _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6849__I _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ _1920_ _1934_ _1110_ _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_3_clk clknet_4_4_0_clk clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8414__A2 _4051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I inst[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7971_ reg_file.reg_storage\[3\]\[0\] _3758_ _3759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6922_ _2805_ _2806_ _2812_ _2813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9641_ _0427_ clknet_leaf_50_clk reg_file.reg_storage\[4\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6853_ _2742_ _2745_ _2746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_92_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5804_ _1719_ _1720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6533__B _2437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6784_ _2165_ _2678_ _2679_ _2680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_9572_ _0358_ clknet_leaf_119_clk reg_file.reg_storage\[9\]\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5400__A2 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8523_ _4015_ _4118_ _4119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5735_ _1579_ _1602_ _1621_ _1650_ _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5666_ _1581_ _1582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8454_ reg_file.reg_storage\[13\]\[2\] _3926_ _4079_ _4080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7405_ _3213_ _3229_ _3239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4617_ reg_file.reg_storage\[12\]\[3\] reg_file.reg_storage\[13\]\[3\] reg_file.reg_storage\[14\]\[3\]
+ reg_file.reg_storage\[15\]\[3\] _0481_ _0539_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_142_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5597_ _1464_ reg_file.reg_storage\[3\]\[28\] _1513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8385_ reg_file.reg_storage\[14\]\[8\] _3943_ _4035_ _4037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5703__A3 _1618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4911__A1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7336_ _3173_ _3175_ _3176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7267_ net93 net94 _3098_ _3112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__9071__S _4466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6218_ _2046_ _2130_ _2131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9006_ reg_file.reg_storage\[1\]\[13\] _3597_ _4414_ _4429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7198_ _0608_ _3048_ _3049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8405__A2 _4038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6149_ _2062_ _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6719__A2 _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4742__I _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7144__A2 _3010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__A1 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_53_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5250__S1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6655__B2 _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_68_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5069__S1 _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4652__I _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7907__B2 _1881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7383__A2 _3205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_126_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5520_ reg_file.reg_storage\[8\]\[27\] reg_file.reg_storage\[9\]\[27\] reg_file.reg_storage\[10\]\[27\]
+ reg_file.reg_storage\[11\]\[27\] _1419_ _1423_ _1436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_80_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8332__A1 reg_file.reg_storage\[7\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5451_ reg_file.reg_storage\[1\]\[26\] _1366_ _1364_ _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8995__S _4421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5241__S1 _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8170_ reg_file.reg_storage\[6\]\[10\] _3557_ _3879_ _3884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6894__A1 _2777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5382_ _1242_ _1267_ _1297_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7121_ _1690_ _2995_ _2996_ net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_1_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7052_ _2937_ _2304_ _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6003_ _1916_ _1917_ _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6528__B _2076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7071__A1 _2217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7954_ _3715_ _3370_ _3743_ _3744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6905_ _1379_ _1881_ _1882_ _2797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_49_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7885_ _3660_ _3682_ _3683_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4562__I _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9624_ _0410_ clknet_leaf_82_clk reg_file.reg_storage\[1\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6836_ _2637_ _2729_ _2040_ _2730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7374__A2 _3202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ _2623_ _2598_ _2630_ _2652_ _2663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_9555_ _0341_ clknet_leaf_76_clk reg_file.reg_storage\[10\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8506_ _3993_ _4069_ _4108_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5480__S1 _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5718_ _0680_ _1583_ _1633_ _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__8323__A1 reg_file.reg_storage\[7\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9486_ _0272_ clknet_leaf_66_clk reg_file.reg_storage\[8\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6698_ _2593_ _2595_ _2597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_72_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8437_ reg_file.reg_storage\[14\]\[31\] _4017_ _4066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5649_ _1386_ _1564_ _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8368_ reg_file.reg_storage\[14\]\[1\] _4026_ _4027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output166_I net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7319_ _3159_ _3151_ _3160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8299_ _3970_ _3959_ _3972_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5342__B _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5860__A2 _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__S _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7984__S _3769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__B _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8865__A2 _4338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5128__A1 _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6628__A1 _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5151__I1 reg_file.reg_storage\[13\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4734__S0 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4647__I _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 inst[15] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_69_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4951_ _0856_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4882_ _0748_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7670_ _3484_ _3485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6621_ _1149_ _1164_ _2523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5367__A1 _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9340_ _0126_ clknet_leaf_103_clk reg_file.reg_storage\[6\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6552_ _2240_ _2236_ _2241_ _2279_ _2456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_125_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5503_ _1418_ _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5119__A1 _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8856__A2 _4331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9271_ _0057_ clknet_leaf_81_clk reg_file.reg_storage\[3\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6483_ _2387_ _1832_ _2373_ _2388_ _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_42_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5427__B _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8222_ _3913_ _3914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6102__I _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5914__I0 _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5434_ _1338_ _1347_ _0733_ _1349_ _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8153_ _3874_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7104_ _2984_ _2983_ _2980_ net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8608__A2 _4171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5365_ _1280_ _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5296_ reg_file.reg_storage\[8\]\[9\] reg_file.reg_storage\[9\]\[9\] reg_file.reg_storage\[10\]\[9\]
+ reg_file.reg_storage\[11\]\[9\] _0778_ _0803_ _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8084_ _3816_ _3831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5162__B _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7035_ _2135_ _2710_ _2922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9033__A2 _4406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5842__A2 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8986_ reg_file.reg_storage\[1\]\[4\] _4412_ _4418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7937_ _3547_ _3729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_77_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7868_ _3660_ _3667_ _3668_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6819_ _2697_ _1542_ _2373_ _2713_ _2714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_9607_ _0393_ clknet_leaf_22_clk reg_file.reg_storage\[1\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7347__A2 _3183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7799_ _3024_ _3602_ _3604_ _3537_ _3605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_108_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9538_ _0324_ clknet_leaf_121_clk reg_file.reg_storage\[10\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8847__A2 _4331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9469_ _0255_ clknet_leaf_88_clk reg_file.reg_storage\[12\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6858__A1 _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__B _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9024__A2 _4437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6682__I _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7035__A1 _2135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5597__A1 _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7338__A2 net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6546__C2 _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4578__S _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_102_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5150_ reg_file.reg_storage\[1\]\[25\] _1065_ _1063_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5081_ _0996_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_47_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9015__A2 _4424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7688__I _3501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8840_ _4328_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_48_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8771_ _4220_ _4281_ _4285_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5132__S0 _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6624__I1 _2525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5983_ _1896_ _1897_ _1898_ _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_7722_ net64 net41 _3412_ _3533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4934_ _0695_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4865_ _0760_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4840__I _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5936__I _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7653_ _3469_ _3470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7584_ _2970_ _1981_ _3404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_74_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6604_ _2259_ _2493_ _2499_ _2506_ _2507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4796_ net6 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_7_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6535_ _2153_ _2439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9323_ _0109_ clknet_leaf_9_clk reg_file.reg_storage\[6\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9254_ _0040_ clknet_leaf_42_clk reg_file.reg_storage\[3\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8205_ _3860_ _3903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6466_ _2080_ _2373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput130 net130 mem_ld_mask[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput141 net141 mem_st_dat[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput152 net152 mem_st_dat[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_120_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5671__I _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9185_ _4516_ _4538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6397_ _2303_ _2169_ _2305_ _2306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5417_ _1014_ _1332_ _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input42_I mem_ld_dat[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput163 net163 mem_st_dat[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_8136_ _3388_ _3809_ _3860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput174 net174 pc_next[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput185 net185 pc_next[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_11_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5348_ _1254_ _1263_ _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_100_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8067_ _3815_ _3821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7265__B2 _3110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput196 net196 pc_next[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7018_ _1010_ _2905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5279_ net66 _0888_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7017__A1 _2725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5371__S0 _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output129_I net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5123__S0 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5579__A1 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8969_ _4404_ _4405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_104_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8517__A1 reg_file.reg_storage\[13\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8222__I _3913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5782__S _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5581__I net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7559__A2 _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6231__A2 _1902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8508__A1 reg_file.reg_storage\[13\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5756__I _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5990__A1 _1795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4650_ net14 _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput10 inst[18] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput21 inst[28] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput43 mem_ld_dat[19] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput54 mem_ld_dat[29] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4581_ reg_file.reg_storage\[8\]\[0\] reg_file.reg_storage\[9\]\[0\] reg_file.reg_storage\[10\]\[0\]
+ reg_file.reg_storage\[11\]\[0\] _0497_ _0500_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput32 inst[9] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6320_ _2229_ _0669_ _1354_ _1759_ _2230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_141_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput76 pc[1] net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput65 pc[0] net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput87 pc[2] net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4928__S0 _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6251_ _2161_ _2162_ _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7495__A1 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6182_ _2093_ _2094_ _2095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5202_ _1114_ _1108_ _1117_ _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5133_ _0778_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5064_ _0979_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6470__A2 _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8823_ reg_file.reg_storage\[10\]\[4\] _4313_ _4319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_88_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8754_ _4202_ _4262_ _4276_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5966_ _1351_ _1457_ _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7705_ _3022_ _3517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8685_ reg_file.reg_storage\[8\]\[20\] _4223_ _4229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4917_ _0797_ _0832_ _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5897_ _1756_ _1812_ _1813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_23_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4848_ _0763_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_63_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7636_ _2085_ _3446_ _3450_ _3452_ _3453_ _3454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__4570__I _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9306_ _0092_ clknet_leaf_85_clk reg_file.reg_storage\[2\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5733__A1 _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7567_ net2 _3387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_62_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4779_ _0694_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6518_ _2246_ _2145_ _2423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7498_ _3272_ net114 _3325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6289__A2 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9237_ _0023_ clknet_leaf_119_clk reg_file.reg_storage\[5\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6449_ _2343_ _2319_ _2321_ _2356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9168_ _4528_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8119_ _3705_ _3812_ _3850_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7238__B2 _3085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9099_ _3966_ _4481_ _4485_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_110_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5777__S _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5647__S1 _1537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8887__I _4354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5575__I1 reg_file.reg_storage\[9\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7477__A1 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5583__S0 _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5820_ reg_file.reg_storage\[8\]\[8\] reg_file.reg_storage\[9\]\[8\] reg_file.reg_storage\[10\]\[8\]
+ reg_file.reg_storage\[11\]\[8\] _1605_ _1361_ _1736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_88_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4591__S _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5963__A1 _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5751_ _1666_ _1667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8470_ reg_file.reg_storage\[13\]\[9\] _4088_ _4089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _0617_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5682_ _1597_ _0490_ _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7421_ _0952_ _3253_ _3254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_127_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4633_ _0543_ _0549_ _0554_ _0487_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_130_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5810__S1 _1672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7352_ _3157_ net101 _3158_ _3190_ _3191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4564_ _0489_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_69_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6303_ _2016_ _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7283_ _3124_ _3126_ _3127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_110_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9022_ _3973_ _4437_ _4438_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6234_ _2133_ _2141_ _2146_ _2147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5574__S0 _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6140__A1 _2046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8968__A1 _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6165_ _2004_ _2079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5116_ reg_file.reg_storage\[4\]\[30\] reg_file.reg_storage\[5\]\[30\] reg_file.reg_storage\[6\]\[30\]
+ reg_file.reg_storage\[7\]\[30\] _0811_ _0761_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6096_ _2003_ _2010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5047_ reg_file.reg_storage\[8\]\[19\] reg_file.reg_storage\[9\]\[19\] reg_file.reg_storage\[10\]\[19\]
+ reg_file.reg_storage\[11\]\[19\] _0921_ _0961_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4565__I _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8196__A2 _3895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8806_ _4305_ _4306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6998_ _2860_ _2838_ _2886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5629__S1 _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5949_ _1635_ _1636_ _1580_ _1601_ _1865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_48_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8737_ reg_file.reg_storage\[11\]\[2\] _4185_ _4266_ _4267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_36_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8668_ reg_file.reg_storage\[8\]\[15\] _4216_ _4186_ _4217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8599_ _4004_ _4164_ _4166_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5557__I1 reg_file.reg_storage\[9\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7619_ _3437_ _3438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5182__A2 _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8120__A2 _3813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5890__B1 _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7631__A1 _3447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5945__A1 _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9136__A1 reg_file.reg_storage\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8410__I _4029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_144_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8111__A2 _3844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5556__S0 _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5308__S0 _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7622__A1 _3436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7970_ _3755_ _3758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6921_ _2810_ _2811_ _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9640_ _0426_ clknet_leaf_58_clk reg_file.reg_storage\[4\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_85_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6852_ _1844_ _2744_ _2745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_76_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5803_ _0671_ _1710_ _1718_ _1719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5210__S _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9571_ _0357_ clknet_leaf_134_clk reg_file.reg_storage\[9\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9127__A1 _4006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _2668_ _2677_ _2679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_71_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8522_ _3395_ _4117_ _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_33_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5734_ _1635_ _1636_ _1649_ _1650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_45_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8453_ _4078_ _4079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5665_ _0728_ _0681_ _0683_ _1581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_8384_ _4036_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7404_ net74 _1603_ _3238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4616_ _0498_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__S0 _1607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5596_ reg_file.reg_storage\[4\]\[28\] reg_file.reg_storage\[5\]\[28\] reg_file.reg_storage\[6\]\[28\]
+ reg_file.reg_storage\[7\]\[28\] _1418_ _1447_ _1512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7335_ _3124_ _3126_ _3129_ _3174_ _3175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__8102__A2 _3831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7266_ _3077_ _3099_ _3111_ net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9005_ _4428_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6217_ _2128_ _2129_ _2022_ _2130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7197_ _3047_ _3048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6148_ _1241_ _2062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6079_ _0696_ _1905_ _1993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output111_I net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8169__A2 _3869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6352__A1 _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5538__S0 _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7852__A1 _3255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4666__A1 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4933__I _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9109__A1 _3980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8580__A2 _4152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5450_ reg_file.reg_storage\[2\]\[26\] reg_file.reg_storage\[3\]\[26\] _1359_ _1366_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6796__S _2183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5381_ _1269_ _1283_ _1296_ _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7120_ net160 _2992_ _2996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_100_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7051_ _2926_ _1874_ _2937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7843__A1 _3228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6002_ _0849_ _0796_ _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8399__A2 _4038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5004__I _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5701__S0 _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7953_ _1481_ _3505_ _3743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6904_ _2061_ _2681_ _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4843__I _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5082__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7884_ reg_file.reg_storage\[5\]\[21\] _3658_ _3683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9623_ _0409_ clknet_leaf_81_clk reg_file.reg_storage\[1\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6835_ _2690_ _2728_ _2007_ _2729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8571__A2 _4147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9554_ _0340_ clknet_leaf_67_clk reg_file.reg_storage\[10\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6766_ _2643_ _2648_ _2662_ net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_46_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8505_ reg_file.reg_storage\[13\]\[25\] _4070_ _4108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5717_ net9 _0701_ _0682_ _0684_ _1633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_127_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6697_ _2593_ _2595_ _2596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5674__I _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9485_ _0271_ clknet_leaf_11_clk reg_file.reg_storage\[8\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9146__I _4515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8436_ _4010_ _4061_ _4065_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5648_ _1445_ _1563_ _1564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input72_I pc[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5768__S0 _1606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4896__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8367_ _4022_ _4026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5579_ _1114_ _1481_ _1494_ _1495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_14_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8298_ reg_file.reg_storage\[7\]\[18\] _3971_ _3972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7318_ _3145_ _1671_ _3159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4991__S1 _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7249_ _3059_ net124 _3061_ _3095_ _3096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_output159_I net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7062__A2 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5073__A1 _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4753__I _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_16_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6573__A1 _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5128__A2 _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6325__A1 _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8895__I _4361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7825__A1 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5025__S _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5687__I0 _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7840__A4 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5151__I2 reg_file.reg_storage\[14\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4734__S1 _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput8 inst[16] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_69_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4950_ _0854_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_129_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4881_ _0791_ _0796_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9167__S _4522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6620_ _2254_ _2407_ _2520_ _2521_ _2522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_52_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8071__S _3822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6551_ _2236_ _2279_ _2455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5502_ _1390_ _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_82_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9270_ _0056_ clknet_leaf_116_clk reg_file.reg_storage\[3\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6482_ _2387_ _1832_ _2077_ _2388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6316__A1 _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8221_ _3388_ _3754_ _3913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6867__A2 _2269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5914__I1 _1829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5433_ _0697_ _1348_ _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8152_ reg_file.reg_storage\[6\]\[2\] _3456_ _3873_ _3874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5364_ _1279_ _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7103_ _2984_ _2974_ _2980_ net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7816__A1 _3547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8083_ _3830_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5295_ reg_file.reg_storage\[12\]\[9\] reg_file.reg_storage\[13\]\[9\] reg_file.reg_storage\[14\]\[9\]
+ reg_file.reg_storage\[15\]\[9\] _0778_ _0803_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7034_ _2245_ _2819_ _2920_ _2424_ _2921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_97_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5055__A1 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8985_ _4417_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7936_ _3417_ _3728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_78_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_52_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7867_ reg_file.reg_storage\[5\]\[19\] _3658_ _3668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9606_ _0392_ clknet_leaf_43_clk reg_file.reg_storage\[1\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6818_ _2697_ _1542_ _2374_ _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8544__A2 _4128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7798_ _3410_ _3603_ _3604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_102_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6749_ _2645_ _2578_ _2646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9537_ _0323_ clknet_leaf_127_clk reg_file.reg_storage\[10\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9468_ _0254_ clknet_leaf_90_clk reg_file.reg_storage\[12\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_67_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6307__A1 _2052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_110_clk_I clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8419_ reg_file.reg_storage\[14\]\[23\] _4024_ _4056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_21_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9399_ _0185_ clknet_leaf_88_clk reg_file.reg_storage\[14\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_131_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7807__A1 _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7995__S _3775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8783__A2 _4288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8535__A2 _4129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4580__I0 reg_file.reg_storage\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5080_ _0995_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7274__A2 _3116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8770_ reg_file.reg_storage\[11\]\[17\] _4275_ _4285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8774__A2 _4281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5132__S1 _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5982_ _1895_ _1871_ _1894_ _1898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7721_ _3532_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4933_ _0848_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_75_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4864_ _0779_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6537__A1 _2439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7652_ _3468_ _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6603_ _2193_ _2505_ _2506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7583_ _3402_ _3403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4795_ net5 _0709_ _0710_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6534_ _2438_ net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_9322_ _0108_ clknet_leaf_7_clk reg_file.reg_storage\[6\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4643__S0 _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9253_ _0039_ clknet_leaf_38_clk reg_file.reg_storage\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6465_ _2173_ _2372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8204_ _3710_ _3862_ _3902_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5416_ _1325_ _1329_ _1330_ _1331_ _0648_ _0823_ _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
Xoutput142 net142 mem_st_dat[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput120 net120 mem_addr[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput131 net131 mem_ld_mask[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_140_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9184_ _3969_ _4531_ _4537_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6396_ _2303_ _2304_ _2305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput164 net164 mem_st_dat[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput153 net153 mem_st_dat[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_101_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8135_ _3751_ _3813_ _3859_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4568__I _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5347_ _0890_ _1262_ _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput175 net175 pc_next[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput186 net186 pc_next[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8066_ _3443_ _3818_ _3820_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5278_ _1193_ _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7265__A2 net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput197 net197 pc_next[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input35_I mem_ld_dat[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7017_ _2725_ _2891_ _2899_ _2904_ net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__5276__A1 _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8214__A1 _3740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5371__S1 _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8765__A2 _4281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5123__S1 _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8968_ _3397_ _3753_ _4404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__A2 _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7919_ _3631_ _3713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_104_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8899_ _4359_ _4365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_26_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6528__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9190__A2 _4536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire203 _2088_ net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_133_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6700__A1 _2573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5019__A1 _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4873__S0 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4941__I _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9181__A2 _4531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4580_ reg_file.reg_storage\[12\]\[0\] reg_file.reg_storage\[13\]\[0\] reg_file.reg_storage\[14\]\[0\]
+ reg_file.reg_storage\[15\]\[0\] _0497_ _0500_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_83_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 inst[19] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 inst[29] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_25_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput33 mem_ld_dat[0] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput44 mem_ld_dat[1] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput55 mem_ld_dat[2] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput66 pc[10] net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput77 pc[20] net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput88 pc[30] net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4928__S1 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6250_ _1292_ _2156_ _2159_ _2162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_110_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5050__S0 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6181_ _1992_ _1993_ _1994_ _2094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5201_ net159 _1116_ _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5132_ reg_file.reg_storage\[4\]\[24\] reg_file.reg_storage\[5\]\[24\] reg_file.reg_storage\[6\]\[24\]
+ reg_file.reg_storage\[7\]\[24\] _0767_ _1047_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_58_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5258__A1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5063_ _0533_ _0977_ _0978_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8822_ _4318_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4851__I _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8753_ reg_file.reg_storage\[11\]\[9\] _4275_ _4276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5965_ _0740_ _1381_ _1480_ _1881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_4
XANTENNA__5430__A1 _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7704_ net63 net40 _3027_ _3516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8684_ _3674_ _4228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4916_ _0829_ _0831_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5896_ _1802_ _1775_ _1808_ _1773_ _1811_ _1812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_75_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4847_ _0623_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7635_ _3066_ _3401_ _1238_ _3402_ _3453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_105_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9305_ _0091_ clknet_leaf_85_clk reg_file.reg_storage\[2\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7566_ _3045_ _3381_ _3382_ _3386_ net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4778_ _0680_ _0689_ _0693_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_132_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6517_ _2113_ _2328_ _2420_ _2421_ _2422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7497_ _3041_ _3324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_31_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9236_ _0022_ clknet_leaf_26_clk reg_file.reg_storage\[5\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6448_ _1215_ _1753_ _2354_ _2355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_9167_ reg_file.reg_storage\[15\]\[11\] _3567_ _4522_ _4528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6379_ _2016_ _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8118_ reg_file.reg_storage\[2\]\[24\] _3813_ _3850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7238__A2 net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output141_I net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9098_ reg_file.reg_storage\[4\]\[17\] _4475_ _4485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8986__A2 _4412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8049_ reg_file.reg_storage\[3\]\[31\] _3756_ _3806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5344__S1 _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4761__I _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9163__A2 _4525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8910__A2 _4362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5280__S0 _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9064__I _4465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_100_clk clknet_4_15_0_clk clknet_leaf_100_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_0_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5583__S1 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6637__B _2537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6988__A1 _2113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5660__A1 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5099__S0 _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7401__A2 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4846__S0 _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5750_ _0735_ _1656_ _1665_ _1666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__4671__I net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5681_ _1589_ _1592_ _1593_ _1594_ _1595_ _1596_ _1597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_56_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4701_ _0609_ _0587_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7420_ _1637_ _3253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4632_ _0551_ _0553_ _0543_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5271__S0 _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5715__A2 _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6912__A1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7351_ _3187_ _3189_ _3190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_25_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4563_ _0488_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_111_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6302_ _2211_ _2212_ _2045_ _2213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7282_ _3105_ _3104_ _3108_ _3125_ _3126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_4_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9021_ reg_file.reg_storage\[1\]\[19\] _4435_ _4438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6233_ _2069_ _2145_ _2146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5574__S1 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9534__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6164_ _1947_ _2064_ _2077_ _2078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8968__A2 _3753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6095_ _1012_ _1101_ _2008_ _2009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5115_ net88 _0889_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5046_ reg_file.reg_storage\[12\]\[19\] reg_file.reg_storage\[13\]\[19\] reg_file.reg_storage\[14\]\[19\]
+ reg_file.reg_storage\[15\]\[19\] _0896_ _0961_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5651__A1 _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8805_ _4304_ _4305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6997_ _2883_ _2884_ _2885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_48_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8053__I _3808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5948_ _1862_ _1863_ _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8736_ _4265_ _4266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_36_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7156__B2 _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7156__A1 _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9085__S _4472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8667_ _3622_ _4216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5879_ net76 _0747_ _0752_ _1332_ _1795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_8598_ reg_file.reg_storage\[12\]\[28\] _4162_ _4166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5557__I2 reg_file.reg_storage\[10\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7618_ _0594_ _3034_ _3437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_output189_I net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7549_ _3248_ net120 _3371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9219_ _0005_ clknet_leaf_0_clk reg_file.reg_storage\[5\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5890__B2 _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9059__I _4461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A2 _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7147__A1 _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7751__B net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5556__S1 _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5308__S1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6920_ _1878_ _2809_ _2811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_85_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6851_ _2743_ _2721_ _2744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5802_ _1670_ _1717_ _1718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9570_ _0356_ clknet_leaf_120_clk reg_file.reg_storage\[9\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9127__A2 _4498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6782_ _2668_ _2677_ _2678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8521_ net31 _3390_ _4117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7138__A1 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5733_ _0968_ net238 _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_143_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8886__A1 _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5664_ _0933_ _1580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8452_ _4072_ _4078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7689__A2 _3444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8383_ reg_file.reg_storage\[14\]\[7\] _3940_ _4035_ _4036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7403_ _0936_ _3233_ _3237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_26_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4615_ reg_file.reg_storage\[1\]\[3\] _0537_ _0535_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5595_ _1413_ _1510_ _1511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5795__S1 _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8638__A1 reg_file.reg_storage\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7334_ _3137_ _3169_ _3174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6121__I _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8249__S _3928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7265_ _3100_ net125 _3101_ _3110_ _3111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9004_ reg_file.reg_storage\[1\]\[12\] _3584_ _4421_ _4428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6216_ _1957_ _1964_ _2028_ _2129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7196_ _0613_ _3047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6147_ _2060_ _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4576__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5872__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6821__B1 _2712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8810__A1 _3865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5624__A1 _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6078_ _1334_ _1985_ _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5029_ reg_file.reg_storage\[8\]\[18\] reg_file.reg_storage\[9\]\[18\] reg_file.reg_storage\[10\]\[18\]
+ reg_file.reg_storage\[11\]\[18\] _0810_ _0942_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__7377__A1 _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output104_I net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5200__I _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8719_ _3750_ _4252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5538__S1 _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__I _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5870__I _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_79_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9054__A1 reg_file.reg_storage\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4666__A2 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7604__A2 _3421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_88_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9109__A2 _4488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5226__S0 _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_97_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5380_ _1294_ _1295_ _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8096__A2 _3831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8069__S _3822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7050_ _2930_ _2934_ _2935_ _2936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9045__A1 _4006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6001_ _1847_ _1148_ _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5854__A1 _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7952_ _3712_ _3603_ _3700_ _3742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_89_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7500__I net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5701__S1 _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6903_ _2284_ _2341_ _2794_ _2610_ _2795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5082__A2 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9622_ _0408_ clknet_leaf_81_clk reg_file.reg_storage\[1\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7883_ _3681_ _3682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_18_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8020__A2 _3789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6834_ _1852_ _2106_ _0832_ _2728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_9_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6031__A1 _1795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9553_ _0339_ clknet_leaf_67_clk reg_file.reg_storage\[10\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ _2404_ _2654_ _2661_ _2641_ _2662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_58_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9484_ _0270_ clknet_leaf_65_clk reg_file.reg_storage\[8\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8504_ _3990_ _4069_ _4107_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8331__I _3913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5716_ _0734_ _1631_ _1632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_73_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6052__S _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8435_ reg_file.reg_storage\[14\]\[30\] _4017_ _4065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5176__B _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6696_ _1863_ _2594_ _2595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5647_ _1558_ _1560_ _1561_ _1562_ _1534_ _1537_ _1563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5768__S1 _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8366_ _4024_ _4025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5578_ _1386_ _1493_ _1494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input65_I pc[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5690__I _1605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8297_ _3921_ _3971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__9162__I _4510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7317_ _3052_ _3158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7248_ _3087_ _3090_ _3094_ _3095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__9036__A1 _3992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5845__A1 _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7179_ _1982_ _3032_ _3033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9252__CLK clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8011__A2 _3778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8241__I _3468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5208__S0 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6325__A2 _2234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8078__A2 _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5687__I1 _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5836__A1 _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5105__I _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4944__I _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput9 inst[17] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_69_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_71_clk clknet_4_9_0_clk clknet_leaf_71_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6013__A1 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4880_ _0795_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5775__I _1690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8151__I _3872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6564__A2 _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6550_ _1991_ _2452_ _2453_ _2090_ _2454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_28_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5501_ _1385_ _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_131_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6481_ _1959_ _2387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_8220_ _3911_ _3912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_124_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5432_ _0731_ _1345_ _1348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8151_ _3872_ _3873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_11_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5363_ _1270_ _0620_ _0834_ _1278_ _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_7102_ _1982_ _2984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_140_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5390__I3 reg_file.reg_storage\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7667__I2 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8082_ reg_file.reg_storage\[2\]\[8\] _3531_ _3828_ _3830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5294_ reg_file.reg_storage\[1\]\[9\] _1209_ _0803_ _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7816__A2 _3618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7033_ _2362_ _2917_ _2919_ _2920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8326__I _3992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8984_ reg_file.reg_storage\[1\]\[3\] _3469_ _4415_ _4417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7230__I net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7935_ _3722_ _3726_ _3727_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62_clk clknet_4_11_0_clk clknet_leaf_62_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7866_ _3666_ _3667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9605_ _0391_ clknet_leaf_38_clk reg_file.reg_storage\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6817_ _2704_ _2140_ _2224_ _2705_ _2711_ _2712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7797_ _3518_ _3032_ net56 _3603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_102_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9157__I _4510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8061__I _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9536_ _0322_ clknet_leaf_128_clk reg_file.reg_storage\[10\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6748_ _2644_ net239 _2645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9467_ _0253_ clknet_leaf_97_clk reg_file.reg_storage\[12\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6679_ _2575_ _2578_ _2579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9398_ _0184_ clknet_leaf_87_clk reg_file.reg_storage\[14\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8418_ _3984_ _4051_ _4055_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_21_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8349_ reg_file.reg_storage\[7\]\[30\] _3914_ _4011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7807__A2 _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9009__A1 reg_file.reg_storage\[1\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6491__A1 _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8236__I _3454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5677__S0 _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5796__S _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_53_clk clknet_4_10_0_clk clknet_leaf_53_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8172__S _3879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_40_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8299__A2 _3959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5601__S0 _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4939__I _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4580__I1 reg_file.reg_storage\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8471__A2 _4075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8146__I _3868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_139_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6785__A2 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5981_ _1782_ _0718_ _1789_ _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
Xclkbuf_leaf_44_clk clknet_4_8_0_clk clknet_leaf_44_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7720_ reg_file.reg_storage\[5\]\[8\] _3531_ _3492_ _3532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8082__S _3828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4932_ _0835_ _0846_ _0847_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7651_ _2148_ _3460_ _3463_ _3467_ _3468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_129_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4863_ _0778_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6602_ _2017_ _2224_ _2504_ _2505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4794_ _0699_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7582_ _3392_ _3402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_144_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9321_ _0107_ clknet_leaf_50_clk reg_file.reg_storage\[6\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6533_ _2087_ _2419_ _2437_ _2438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_55_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4643__S1 _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9252_ _0038_ clknet_4_7_0_clk reg_file.reg_storage\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6464_ _1217_ _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xoutput110 net110 mem_addr[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_141_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4849__I _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8203_ reg_file.reg_storage\[6\]\[25\] _3863_ _3902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5415_ reg_file.reg_storage\[8\]\[1\] reg_file.reg_storage\[9\]\[1\] reg_file.reg_storage\[10\]\[1\]
+ reg_file.reg_storage\[11\]\[1\] _0770_ _1271_ _1331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput132 net132 mem_ld_mask[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput143 net143 mem_st_dat[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput121 net211 mem_addr[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_113_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9183_ reg_file.reg_storage\[15\]\[18\] _4536_ _4537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6395_ _2170_ _2304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput165 net165 mem_st_dat[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput154 net154 mem_st_dat[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8134_ reg_file.reg_storage\[2\]\[31\] _3811_ _3859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5346_ _1255_ _1259_ _1260_ _1261_ _0785_ _0825_ _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput176 net176 pc_next[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8257__S _3941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8462__A2 _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8065_ reg_file.reg_storage\[2\]\[1\] _3819_ _3820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5277_ _1192_ _1193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput198 net198 pc_next[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput187 net187 pc_next[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7016_ _2903_ _2904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_34_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input28_I inst[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6225__A1 _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8967_ _4252_ _4357_ _4403_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5659__S0 _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7918_ _2977_ _3712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_104_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_35_clk clknet_4_2_0_clk clknet_leaf_35_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_26_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8898_ _4177_ _4362_ _4364_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7849_ _3010_ _3449_ _3651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_133_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9519_ _0305_ clknet_leaf_64_clk reg_file.reg_storage\[11\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6700__A2 _2566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_52_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7661__B1 _3474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4873__S1 _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_26_clk clknet_4_3_0_clk clknet_leaf_26_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7716__A1 _3526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput12 inst[1] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput34 mem_ld_dat[10] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput45 mem_ld_dat[20] net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput23 inst[2] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput56 mem_ld_dat[30] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8141__A1 _3421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput67 pc[11] net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput78 pc[21] net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput89 pc[31] net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8692__A2 _4226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5050__S1 _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5200_ _1115_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6180_ _1309_ _1989_ _2093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_51_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5131_ _0983_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_58_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5258__A2 _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _0680_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_66_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8821_ reg_file.reg_storage\[10\]\[3\] _4189_ _4316_ _4318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7955__A1 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8752_ _4260_ _4275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6758__A2 _2429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7703_ _3514_ _3515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_17_clk clknet_4_0_0_clk clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5964_ _1878_ _1879_ _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8683_ _4225_ _4226_ _4227_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_23_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5895_ _1810_ _1772_ _1811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4915_ _0830_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5981__A3 _1789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7634_ _3024_ _3451_ _3414_ _3452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_118_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4846_ reg_file.reg_storage\[4\]\[20\] reg_file.reg_storage\[5\]\[20\] reg_file.reg_storage\[6\]\[20\]
+ reg_file.reg_storage\[7\]\[20\] _0758_ _0761_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_8_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7565_ _3209_ net121 _3385_ _3386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9304_ _0090_ clknet_leaf_82_clk reg_file.reg_storage\[2\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6516_ _1999_ _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4777_ _0690_ _0511_ _0691_ _0692_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_132_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer20_I _1506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7496_ _3317_ _3322_ _3323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__8683__A2 _4226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9235_ _0021_ clknet_leaf_78_clk reg_file.reg_storage\[5\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6447_ _2318_ _2353_ _2354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9166_ _4527_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6378_ _2116_ _2285_ _2286_ _2287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_clkbuf_leaf_19_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5329_ reg_file.reg_storage\[1\]\[7\] _1244_ _0642_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8117_ _3696_ _3819_ _3849_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9097_ _3963_ _4481_ _4484_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8048_ _3746_ _3801_ _3805_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_110_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output134_I net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__I _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7946__A1 _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7574__B net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5575__I3 reg_file.reg_storage\[11\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5280__S1 _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4932__A1 _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8674__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7882__B1 _3678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9080__I _4460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6988__A2 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5099__S1 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4846__S1 _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5680_ _1235_ _1596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_84_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4700_ _0615_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7165__A2 _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5176__A1 _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8362__A1 _3760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ _0528_ _0552_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6912__A2 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5271__S1 _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7350_ _3168_ _3176_ _3188_ _3189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4562_ _0487_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8665__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6301_ _2004_ _1926_ _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_40_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7281_ _3113_ _3116_ _3102_ _3097_ _3125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5023__S1 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9020_ _4415_ _4437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_6_clk clknet_4_6_0_clk clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6232_ _2035_ _2143_ _2144_ _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_110_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8417__A2 _4024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6163_ _2076_ _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6094_ _2007_ _2008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5114_ _0909_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5045_ _0836_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_108_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8334__I _3725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__I _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8804_ _3809_ _4171_ _4304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6996_ _2879_ _2882_ _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5947_ _1632_ _1634_ _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_8735_ _4259_ _4265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_36_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8666_ _4213_ _4214_ _4215_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7617_ net129 _3435_ _3436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8353__A1 reg_file.reg_storage\[7\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5167__A1 _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input95_I pc[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5878_ _1343_ _1350_ _1793_ _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8597_ _4000_ _4164_ _4165_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_117_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5557__I3 reg_file.reg_storage\[11\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__I _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4829_ _0744_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_133_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7548_ _3368_ _3369_ _3370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7479_ net81 _1444_ _3307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_102_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6667__A1 _1580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9218_ _0004_ clknet_leaf_18_clk reg_file.reg_storage\[5\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8408__A2 _4049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5134__S _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9149_ reg_file.reg_storage\[15\]\[3\] _3469_ _4516_ _4518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_126_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9081__A2 _4475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7092__A1 _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8244__I _3477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7395__A2 _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_135_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5158__A1 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9075__I _4460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6850_ _1577_ _2439_ _2743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5801_ _1604_ _1716_ _1717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6781_ _1849_ _2676_ _2677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_69_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8520_ _4013_ _4070_ _4116_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5732_ _1647_ _1648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_57_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8886__A2 _4171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5663_ _1543_ _1556_ _1567_ _1578_ _1579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_44_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8451_ _3919_ _4075_ _4077_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_143_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8382_ _4023_ _4035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7402_ _3226_ _3232_ _3235_ _3179_ _3236_ net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_TAPCELL_ROW_13_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4614_ reg_file.reg_storage\[2\]\[3\] reg_file.reg_storage\[3\]\[3\] _0496_ _0537_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5594_ net21 _1402_ _1510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7333_ _3154_ _3161_ _3170_ _3172_ _3173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_13_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9003_ _4427_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6558__B _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7264_ _3104_ _3109_ _3110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4857__I _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6215_ _2104_ _1908_ _1909_ _2127_ _2128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7195_ _0606_ _3042_ _3043_ _3046_ net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7233__I _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5321__A1 _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6146_ _2059_ _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5624__A2 _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6077_ _1986_ _1987_ _1990_ _1991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5180__S0 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5688__I _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ reg_file.reg_storage\[12\]\[18\] reg_file.reg_storage\[13\]\[18\] reg_file.reg_storage\[14\]\[18\]
+ reg_file.reg_storage\[15\]\[18\] _0810_ _0942_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_input10_I inst[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6293__B _2153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8064__I _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7377__A2 _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6979_ _2064_ _2866_ _2867_ _2017_ _2868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8718_ _4250_ _4244_ _4251_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8649_ reg_file.reg_storage\[8\]\[9\] _4203_ _4204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5129__S _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6468__B _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7301__A2 _3136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9054__A2 _4457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5863__A2 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6812__A1 _2684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8903__S _4366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5226__S1 _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5551__A1 _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4677__I _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6000_ _1544_ _0851_ _1914_ _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5854__A2 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9045__A2 _4407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I inst[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7951_ _3722_ _3740_ _3741_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7882_ net110 _3661_ _3678_ _3680_ _3681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_77_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _2585_ _2792_ _2793_ _2492_ _2794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5301__I _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6833_ _2725_ _2726_ _2727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9621_ _0407_ clknet_leaf_23_clk reg_file.reg_storage\[1\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7359__A2 _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9552_ _0338_ clknet_leaf_68_clk reg_file.reg_storage\[10\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _2463_ _2423_ _2655_ _2660_ _2661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_8503_ reg_file.reg_storage\[13\]\[24\] _4070_ _4107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5715_ _1630_ _1622_ _1631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8859__A2 _4338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _1601_ _2398_ _2565_ _2594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9483_ _0269_ clknet_leaf_2_clk reg_file.reg_storage\[8\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8434_ _4007_ _4061_ _4064_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5646_ reg_file.reg_storage\[4\]\[20\] reg_file.reg_storage\[5\]\[20\] reg_file.reg_storage\[6\]\[20\]
+ reg_file.reg_storage\[7\]\[20\] _1428_ _1422_ _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_98_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6132__I _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7531__A2 _3346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5577_ _1462_ _1492_ _1493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8365_ _4023_ _4024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5542__A1 _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8296_ _3969_ _3970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7316_ _3050_ _3157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input58_I mem_ld_dat[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4587__I _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7247_ _3091_ _3093_ _3094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5845__A2 _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7178_ _3031_ _3032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7598__A2 _3417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6129_ _2027_ _2033_ _2042_ _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5153__S0 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5208__S1 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__I1 reg_file.reg_storage\[13\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7589__A2 _3408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7601__I _3420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5500_ _1414_ _1415_ _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_27_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6480_ _2288_ _2380_ _2385_ _2386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_43_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7513__A2 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5524__A1 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5431_ _1344_ _1346_ _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_77_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8150_ _3866_ _3872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_10_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5362_ _1277_ _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7101_ net108 _2983_ _2980_ net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_93_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8081_ _3829_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7667__I3 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5293_ reg_file.reg_storage\[2\]\[9\] reg_file.reg_storage\[3\]\[9\] _0638_ _1209_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7032_ _2029_ _2918_ _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5827__A2 _1742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9018__A2 _4435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7029__A1 _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8983_ _4416_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6127__I _2040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7934_ reg_file.reg_storage\[5\]\[27\] _3720_ _3727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7865_ net107 _3661_ _3663_ _3665_ _3666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_7796_ net38 net47 _3412_ _3602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4870__I _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ _2061_ _2710_ _2026_ _2711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9604_ _0390_ clknet_leaf_19_clk reg_file.reg_storage\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5063__I0 _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5763__A1 _1604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6747_ _0969_ _2644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9535_ _0321_ clknet_leaf_123_clk reg_file.reg_storage\[10\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9466_ _0252_ clknet_leaf_97_clk reg_file.reg_storage\[12\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6678_ _2304_ _2578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9173__I _4511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8417_ reg_file.reg_storage\[14\]\[22\] _4024_ _4055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9397_ _0183_ clknet_leaf_20_clk reg_file.reg_storage\[14\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5629_ reg_file.reg_storage\[8\]\[23\] reg_file.reg_storage\[9\]\[23\] reg_file.reg_storage\[10\]\[23\]
+ reg_file.reg_storage\[11\]\[23\] _1471_ _1465_ _1545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_21_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8348_ _4009_ _4010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output164_I net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8279_ _3610_ _3957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_53_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5206__I _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9009__A2 _4424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5677__S1 _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7743__A2 _3146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__S1 _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5317__S _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__I2 reg_file.reg_storage\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6482__A2 _1832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4955__I _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5980_ _1871_ _1894_ _1895_ _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_144_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5993__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4931_ net79 _0798_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_118_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4862_ _0632_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8162__I _3867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7650_ _3069_ _3464_ _3465_ _3466_ _3467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__4690__I net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7734__A2 _3544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6601_ _2288_ _2503_ _2504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9320_ _0106_ clknet_leaf_49_clk reg_file.reg_storage\[6\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4793_ _0698_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7581_ _3034_ _3401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_27_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6532_ _2259_ _2422_ _2436_ _2437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _2289_ _2361_ _2369_ _2370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_70_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9251_ _0037_ clknet_leaf_3_clk reg_file.reg_storage\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput100 net100 mem_addr[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9182_ _4510_ _4536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8202_ _3705_ _3862_ _3901_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6170__A1 _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5414_ reg_file.reg_storage\[12\]\[1\] reg_file.reg_storage\[13\]\[1\] reg_file.reg_storage\[14\]\[1\]
+ reg_file.reg_storage\[15\]\[1\] _0770_ _1271_ _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput122 net122 mem_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput111 net111 mem_addr[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput133 net133 mem_ld_mask[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_140_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8133_ _3746_ _3854_ _3858_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6394_ _1252_ _1772_ _2303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput166 net166 mem_st_en vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput144 net144 mem_st_dat[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput155 net155 mem_st_dat[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_140_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5026__I _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5345_ reg_file.reg_storage\[8\]\[6\] reg_file.reg_storage\[9\]\[6\] reg_file.reg_storage\[10\]\[6\]
+ reg_file.reg_storage\[11\]\[6\] _0860_ _0837_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_2_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput177 net177 pc_next[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8064_ _3815_ _3819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5276_ _0835_ _1190_ _1191_ _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput199 net199 pc_next[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput188 net188 pc_next[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5356__S0 _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4865__I _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7015_ _2180_ _2849_ _2902_ _2351_ _2903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5108__S0 _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6225__A2 _2137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7422__A1 _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8966_ reg_file.reg_storage\[9\]\[31\] _4355_ _4403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5659__S1 _1537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7917_ _3400_ _3710_ _3711_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5984__A1 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8897_ reg_file.reg_storage\[9\]\[1\] _4363_ _4364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7848_ _3600_ _3649_ _3650_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7779_ _3586_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9518_ _0304_ clknet_leaf_60_clk reg_file.reg_storage\[11\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9449_ _0235_ clknet_leaf_51_clk reg_file.reg_storage\[12\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7489__A1 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7661__B2 _3476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7661__A1 net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7964__A2 _3751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A2 _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7716__A2 _3527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8710__I _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_8_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 inst[20] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6431__S _2183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput35 mem_ld_dat[11] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 mem_ld_dat[21] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput24 inst[30] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput57 mem_ld_dat[31] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput68 pc[12] net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput79 pc[22] net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6152__A1 _1789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5130_ net81 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_20_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4685__I _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5061_ _0509_ _0976_ net236 _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8093__S _3821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8820_ _4317_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8751_ _4274_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5963_ _1400_ _1403_ _1405_ _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7702_ _3513_ _3514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4914_ _0695_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8682_ reg_file.reg_storage\[8\]\[19\] _4223_ _4227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8821__S _4316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5894_ _1809_ _1810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_23_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7633_ net55 net34 _3412_ _3451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4845_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8380__A2 _4026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8620__I _4179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7564_ _3075_ _3384_ _3385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4776_ _0674_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9303_ _0089_ clknet_leaf_81_clk reg_file.reg_storage\[2\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6515_ _2130_ _2102_ _2179_ _2420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7495_ _1046_ _3304_ _3322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_101_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9234_ _0020_ clknet_leaf_79_clk reg_file.reg_storage\[5\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6446_ _1744_ _2157_ _2353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_9165_ reg_file.reg_storage\[15\]\[10\] _3556_ _4522_ _4527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8268__S _3941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6377_ _2079_ _2108_ _2179_ _2286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9096_ reg_file.reg_storage\[4\]\[16\] _4475_ _4484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5328_ reg_file.reg_storage\[2\]\[7\] reg_file.reg_storage\[3\]\[7\] _0755_ _1244_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8116_ reg_file.reg_storage\[2\]\[23\] _3817_ _3849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input40_I mem_ld_dat[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8047_ reg_file.reg_storage\[3\]\[30\] _3756_ _3805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8067__I _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6446__A2 _2157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5259_ _1165_ _0937_ _1174_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_110_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output127_I net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8199__A2 _3868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7946__A2 _3505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8949_ _4234_ _4363_ _4393_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5568__S0 _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7882__A1 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7882__B2 _3680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5660__A3 _1575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5948__A1 _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8440__I _4067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8362__A2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ reg_file.reg_storage\[12\]\[4\] reg_file.reg_storage\[13\]\[4\] reg_file.reg_storage\[14\]\[4\]
+ reg_file.reg_storage\[15\]\[4\] _0513_ _0514_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_37_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8114__A2 _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _1919_ _1932_ _2062_ _2211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4561_ _0484_ _0486_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_123_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7280_ _3113_ _3116_ _3124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__A1 _2038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6231_ _2121_ _1902_ _1946_ _2144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_21_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6162_ _1348_ _2076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5113_ _1028_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__6428__A2 _2335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7720__S _3492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6093_ _2006_ _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5044_ _0954_ _0955_ _0956_ _0959_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6844__B _2737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8803_ _4252_ _4257_ _4303_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7928__A2 _3719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8050__A1 _3751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6995_ _2879_ _2882_ _2883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ _1860_ _1861_ _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6135__I _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8734_ _4177_ _4262_ _4264_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8665_ reg_file.reg_storage\[8\]\[14\] _4203_ _4215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6739__I0 _2586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5877_ _1782_ _0726_ _1792_ _0678_ _1793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_36_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7616_ net44 net64 net41 net50 _3433_ _3434_ _3435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_47_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4828_ _0743_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8596_ reg_file.reg_storage\[12\]\[27\] _4162_ _4165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5798__S0 _1607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5167__A2 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input88_I pc[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8105__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7547_ _3344_ net86 _3356_ _3369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4759_ _0489_ _0511_ _0673_ _0674_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_43_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7478_ _3248_ net113 _3306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6667__A2 _2566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9217_ _0003_ clknet_leaf_126_clk reg_file.reg_storage\[5\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6429_ _2028_ _2336_ _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7864__A1 _3446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9148_ _4517_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9079_ _4474_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6419__A2 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5890__A3 _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7092__A2 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5722__S0 _1614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5150__S _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_50_clk_I clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_65_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9091__I _4461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7607__A1 _3424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5713__S0 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_123_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4963__I _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5800_ _1711_ _1713_ _1714_ _1715_ _1533_ _1536_ _1716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__8583__A2 _4154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6780_ _2671_ _2675_ _2676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5731_ _1586_ _1637_ _1646_ _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_clkbuf_leaf_18_clk_I clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5641__I0 _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5662_ _0849_ _1577_ _1578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6346__A1 _2135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8450_ reg_file.reg_storage\[13\]\[1\] _4076_ _4077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8381_ _3938_ _4025_ _4034_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5593_ _1009_ _1508_ _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7401_ _3209_ net105 _3236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4613_ reg_file.reg_storage\[8\]\[3\] reg_file.reg_storage\[9\]\[3\] reg_file.reg_storage\[10\]\[3\]
+ reg_file.reg_storage\[11\]\[3\] _0534_ _0535_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_25_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7332_ _3159_ _3171_ _3172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7263_ _3105_ _3108_ _3109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9002_ reg_file.reg_storage\[1\]\[11\] _3567_ _4421_ _4427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6214_ _2006_ _1954_ _2127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7861__A4 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7194_ _3045_ _3046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_110_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5034__I _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6145_ _2044_ _2059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_127_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7074__A2 _2550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6076_ _1310_ _1989_ _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5027_ reg_file.reg_storage\[1\]\[18\] _0941_ _0942_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5180__S1 _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8717_ reg_file.reg_storage\[8\]\[30\] _4173_ _4251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6978_ _2005_ _2754_ _2867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5929_ _1843_ _1844_ _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8648_ _4180_ _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8579_ _3974_ _4154_ _4155_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output194_I net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4899__A1 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__A2 _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8456__S _4079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8255__I _3509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6879__A2 _2450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5000__A1 _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6500__A1 _2404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7950_ reg_file.reg_storage\[5\]\[29\] _3720_ _3741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5457__I3 _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4814__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6901_ _2137_ _2588_ _2793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7881_ _3671_ _3277_ _3499_ _3679_ _3680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6832_ _2720_ _2723_ _2726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8556__A2 _4128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9620_ _0406_ clknet_leaf_22_clk reg_file.reg_storage\[1\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9551_ _0337_ clknet_leaf_64_clk reg_file.reg_storage\[10\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8308__A2 _3975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6763_ _2324_ _2659_ _2210_ _2660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5714_ _1624_ _1626_ _1628_ _1629_ _1531_ _1235_ _1630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_6694_ _1862_ _2593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8502_ _3987_ _4076_ _4106_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9482_ _0268_ clknet_leaf_3_clk reg_file.reg_storage\[8\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8433_ reg_file.reg_storage\[14\]\[29\] _4059_ _4064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5645_ reg_file.reg_storage\[12\]\[20\] reg_file.reg_storage\[13\]\[20\] reg_file.reg_storage\[14\]\[20\]
+ reg_file.reg_storage\[15\]\[20\] _1463_ _1422_ _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_98_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ _1484_ _1488_ _1490_ _1491_ _1455_ _1438_ _1492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_8364_ _4022_ _4023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5542__A2 _1457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8295_ _3656_ _3969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4868__I _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7315_ _3154_ _3155_ _3156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7246_ _3092_ _3084_ _3093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7177_ _2975_ _1901_ _3031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6128_ _2036_ _1323_ _2039_ _2041_ _2042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5699__I _1614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5153__S1 _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6059_ _1972_ _1973_ _1974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_107_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8547__A2 _4129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4664__S0 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5230__A1 _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8914__S _4372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8713__I _3739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4655__S0 _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5430_ _0729_ _1345_ _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5524__A2 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5361_ _1272_ _1274_ _1275_ _1276_ _0625_ _0823_ _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_7100_ net97 _2982_ _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_93_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5292_ reg_file.reg_storage\[4\]\[9\] reg_file.reg_storage\[5\]\[9\] reg_file.reg_storage\[6\]\[9\]
+ reg_file.reg_storage\[7\]\[9\] _0919_ _0856_ _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8080_ reg_file.reg_storage\[2\]\[7\] _3511_ _3828_ _3829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7031_ _1929_ _1922_ _2918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7029__A2 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8777__A2 _4288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7013__B _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8982_ reg_file.reg_storage\[1\]\[2\] _3455_ _4415_ _4416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5312__I _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7933_ _3725_ _3726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8623__I _3454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7864_ _3446_ _3664_ _3665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7795_ _3472_ _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_93_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6815_ _2606_ _2709_ _2101_ _2710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9603_ _0389_ clknet_leaf_136_clk reg_file.reg_storage\[1\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9534_ _0320_ clknet_4_13_0_clk reg_file.reg_storage\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6746_ _2115_ _2571_ _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5763__A2 _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6960__A1 _2841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9465_ _0251_ clknet_leaf_96_clk reg_file.reg_storage\[12\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6677_ _2576_ _2577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8416_ _3981_ _4051_ _4054_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9396_ _0182_ clknet_leaf_28_clk reg_file.reg_storage\[14\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6712__A1 _1635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5628_ _0874_ _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input70_I pc[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8347_ _3745_ _4009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5559_ _1462_ _1474_ _1475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_60_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8278_ _3956_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5279__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output157_I net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7229_ _3076_ _3077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8768__A2 _4275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6228__B1 _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8533__I _4127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9193__A2 _4538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8940__A2 _4386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4637__S0 _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_130_clk clknet_4_5_0_clk clknet_leaf_130_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_122_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7259__A2 _3090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4580__I3 reg_file.reg_storage\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_4_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4930_ _0845_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4861_ _0765_ _0766_ _0769_ _0776_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__9184__A2 _4531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7195__A1 _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6600_ _2366_ _2502_ _2185_ _2503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7580_ _3399_ _3400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4792_ _0600_ _0605_ _0613_ _0608_ _0707_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_6531_ _2193_ _2431_ _2435_ _2436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6462_ _2333_ _2368_ _2369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9250_ _0036_ clknet_leaf_19_clk reg_file.reg_storage\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_121_clk clknet_4_7_0_clk clknet_leaf_121_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7498__A2 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput101 net101 mem_addr[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9181_ _3966_ _4531_ _4535_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8201_ reg_file.reg_storage\[6\]\[24\] _3863_ _3901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6393_ _2261_ _2301_ _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8819__S _4316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5413_ _1326_ _0624_ _1327_ _1328_ _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput123 net123 mem_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput112 net112 mem_addr[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput134 net134 mem_st_dat[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8132_ reg_file.reg_storage\[2\]\[30\] _3811_ _3858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5344_ reg_file.reg_storage\[12\]\[6\] reg_file.reg_storage\[13\]\[6\] reg_file.reg_storage\[14\]\[6\]
+ reg_file.reg_storage\[15\]\[6\] _0860_ _0837_ _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput167 net167 mem_st_mask[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput156 net156 mem_st_dat[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput145 net145 mem_st_dat[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_130_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8618__I _4180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8998__A2 _4424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8063_ _3817_ _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5275_ net67 _0888_ _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput178 net178 pc_next[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput189 net189 pc_next[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5356__S1 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7522__I _1511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7014_ _0996_ _1890_ _2900_ _2901_ _2902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_128_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5042__I _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5108__S1 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8965_ _4250_ _4398_ _4402_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4867__S0 _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5433__A1 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7916_ reg_file.reg_storage\[5\]\[25\] _3422_ _3711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8896_ _4359_ _4363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9175__A2 _4531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7847_ reg_file.reg_storage\[5\]\[17\] _3544_ _3650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5292__S0 _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7778_ reg_file.reg_storage\[5\]\[12\] _3585_ _3569_ _3586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6729_ _2564_ _2626_ _2627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9517_ _0303_ clknet_leaf_12_clk reg_file.reg_storage\[11\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5926__B _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9448_ _0234_ clknet_leaf_48_clk reg_file.reg_storage\[12\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_112_clk clknet_4_13_0_clk clknet_leaf_112_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7489__A2 _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8438__A1 _4013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9379_ _0165_ clknet_leaf_136_clk reg_file.reg_storage\[14\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7110__A1 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7413__A2 net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8263__I _3945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6924__A1 _2404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5328__S _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput36 mem_ld_dat[12] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_103_clk clknet_4_15_0_clk clknet_leaf_103_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput14 inst[21] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput25 inst[31] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput58 mem_ld_dat[3] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput47 mem_ld_dat[22] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput69 pc[13] net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_122_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8429__A1 reg_file.reg_storage\[14\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7101__A1 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5063__S _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5060_ _0975_ _0709_ _0710_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8374__S _4029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7404__A2 _1603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8750_ reg_file.reg_storage\[11\]\[8\] _4200_ _4272_ _4274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_88_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5962_ _1406_ _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7701_ _1709_ _0714_ _2986_ _3513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4913_ _0828_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5966__A2 _1457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8681_ _4187_ _4226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5893_ _1251_ _1809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_23_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7632_ _3405_ _3449_ _3450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_118_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4844_ _0759_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7563_ net89 _3383_ _3384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_16_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4775_ _0673_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_133_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9302_ _0088_ clknet_leaf_116_clk reg_file.reg_storage\[2\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6514_ _2415_ _2418_ _2419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9233_ _0019_ clknet_leaf_70_clk reg_file.reg_storage\[5\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7494_ _3319_ _3320_ _3321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6445_ _2351_ _2352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9164_ _3945_ _4512_ _4526_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6376_ _2098_ _2111_ _2003_ _2285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8348__I _4009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8115_ _3689_ _3844_ _3848_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5327_ reg_file.reg_storage\[4\]\[7\] reg_file.reg_storage\[5\]\[7\] reg_file.reg_storage\[6\]\[7\]
+ reg_file.reg_storage\[7\]\[7\] _0633_ _0642_ _1243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_9095_ _4483_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4876__I _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8046_ _3740_ _3801_ _3804_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input33_I mem_ld_dat[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5258_ _0800_ _1173_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_110_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5189_ _0510_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_97_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5406__A1 _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8948_ reg_file.reg_storage\[9\]\[23\] _4361_ _4393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7159__A1 _3019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7159__B2 _1664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8879_ _4246_ _4348_ _4350_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8811__I _4309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__S1 _1483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7882__A2 _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5611__S _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6950__B _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5256__S0 _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4560_ _0485_ net16 net17 _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_37_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7873__A2 _3262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6230_ _2134_ _2142_ _1948_ _2143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_110_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6161_ _2074_ _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5112_ _1013_ _1027_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5636__A1 _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6092_ _1977_ _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5487__I1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5043_ _0957_ reg_file.reg_storage\[2\]\[19\] _0958_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8802_ reg_file.reg_storage\[11\]\[31\] _4255_ _4303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8832__S _4322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6994_ _1521_ _2881_ _2882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5320__I net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ _0891_ _0907_ _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8733_ reg_file.reg_storage\[11\]\[1\] _4263_ _4264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8664_ _4181_ _4214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6739__I1 _2636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8631__I _3477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5876_ _1253_ _1784_ _1785_ _1791_ _1792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_36_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7615_ _3023_ _3434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ _0736_ _0741_ _0742_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_7_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8595_ _4120_ _4164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5798__S1 _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6151__I _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7546_ net88 _3368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4758_ _0667_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_114_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4689_ _0597_ _0600_ _0605_ net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7477_ net81 _3304_ _3305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA_clkbuf_4_12_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9216_ _0002_ clknet_leaf_129_clk reg_file.reg_storage\[5\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6428_ _1810_ _2335_ _1229_ _2336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_112_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9147_ reg_file.reg_storage\[15\]\[2\] _3455_ _4516_ _4517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6359_ _2170_ _2269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9078_ reg_file.reg_storage\[4\]\[8\] _3530_ _4472_ _4474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8029_ reg_file.reg_storage\[3\]\[22\] _3764_ _3795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_141_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5722__S1 _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8041__A2 _3799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6355__A2 _2264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8804__A1 _3809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7607__A2 _3425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8716__I _3745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5713__S1 _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6236__I _2148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8652__S _4198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8032__A2 _3766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5477__S0 _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ _0734_ _1645_ _1646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5661_ _0672_ _1568_ _1576_ _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_72_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7400_ _3233_ _3234_ _3235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_111_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8380_ reg_file.reg_storage\[14\]\[6\] _4026_ _4034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5592_ _1417_ _1498_ _1507_ _1508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_4_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4612_ _0482_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_142_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7331_ _3154_ _3161_ _3171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7262_ _3092_ _3084_ _3107_ _3108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_1_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9001_ _1197_ _4406_ _4426_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6213_ _2079_ _2119_ _2125_ _2126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5857__A1 _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7193_ _3044_ _3045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6144_ _2000_ _2025_ _2055_ _2057_ _2058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_0_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _0979_ _1988_ _1989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_127_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ _0856_ _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_92_clk clknet_4_14_0_clk clknet_leaf_92_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8023__A2 _3789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__I _1900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6977_ _2030_ _2817_ _2865_ _2866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8716_ _3745_ _4250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ _1555_ _1844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8647_ _3542_ _4202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6337__A2 _2032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5859_ _1761_ _1764_ _1774_ _1775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_138_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8578_ reg_file.reg_storage\[12\]\[19\] _4152_ _4155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output187_I net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7529_ _3350_ _3352_ _3353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5225__I _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8737__S _4266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7641__S _3458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9211__A1 _4009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8472__S _4085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_83_clk clknet_4_14_0_clk clknet_leaf_83_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6025__A1 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7773__A1 _1692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6500__A2 _2405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8253__A2 _3924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4814__A2 _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9202__A1 _3995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_74_clk clknet_4_9_0_clk clknet_leaf_74_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6900_ _2245_ _2691_ _2791_ _2792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7880_ _3278_ _3645_ _3679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6831_ _2404_ _2725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_18_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9550_ _0336_ clknet_leaf_60_clk reg_file.reg_storage\[10\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6567__A2 _2470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_75_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8501_ reg_file.reg_storage\[13\]\[23\] _4074_ _4106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6762_ _2548_ _2658_ _2101_ _2659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9481_ _0267_ clknet_leaf_52_clk reg_file.reg_storage\[8\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5713_ reg_file.reg_storage\[4\]\[17\] reg_file.reg_storage\[5\]\[17\] reg_file.reg_storage\[6\]\[17\]
+ reg_file.reg_storage\[7\]\[17\] _0658_ _1627_ _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6693_ _2592_ net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_72_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7516__A1 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8432_ _4004_ _4061_ _4063_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5644_ reg_file.reg_storage\[1\]\[20\] _1559_ _1422_ _1560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_98_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5622__S0 _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8363_ _3865_ _4021_ _4022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5575_ reg_file.reg_storage\[8\]\[30\] reg_file.reg_storage\[9\]\[30\] reg_file.reg_storage\[10\]\[30\]
+ reg_file.reg_storage\[11\]\[30\] _1482_ _1483_ _1491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7314_ _3145_ _3133_ _3155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8294_ _3967_ _3959_ _3968_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8557__S _4138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5045__I _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7245_ _3078_ _3081_ _3092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7176_ net108 _3030_ _2971_ net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6127_ _2040_ _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_99_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _0721_ _1783_ _1973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_65_clk clknet_4_11_0_clk clknet_leaf_65_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_64_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5009_ _0906_ _0918_ _0924_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_107_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output102_I net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6558__A2 _2461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7755__A1 _3484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9679_ _0465_ clknet_leaf_54_clk reg_file.reg_storage\[15\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_79_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4664__S1 _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8180__A1 _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8467__S _4085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5836__A4 _1751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8235__A2 _3923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__A1 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_56_clk clknet_4_10_0_clk clknet_leaf_56_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_69_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8930__S _4365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4655__S1 _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_0_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4969__I _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5524__A3 _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7345__I _3183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5360_ reg_file.reg_storage\[8\]\[5\] reg_file.reg_storage\[9\]\[5\] reg_file.reg_storage\[10\]\[5\]
+ reg_file.reg_storage\[11\]\[5\] _0637_ _0634_ _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_93_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5291_ net96 _0749_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7030_ _2036_ _2864_ _2917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5288__A2 _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8226__A2 _3915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8981_ _4414_ _4415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7948__C _3738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7932_ net116 _3698_ _3699_ _3723_ _3724_ _3725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_78_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5460__A2 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7588__I1 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7863_ _3401_ _3252_ _3439_ _3253_ _3664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7794_ _3427_ _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6424__I _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6814_ _2038_ _2707_ _2708_ _2709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9602_ _0388_ clknet_leaf_19_clk reg_file.reg_storage\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9533_ _0319_ clknet_leaf_108_clk reg_file.reg_storage\[11\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6745_ _2615_ _2620_ _2642_ net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_9464_ _0250_ clknet_leaf_89_clk reg_file.reg_storage\[12\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_102_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8415_ reg_file.reg_storage\[14\]\[21\] _4049_ _4054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6676_ _2167_ _2576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9395_ _0181_ clknet_leaf_75_clk reg_file.reg_storage\[14\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6712__A2 _2171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5627_ _0828_ _1542_ _1543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input63_I mem_ld_dat[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8346_ _4007_ _4001_ _4008_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5558_ _1466_ _1470_ _1472_ _1473_ _1437_ _1438_ _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_8277_ reg_file.reg_storage\[7\]\[13\] _3955_ _3927_ _3956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5489_ _1378_ _1397_ _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5279__A2 _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7228_ _3075_ _3076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7159_ _3019_ _3018_ _3017_ _1664_ _2994_ net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__5503__I _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6228__A1 _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6228__B2 _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8814__I _4309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_38_clk clknet_4_2_0_clk clknet_leaf_38_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8750__S _4272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__S0 _1590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6400__B2 _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6400__A1 _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4789__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6703__A2 _2368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8925__S _4365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7967__A1 _3753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4860_ _0773_ reg_file.reg_storage\[2\]\[20\] _0775_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__S0 _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6530_ _2432_ _1835_ _2173_ _2434_ _2435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_7_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4791_ _0597_ _0599_ _0611_ _0664_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_28_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6461_ _2362_ _2223_ _2367_ _2368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_141_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9180_ reg_file.reg_storage\[15\]\[17\] _4525_ _4535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8200_ _3696_ _3870_ _3900_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6392_ _2145_ _2300_ _2185_ _2301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5412_ reg_file.reg_storage\[2\]\[1\] _0771_ _0624_ _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput124 net124 mem_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput102 net102 mem_addr[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput113 net113 mem_addr[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_140_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8131_ _3740_ _3854_ _3857_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5343_ _1256_ _0807_ _1257_ _1258_ _1259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_51_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput168 net168 mem_st_mask[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput135 net135 mem_st_dat[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput146 net146 mem_st_dat[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput157 net157 mem_st_dat[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_130_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6458__A1 _2018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8062_ _3816_ _3817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5274_ _1189_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput179 net179 pc_next[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7013_ _2879_ _1521_ _2168_ _2173_ _2901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__8634__I _3489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8964_ reg_file.reg_storage\[9\]\[30\] _4355_ _4402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4867__S1 _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7915_ _3709_ _3710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8895_ _4361_ _4362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7846_ _3648_ _3649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7186__A2 _3037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4989_ reg_file.reg_storage\[8\]\[17\] reg_file.reg_storage\[9\]\[17\] reg_file.reg_storage\[10\]\[17\]
+ reg_file.reg_storage\[11\]\[17\] _0861_ _0893_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_92_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6933__A2 _2370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7777_ _3584_ _3585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9516_ _0302_ clknet_leaf_64_clk reg_file.reg_storage\[11\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8135__A1 _3751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5292__S1 _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6728_ _1600_ _1863_ _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4603__S _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8686__A2 _4226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9447_ _0233_ clknet_leaf_34_clk reg_file.reg_storage\[12\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6659_ _2532_ _2540_ _2559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9378_ _0164_ clknet_leaf_4_clk reg_file.reg_storage\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8329_ _3718_ _3995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5807__S0 _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput37 mem_ld_dat[13] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput26 inst[3] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput15 inst[22] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput59 mem_ld_dat[4] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 mem_ld_dat[23] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5408__I net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8719__I _3750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8655__S _4198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5112__A1 _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6860__A1 _2122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5961_ _1085_ _1376_ _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8390__S _4035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8680_ _3666_ _4225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7700_ _3512_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4912_ _0799_ _0827_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7631_ _3447_ _3028_ _3448_ _3449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_114_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5892_ _1761_ _1806_ _1807_ _1808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4843_ _0640_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4774_ _0488_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7562_ _3344_ net86 _3368_ _3356_ _3383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_28_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9301_ _0087_ clknet_leaf_24_clk reg_file.reg_storage\[2\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6513_ _2417_ _2405_ _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7493_ _3309_ _3313_ _3307_ _3320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_114_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7961__C _3749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9232_ _0018_ clknet_leaf_32_clk reg_file.reg_storage\[5\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6444_ _1907_ _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_9_clk clknet_4_6_0_clk clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9163_ reg_file.reg_storage\[15\]\[9\] _4525_ _4526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6375_ _2189_ _2284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_3_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5351__A1 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9093__A2 _4481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8114_ reg_file.reg_storage\[2\]\[22\] _3817_ _3848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9094_ reg_file.reg_storage\[4\]\[15\] _3623_ _4465_ _4483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5326_ _1183_ _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8045_ reg_file.reg_storage\[3\]\[29\] _3799_ _3804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5103__A1 _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5257_ _1166_ _1170_ _1171_ _1172_ _0822_ _0825_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__5053__I _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5188_ _1045_ _1102_ _1103_ _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_3_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input26_I inst[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8947_ _4232_ _4388_ _4392_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5406__A2 _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8878_ reg_file.reg_storage\[10\]\[28\] _4346_ _4350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8356__A1 _3809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7829_ _3626_ _3632_ _3539_ _3633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5965__I0 _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8903__I0 reg_file.reg_storage\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7331__A2 _3161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7398__A2 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8898__A2 _4362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5256__S1 _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4977__I _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6530__B1 _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6160_ _2073_ _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8385__S _4035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5111_ _1014_ _1026_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6833__A1 _2725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6091_ _2004_ _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_109_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5042_ _0763_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8801_ _4250_ _4298_ _4302_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8586__A1 reg_file.reg_storage\[12\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7389__A2 net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6993_ _2836_ _2857_ _2880_ _2881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8732_ _4259_ _4263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5944_ net73 _0889_ _1860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8663_ _3610_ _4213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5875_ _1119_ _1786_ _1790_ _1791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7614_ _3411_ _3433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8594_ _3996_ _4121_ _4163_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4826_ _0555_ _0671_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7545_ _3045_ _3364_ _3366_ _3324_ _3367_ net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_28_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5048__I _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4757_ _0666_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4688_ _0604_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7476_ net79 net80 _3274_ _3304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8359__I _4016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4887__I _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9215_ _0001_ clknet_leaf_18_clk reg_file.reg_storage\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6427_ _1924_ _2335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_112_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6358_ _2167_ _2268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9146_ _4515_ _4516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_8_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5875__A2 _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5309_ _1224_ _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9077_ _4473_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5627__A2 _1542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6289_ _2140_ _2200_ _2201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6824__B2 _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8028_ _3682_ _3791_ _3794_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6607__I _1955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5667__B net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7552__A2 _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__A2 _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8804__A2 _4171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__S1 _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8732__I _4259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5660_ _1445_ _1385_ _1575_ _1576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_57_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ _0513_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_143_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4988__S0 _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5554__A1 _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5591_ _1351_ _1506_ _1507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7330_ _3139_ _3147_ _3169_ _3148_ _3170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_13_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7083__I _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7261_ _3091_ _3106_ _3107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6354__I0 _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9000_ _3556_ _4405_ _4426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5857__A2 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6212_ _2117_ _1945_ _2124_ _2125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7192_ _3039_ _3044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6143_ _2056_ _2057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__9004__S _4421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5165__S0 _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6806__A1 _2684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6074_ _1182_ _0694_ _1903_ _0730_ _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_5025_ reg_file.reg_storage\[2\]\[18\] reg_file.reg_storage\[3\]\[18\] _0940_ _0941_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8843__S _4315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6976_ _2008_ _2864_ _2865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7231__A1 _3058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8715_ _4248_ _4244_ _4249_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5927_ _1544_ _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8646_ _4201_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input93_I pc[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7534__A2 net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5858_ _1767_ _1768_ _1773_ _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_138_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8577_ _4132_ _4154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5789_ _1584_ _1705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4809_ _0703_ _0724_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7528_ _3338_ _3351_ _3336_ _3352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7459_ _3270_ _3287_ _3288_ _3289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_31_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5848__A2 _1763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9129_ _4009_ _4498_ _4502_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8817__I _4309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7470__A1 _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__S0 _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8722__A1 _3754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7525__A2 _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_80_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7289__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4990__I _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6830_ _2720_ _2723_ _2724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_18_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5075__I0 reg_file.reg_storage\[12\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6761_ _2012_ _2604_ _2657_ _2658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5712_ reg_file.reg_storage\[12\]\[17\] reg_file.reg_storage\[13\]\[17\] reg_file.reg_storage\[14\]\[17\]
+ reg_file.reg_storage\[15\]\[17\] _0658_ _1627_ _1628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_92_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8500_ _3984_ _4101_ _4105_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9480_ _0266_ clknet_leaf_56_clk reg_file.reg_storage\[8\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6692_ _2569_ _2572_ _2581_ _2591_ _2592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_8431_ reg_file.reg_storage\[14\]\[28\] _4059_ _4063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5643_ reg_file.reg_storage\[2\]\[20\] reg_file.reg_storage\[3\]\[20\] _1369_ _1559_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_98_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5574_ reg_file.reg_storage\[12\]\[30\] reg_file.reg_storage\[13\]\[30\] reg_file.reg_storage\[14\]\[30\]
+ reg_file.reg_storage\[15\]\[30\] _1482_ _1489_ _1490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_98_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5622__S1 _1537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8362_ _3760_ net2 _4021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7313_ net67 _3154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8293_ reg_file.reg_storage\[7\]\[17\] _3947_ _3968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5386__S0 _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7244_ _3078_ _3081_ _3091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7175_ _2972_ net97 _3030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8637__I _3501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__S0 _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6126_ _2021_ _2040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6057_ _1795_ _1242_ _1972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5008_ _0906_ _0923_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_107_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6007__A2 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7204__A1 _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7755__A2 _3156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6959_ _2333_ _2570_ _2849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_64_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9678_ _0464_ clknet_leaf_62_clk reg_file.reg_storage\[15\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5518__A1 _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8629_ reg_file.reg_storage\[8\]\[3\] _4189_ _4187_ _4190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8180__A2 _3888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8748__S _4272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6067__I _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7443__A1 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__A2 _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__8483__S _4078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_82_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9120__A1 _3995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8658__S _4186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5290_ _1194_ _0951_ _1205_ _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5368__S0 _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8980_ _4409_ _4414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5540__S0 _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5996__A1 _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7931_ _3702_ _3342_ _3496_ _1416_ _3724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_89_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7862_ _3640_ _3662_ _3652_ _3663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_77_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9601_ _0387_ clknet_leaf_126_clk reg_file.reg_storage\[1\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5748__A1 _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7793_ _3599_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6813_ _2122_ _2656_ _2708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9532_ _0318_ clknet_leaf_101_clk reg_file.reg_storage\[11\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6744_ _2631_ _2633_ _2640_ _2641_ _2642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_58_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9463_ _0249_ clknet_leaf_89_clk reg_file.reg_storage\[12\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_102_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6675_ _2573_ _2562_ _2575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8414_ _3978_ _4051_ _4053_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5626_ _1541_ _1542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7536__I net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9394_ _0180_ clknet_leaf_75_clk reg_file.reg_storage\[14\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8345_ reg_file.reg_storage\[7\]\[29\] _3997_ _4008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5557_ reg_file.reg_storage\[8\]\[31\] reg_file.reg_storage\[9\]\[31\] reg_file.reg_storage\[10\]\[31\]
+ reg_file.reg_storage\[11\]\[31\] _1464_ _1465_ _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__8568__S _4131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _1403_ _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5359__S0 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8276_ _3596_ _3955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input56_I mem_ld_dat[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7227_ _3040_ _3075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7673__A1 _3090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7158_ _3006_ net219 _3019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_67_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7089_ _2968_ _2971_ _2972_ _2973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6109_ _2019_ _2020_ _2022_ _2023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5739__A1 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5834__S1 _1642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6400__A2 _2283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7900__A2 _3458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6164__A1 _1947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_94_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_20_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8478__S _4078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4714__A2 _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7664__A1 _3428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7967__A2 _3754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__S1 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4790_ _0617_ _0615_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_129_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5589__S0 _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6155__A1 _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6460_ _2110_ _2366_ _2367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6391_ _2297_ _2222_ _2299_ _2300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5411_ reg_file.reg_storage\[3\]\[1\] _0628_ _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput125 net125 mem_addr[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput103 net103 mem_addr[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput114 net114 mem_addr[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_63_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8130_ reg_file.reg_storage\[2\]\[29\] _3852_ _3857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5342_ reg_file.reg_storage\[2\]\[6\] _0813_ _0774_ _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput136 net136 mem_st_dat[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput158 net158 mem_st_dat[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput147 net147 mem_st_dat[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_130_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8187__I _3867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8061_ _3815_ _3816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput169 net169 mem_st_mask[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_130_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7091__I _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5273_ _1184_ _1186_ _1187_ _1188_ _0964_ _0946_ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_7012_ _0996_ _1890_ _2374_ _2900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5761__S0 _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_78_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7958__A2 _3746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_121_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8963_ _4248_ _4398_ _4401_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6435__I _1734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7914_ net114 _3698_ _3699_ _3707_ _3708_ _3709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_8894_ _4360_ _4361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7845_ net105 _3601_ _3644_ _3647_ _3648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_77_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_136_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6394__A1 _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4988_ reg_file.reg_storage\[12\]\[17\] reg_file.reg_storage\[13\]\[17\] reg_file.reg_storage\[14\]\[17\]
+ reg_file.reg_storage\[15\]\[17\] _0861_ _0903_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_clkbuf_leaf_16_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9515_ _0301_ clknet_leaf_1_clk reg_file.reg_storage\[11\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7776_ _3583_ _3584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8135__A2 _3813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6727_ _2597_ _2622_ _2624_ _2560_ _2625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9446_ _0232_ clknet_leaf_42_clk reg_file.reg_storage\[12\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6658_ _2532_ _2540_ _2558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6697__A2 _2595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5609_ _1423_ _1352_ _1479_ _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9377_ _0163_ clknet_leaf_132_clk reg_file.reg_storage\[14\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8328_ _3993_ _3915_ _3994_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6589_ _2209_ _2492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output162_I net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8259_ _3529_ _3943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5450__S _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8761__S _4265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5807__S1 _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput27 inst[4] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput16 inst[23] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput38 mem_ld_dat[14] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput49 mem_ld_dat[24] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7885__A1 _3660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8735__I _4259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6860__A2 _2707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5960_ _1409_ _1441_ _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4911_ _0800_ _0826_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5891_ _1265_ _1760_ _1807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7630_ net42 _3433_ _3448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4842_ _0757_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_59_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7086__I _2969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8117__A2 _3819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4773_ _0682_ _0684_ _0688_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7561_ _3378_ _3379_ _3380_ _3382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9300_ _0086_ clknet_leaf_75_clk reg_file.reg_storage\[2\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6512_ _1959_ _2416_ _2417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7492_ _3316_ _3318_ _3319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6128__A1 _2036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9231_ _0017_ clknet_4_10_0_clk reg_file.reg_storage\[5\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6443_ _2350_ net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_82_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9162_ _4510_ _4525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6374_ _2279_ _2282_ _2283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_9093_ _3957_ _4481_ _4482_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8113_ _3682_ _3844_ _3847_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5325_ _1240_ _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8044_ _3734_ _3801_ _3803_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5256_ reg_file.reg_storage\[8\]\[15\] reg_file.reg_storage\[9\]\[15\] reg_file.reg_storage\[10\]\[15\]
+ reg_file.reg_storage\[11\]\[15\] _0802_ _0804_ _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_110_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5270__S _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5187_ _0979_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_143_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8946_ reg_file.reg_storage\[9\]\[22\] _4361_ _4392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input19_I inst[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8877_ _4243_ _4348_ _4349_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8356__A2 _4015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__S _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7828_ _3631_ _3632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_65_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6367__A1 _2231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7759_ _3567_ _3568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8108__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5965__I1 _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_50_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5590__A2 _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9429_ _0215_ clknet_leaf_20_clk reg_file.reg_storage\[13\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5342__A2 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5725__S0 _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4853__A1 _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8044__A1 _3734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5419__I _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7858__A1 _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6530__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5110_ _1015_ _1019_ _1023_ _1024_ _0965_ _1025_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_85_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6090_ _2003_ _2004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5041_ _0772_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5097__A1 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8800_ reg_file.reg_storage\[11\]\[30\] _4255_ _4302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8586__A2 _4127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6597__A1 _2494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6992_ _2856_ _2484_ _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8731_ _4261_ _4262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5943_ _0950_ _1858_ _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8662_ _4212_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5874_ _1787_ _1789_ _0719_ _1790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8593_ reg_file.reg_storage\[12\]\[26\] _4162_ _4163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7613_ _3431_ _3432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4825_ _0737_ _0728_ _0739_ _0740_ _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_7_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7544_ _3051_ net118 _3367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7849__A1 _3010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4756_ _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4687_ _0601_ _0602_ _0603_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_7475_ _3076_ _3294_ _3302_ _3226_ _3303_ net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_114_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9214_ _0000_ clknet_leaf_112_clk reg_file.reg_storage\[5\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6426_ _2037_ _1283_ _1266_ _2334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_31_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9145_ _4509_ _4515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_59_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6357_ _1938_ _2231_ _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_8_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5064__I _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5308_ _1219_ _1221_ _1222_ _1223_ _0821_ _0787_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__7077__A2 _2171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5088__A1 _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9076_ reg_file.reg_storage\[4\]\[7\] _3510_ _4472_ _4473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6288_ _2041_ _2197_ _2199_ _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5239_ _0863_ reg_file.reg_storage\[2\]\[14\] _0958_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8027_ reg_file.reg_storage\[3\]\[21\] _3789_ _3794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4835__A1 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output125_I net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8929_ _4213_ _4381_ _4382_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5260__A1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6760__A1 _2030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8501__A2 _4074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7454__I net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6512__A1 _1959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5079__A1 _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4826__A1 _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4610_ _0533_ net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
X_5590_ _1505_ _1462_ _1506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4988__S1 _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7260_ _3087_ _3090_ _3106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7191_ net65 _0689_ _3043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6211_ _2120_ _2123_ _2124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8396__S _4028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6142_ _1113_ _2056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5165__S1 _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6073_ _1902_ _1905_ _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_127_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _0628_ _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5490__A1 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ _1927_ _1930_ _2864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8714_ reg_file.reg_storage\[8\]\[29\] _4241_ _4249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6443__I _2350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5926_ _1813_ _1841_ _1651_ _1842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8645_ reg_file.reg_storage\[8\]\[8\] _4200_ _4198_ _4201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5857_ _1251_ _1772_ _1773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5059__I net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8576_ _3970_ _4147_ _4153_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6742__A1 _2463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5788_ _1582_ _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input86_I pc[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4808_ _0722_ _0716_ _0708_ _0723_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_133_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__I _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4739_ _0588_ _0598_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7527_ net84 _3335_ _3351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7458_ _3275_ _3278_ _3288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6409_ _2230_ _1771_ _2317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__5723__S _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7389_ _3208_ net104 _3060_ _3224_ _3225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9128_ reg_file.reg_storage\[4\]\[30\] _4455_ _4502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9059_ _4461_ _4462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5522__I _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7470__A2 _3138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5481__A1 _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__S1 _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5233__A1 _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8722__A2 _4171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4992__B1 _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7289__A2 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7461__A2 net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5224__A1 _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5075__I1 reg_file.reg_storage\[13\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6760_ _2030_ _2656_ _2657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_18_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6972__A1 _2841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5711_ _0535_ _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_114_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6691_ _2583_ _2590_ _2591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5808__S _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8430_ _4000_ _4061_ _4062_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5642_ reg_file.reg_storage\[8\]\[20\] reg_file.reg_storage\[9\]\[20\] reg_file.reg_storage\[10\]\[20\]
+ reg_file.reg_storage\[11\]\[20\] _1428_ _1451_ _1558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_98_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_rebuffer9_I _1742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8361_ _3912_ _4018_ _4020_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5573_ _1363_ _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7312_ _3035_ _2413_ _3144_ _3146_ _3153_ net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_13_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8292_ _3966_ _3967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7243_ _1382_ _1383_ _3090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7174_ _3024_ _3029_ net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_123_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8229__A1 _3424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6125_ _2038_ _1283_ _1296_ _2039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5138__S1 _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7452__A2 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6056_ _1299_ _1971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5007_ reg_file.reg_storage\[4\]\[16\] reg_file.reg_storage\[5\]\[16\] reg_file.reg_storage\[6\]\[16\]
+ reg_file.reg_storage\[7\]\[16\] _0921_ _0922_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_107_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7204__A2 _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5215__A1 _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_132_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_120_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6958_ _2176_ _2846_ _2847_ _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_64_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6963__A1 _2841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8704__A2 _4241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6889_ _2719_ _2718_ _2781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_9677_ _0463_ clknet_leaf_13_clk reg_file.reg_storage\[15\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5909_ _1193_ _1825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_106_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8628_ _3468_ _4189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8559_ reg_file.reg_storage\[12\]\[11\] _3951_ _4138_ _4144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output192_I net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_141_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7140__A1 net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7732__I _3542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7443__A2 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__A3 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8943__A2 _4388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6083__I _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8004__S _3775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_133_clk clknet_4_4_0_clk clknet_leaf_133_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_23_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9120__A2 _4456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7131__A1 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5368__S1 _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7434__A2 _3253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7930_ _3712_ _3560_ _3700_ _3723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_117_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7861_ _2968_ _3641_ _3642_ net43 _3662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__9187__A2 _4538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5540__S1 _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8934__A2 _4375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6812_ _2684_ _2706_ _1916_ _2707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9600_ _0386_ clknet_leaf_129_clk reg_file.reg_storage\[1\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7198__A1 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5748__A2 _1663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7792_ reg_file.reg_storage\[5\]\[13\] _3598_ _3569_ _3599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9531_ _0317_ clknet_leaf_99_clk reg_file.reg_storage\[11\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ _2067_ _2641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9462_ _0248_ clknet_leaf_88_clk reg_file.reg_storage\[12\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_102_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6674_ _2345_ _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8413_ reg_file.reg_storage\[14\]\[20\] _4049_ _4053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5625_ _1385_ _1525_ _1540_ _1541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9393_ _0179_ clknet_leaf_31_clk reg_file.reg_storage\[14\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5337__I _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8344_ _4006_ _4007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5556_ reg_file.reg_storage\[12\]\[31\] reg_file.reg_storage\[13\]\[31\] reg_file.reg_storage\[14\]\[31\]
+ reg_file.reg_storage\[15\]\[31\] _1471_ _1465_ _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7122__A1 net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8648__I _4180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9111__A2 _4488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8275_ _3954_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5359__S1 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5487_ _1353_ net18 _1402_ _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7226_ _3042_ _3068_ _3074_ net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7673__A2 _3403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I mem_ld_dat[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4731__I0 reg_file.reg_storage\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__A1 _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7157_ _1374_ _3018_ _3017_ _1679_ _2993_ net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_7088_ net4 _2972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6108_ _2021_ _2022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6039_ _1952_ _1953_ _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9178__A2 _4525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4860__B _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5295__S0 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_115_clk clknet_4_12_0_clk clknet_leaf_115_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5047__S0 _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8759__S _4265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__A3 _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7113__A1 _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9102__A2 _4481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7416__A2 net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__A1 _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6927__A1 _2038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5286__S0 _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_106_clk clknet_4_13_0_clk clknet_leaf_106_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7637__I _3454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5358__S _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5589__S1 _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6390_ _2047_ _2298_ _2299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5410_ reg_file.reg_storage\[1\]\[1\] _1326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput104 net104 mem_addr[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput115 net115 mem_addr[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5341_ reg_file.reg_storage\[3\]\[6\] _0758_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4996__I _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput126 net126 mem_addr[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput159 net159 mem_st_dat[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput148 net148 mem_st_dat[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput137 net137 mem_st_dat[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_130_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8060_ _3753_ _3808_ _3815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5272_ reg_file.reg_storage\[8\]\[11\] reg_file.reg_storage\[9\]\[11\] reg_file.reg_storage\[10\]\[11\]
+ reg_file.reg_storage\[11\]\[11\] _0779_ _1135_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7011_ _2284_ _2472_ _2898_ _2610_ _2899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5821__S _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7407__A2 _3228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8962_ reg_file.reg_storage\[9\]\[29\] _4396_ _4401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5418__A1 _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__I _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7913_ _3702_ _3323_ _3497_ _1384_ _3708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__7748__S _3492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8893_ _4359_ _4360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_104_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7844_ _3607_ _3235_ _3634_ _3646_ _3647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_93_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7775_ _3571_ _3582_ _3583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_135_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ _0902_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_93_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6726_ _2623_ _2598_ _2624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6394__A2 _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9514_ _0300_ clknet_leaf_3_clk reg_file.reg_storage\[11\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__I _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9445_ _0231_ clknet_leaf_40_clk reg_file.reg_storage\[12\]\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6657_ _2557_ net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_33_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6588_ _2215_ _2211_ _2060_ _2491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5608_ _1377_ _1408_ _1461_ _1523_ _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_9376_ _0162_ clknet_leaf_134_clk reg_file.reg_storage\[14\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8327_ reg_file.reg_storage\[7\]\[25\] _3916_ _3994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5539_ _1372_ _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4952__I0 reg_file.reg_storage\[12\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8258_ _3942_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output155_I net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8189_ _3657_ _3888_ _3894_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5016__B _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7209_ _3050_ _3059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5530__I _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5268__S0 _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6385__A2 _2290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6137__A2 _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput17 inst[24] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput28 inst[5] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput39 mem_ld_dat[15] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7885__A2 _3682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5196__I0 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5648__A1 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__A1 _1902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9011__A1 _3623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4910_ _0805_ _0816_ _0819_ _0820_ _0822_ _0825_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5890_ _1803_ _1293_ _0743_ _1805_ _1279_ _1806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_90_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4841_ _0756_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_135_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6271__I _2040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7560_ _3378_ _3379_ _3380_ _3381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4772_ _0687_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_126_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6511_ _1682_ _2401_ _2416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7491_ _3317_ _1404_ _3318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9230_ _0016_ clknet_leaf_60_clk reg_file.reg_storage\[5\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7876__A2 _3658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6442_ _2323_ _2349_ _2350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_140_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9161_ _4524_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5887__A1 _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8112_ reg_file.reg_storage\[2\]\[21\] _3842_ _3847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5615__I _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6373_ _2280_ _2281_ _2282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9092_ reg_file.reg_storage\[4\]\[14\] _4475_ _4482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5639__A1 _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5324_ _1239_ _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8043_ reg_file.reg_storage\[3\]\[28\] _3799_ _3803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5255_ reg_file.reg_storage\[12\]\[15\] reg_file.reg_storage\[13\]\[15\] reg_file.reg_storage\[14\]\[15\]
+ reg_file.reg_storage\[15\]\[15\] _0817_ _0818_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6687__I0 _2523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7830__I _3431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5186_ _1073_ _1101_ _0886_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_143_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8945_ _4230_ _4388_ _4391_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8876_ reg_file.reg_storage\[10\]\[27\] _4346_ _4349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7827_ _2982_ _3630_ _3579_ _3631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_94_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7758_ _3566_ _3567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _2177_ _2607_ _2189_ _2608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6119__A2 _2032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7689_ reg_file.reg_storage\[5\]\[6\] _3444_ _3503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_50_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5178__I0 reg_file.reg_storage\[12\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7867__A2 _3658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9428_ _0214_ clknet_leaf_28_clk reg_file.reg_storage\[13\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9359_ _0145_ clknet_leaf_55_clk reg_file.reg_storage\[7\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5725__S1 _1623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__I _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_62_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_87_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7187__I _3038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_77_clk_I clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_120_clk_I clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5435__I _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9573__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8283__A2 _3959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_135_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5040_ _0768_ reg_file.reg_storage\[3\]\[19\] _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_15_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6046__A1 _1959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6991_ _0997_ _2879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5942_ _1620_ _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8730_ _4260_ _4261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6597__A2 _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5873_ _0703_ _1788_ _0723_ _1789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8661_ reg_file.reg_storage\[8\]\[13\] _4211_ _4186_ _4212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8592_ _4119_ _4162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4824_ net17 _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_7612_ _3430_ _3431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4755_ _0670_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7543_ _3359_ _3365_ _3366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_16_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4780__A1 _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9213_ _4012_ _4507_ _4553_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4686_ _0591_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_4_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7474_ _3272_ net112 _3303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5404__S0 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7761__S _3569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6425_ _2332_ _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_112_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6356_ _2073_ _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_8_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9144_ _3918_ _4512_ _4514_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5307_ reg_file.reg_storage\[8\]\[8\] reg_file.reg_storage\[9\]\[8\] reg_file.reg_storage\[10\]\[8\]
+ reg_file.reg_storage\[11\]\[8\] _0940_ _1062_ _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_9075_ _4460_ _4472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8026_ _3675_ _3791_ _3793_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6287_ _2198_ _2194_ _0677_ _2199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6285__A1 _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5238_ _0892_ reg_file.reg_storage\[3\]\[14\] _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input31_I inst[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_95_clk clknet_4_15_0_clk clknet_leaf_95_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8026__A2 _3791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5169_ _1084_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6037__A1 _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output118_I net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4625__S _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8928_ reg_file.reg_storage\[9\]\[14\] _4375_ _4382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8859_ _4225_ _4338_ _4339_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5166__I3 _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8265__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__I0 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_86_clk clknet_4_14_0_clk clknet_leaf_86_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8017__A2 _3778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_27_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__S0 _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6200__A1 _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7190_ _3041_ _3042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6210_ _1937_ _1939_ _2122_ _2123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_36_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6141_ _2026_ _2043_ _2054_ _2055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_1_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6072_ _1335_ _1985_ _1986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_127_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9205__A1 _3999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5023_ reg_file.reg_storage\[4\]\[18\] reg_file.reg_storage\[5\]\[18\] reg_file.reg_storage\[6\]\[18\]
+ reg_file.reg_storage\[7\]\[18\] _0810_ _0842_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_leaf_77_clk clknet_4_12_0_clk clknet_leaf_77_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6019__A1 _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_45_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9100__I _4460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6974_ _2860_ _2862_ _2863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9693_ _0479_ clknet_leaf_92_clk reg_file.reg_storage\[15\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8713_ _3739_ _4248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5925_ _1814_ _1824_ _1837_ net224 _1840_ _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_118_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8644_ _3529_ _4200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5856_ _1771_ _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_119_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4807_ _0712_ _0709_ _0710_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_35_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8575_ reg_file.reg_storage\[12\]\[18\] _4152_ _4153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5787_ _1670_ _1702_ _1703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4738_ _0607_ _0597_ _0611_ _0653_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7526_ _3307_ _3318_ _3347_ _3349_ _3350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_32_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8495__A2 _4099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input79_I pc[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4669_ _0586_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7457_ net78 _1525_ _3263_ _3260_ _3287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_31_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5148__I3 reg_file.reg_storage\[7\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6408_ _2238_ _2310_ _2313_ _2314_ _2315_ _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_9127_ _4006_ _4498_ _4501_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7388_ _3213_ _3223_ _3224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__S1 _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6339_ _2245_ _2051_ _2247_ _2248_ _2249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8247__A2 _3923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9058_ _4460_ _4461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8009_ _3783_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_68_clk clknet_4_11_0_clk clknet_leaf_68_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4992__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__B2 _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5186__S _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4744__A1 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8486__A2 _4094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4773__B _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6421__A1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5710_ reg_file.reg_storage\[1\]\[17\] _1625_ _1623_ _1626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6690_ _2463_ _2331_ _2584_ _2589_ _2590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_72_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ _1429_ _1352_ _1479_ _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_142_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8360_ reg_file.reg_storage\[14\]\[0\] _4019_ _4020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5572_ _1468_ _1033_ _1485_ _1487_ _1488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4735__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8291_ _3648_ _3966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_124_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7311_ _3060_ _3151_ _3152_ _3153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_25_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7242_ _3087_ _3088_ _3089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_13_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4948__B _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7173_ _3028_ _3029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8229__A2 _3761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5550__I3 reg_file.reg_storage\[7\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6124_ _2037_ _2038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6055_ _0744_ _1935_ _1969_ _1113_ _1970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5006_ _0836_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_107_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6957_ _2189_ _2386_ _2067_ _2847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6412__A1 _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9676_ _0462_ clknet_leaf_62_clk reg_file.reg_storage\[15\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6888_ _2663_ _2779_ _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5908_ _1721_ _1822_ _1823_ _1824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_49_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ _1745_ _1754_ _1755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8627_ _4188_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8558_ _4143_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output185_I net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7509_ _1088_ _1416_ _3334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8489_ _4073_ _4099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4585__S0 _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7600__B1 _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4965__A1 _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8459__A2 _4075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5443__I _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5532__I3 reg_file.reg_storage\[7\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7860_ _3431_ _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _2106_ _2706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6945__A2 _2797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7791_ _3597_ _3598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9530_ _0316_ clknet_leaf_99_clk reg_file.reg_storage\[11\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4723__S _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6742_ _2463_ _2380_ _2635_ _2639_ _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_9_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5618__I _1533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6673_ _1580_ _2573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6223__B _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9461_ _0247_ clknet_leaf_20_clk reg_file.reg_storage\[12\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9392_ _0178_ clknet_leaf_33_clk reg_file.reg_storage\[14\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8412_ _3974_ _4051_ _4052_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5624_ _0736_ _1539_ _1540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8343_ _3739_ _4006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5555_ _1360_ _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_41_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8274_ reg_file.reg_storage\[7\]\[12\] _3953_ _3927_ _3954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5486_ _1355_ _1402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7225_ _3059_ net122 _3061_ _3073_ _3074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7156_ _1397_ _3018_ _3017_ _1828_ _2991_ net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__5684__A2 _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4731__I1 reg_file.reg_storage\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6107_ _1786_ _2021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7087_ _2970_ _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8664__I _4181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8622__A2 _4182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6038_ _0933_ _0970_ _1953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_68_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output100_I net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7989_ _3478_ _3765_ _3772_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5295__S1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9659_ _0445_ clknet_leaf_98_clk reg_file.reg_storage\[4\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8689__A2 _4226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5047__S1 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7361__A2 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6359__I _2170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5124__A1 _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8861__A2 _4338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8574__I _4126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5427__A2 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4730__S0 _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5286__S1 _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8129__A1 _3734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7352__A2 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7653__I _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__A1 _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput105 net105 mem_addr[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput116 net116 mem_addr[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_140_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5340_ reg_file.reg_storage\[1\]\[6\] _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput127 net127 mem_addr[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput138 net138 mem_st_dat[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput149 net149 mem_st_dat[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5271_ reg_file.reg_storage\[12\]\[11\] reg_file.reg_storage\[13\]\[11\] reg_file.reg_storage\[14\]\[11\]
+ reg_file.reg_storage\[15\]\[11\] _0920_ _1135_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5115__A1 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8852__A2 _4325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7010_ _2704_ _2892_ _2897_ _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_10_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8961_ _4246_ _4398_ _4400_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6615__A1 _2494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5418__A2 _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7912_ _2978_ _3535_ _3700_ _3707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_78_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8892_ _3425_ _4178_ _4359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_144_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7843_ _3228_ _3645_ _3646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4986_ _0759_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7774_ _3572_ _3167_ _3573_ _3580_ _3581_ _3582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_9513_ _0299_ clknet_leaf_52_clk reg_file.reg_storage\[11\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6725_ _2567_ _2623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_63_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7049__B _2086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5029__S1 _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6656_ _1997_ _2541_ _2556_ _2557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9444_ _0230_ clknet_leaf_16_clk reg_file.reg_storage\[12\]\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6587_ _2481_ _2489_ _2490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5607_ _1478_ _1496_ _1509_ _1522_ _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_5_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9375_ _0161_ clknet_leaf_4_clk reg_file.reg_storage\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9096__A2 _4475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8326_ _3992_ _3993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5538_ reg_file.reg_storage\[8\]\[24\] reg_file.reg_storage\[9\]\[24\] reg_file.reg_storage\[10\]\[24\]
+ reg_file.reg_storage\[11\]\[24\] _1446_ _1451_ _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_41_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input61_I mem_ld_dat[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8257_ reg_file.reg_storage\[7\]\[7\] _3940_ _3941_ _3942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5083__I _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5469_ _0671_ _1385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7208_ net87 _3058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8188_ reg_file.reg_storage\[6\]\[18\] _3893_ _3894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output148_I net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7139_ _3007_ _3000_ _3008_ net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_100_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A2 _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5268__S1 _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput18 inst[25] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_135_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5196__I1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput29 inst[6] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7098__A1 _2969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8598__A1 reg_file.reg_storage\[12\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9011__A2 _4405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4840_ _0755_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5369__S _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5584__A1 _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4771_ _0686_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6510_ _1192_ _1666_ _2414_ _2415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_126_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7490_ net82 _3317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6441_ _2296_ _2330_ _2341_ _2342_ _2348_ _2349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_3_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9160_ reg_file.reg_storage\[15\]\[8\] _3530_ _4522_ _4524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6372_ _2238_ _2242_ _2236_ _2281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5887__A2 _1763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8111_ _3675_ _3844_ _3846_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5323_ net156 _1238_ _0679_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5832__S _1642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9091_ _4461_ _4481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_61_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_143_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8042_ _3726_ _3801_ _3802_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5254_ _0807_ _1167_ _1168_ _1169_ _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5639__A2 _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6687__I1 _2586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4942__S0 _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5185_ _1087_ _1100_ _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8589__A1 _3990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9103__I _4466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6064__A2 _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8944_ reg_file.reg_storage\[9\]\[21\] _4386_ _4391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8875_ _4305_ _4348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7826_ _3481_ _3628_ _3629_ _3630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7564__A2 _3384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7757_ _2438_ _3504_ _3565_ _3566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_46_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4969_ _0884_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8513__A1 reg_file.reg_storage\[13\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7688_ _3501_ _3502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6708_ _2502_ _2606_ _2198_ _2607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5178__I1 reg_file.reg_storage\[13\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9427_ _0213_ clknet_leaf_27_clk reg_file.reg_storage\[13\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6639_ _2539_ _2540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9358_ _0144_ clknet_leaf_56_clk reg_file.reg_storage\[7\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9069__A2 _4463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9289_ _0075_ clknet_leaf_44_clk reg_file.reg_storage\[2\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8309_ _3681_ _3980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8816__A2 _4312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7252__A1 _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6055__A2 _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5802__A2 _1717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7004__A1 _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__S0 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8504__A1 _3990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5318__A1 _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4620__I _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6294__A2 _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6990_ _2878_ net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_0_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ _0969_ _1647_ _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5400__B _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8660_ _3596_ _4211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5872_ net24 _0701_ _0715_ _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8591_ _3993_ _4121_ _4161_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7611_ _3429_ _3430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4823_ _0738_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4754_ _0669_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7542_ _3344_ _3356_ _3365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7473_ _3296_ _3301_ _3302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9212_ reg_file.reg_storage\[15\]\[31\] _4505_ _4553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4685_ _0590_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5404__S1 _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6424_ _1120_ _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6355_ _2261_ _2264_ _2265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_8_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9143_ reg_file.reg_storage\[15\]\[1\] _4513_ _4514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_112_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5306_ reg_file.reg_storage\[12\]\[8\] reg_file.reg_storage\[13\]\[8\] reg_file.reg_storage\[14\]\[8\]
+ reg_file.reg_storage\[15\]\[8\] _0801_ _0983_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_59_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9074_ _3937_ _4462_ _4471_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6286_ _2109_ _2198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5237_ reg_file.reg_storage\[1\]\[14\] _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8025_ reg_file.reg_storage\[3\]\[20\] _3789_ _3793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5168_ _1074_ _1083_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input24_I inst[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5099_ reg_file.reg_storage\[4\]\[31\] reg_file.reg_storage\[5\]\[31\] reg_file.reg_storage\[6\]\[31\]
+ reg_file.reg_storage\[7\]\[31\] _0896_ _0961_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_75_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7234__A1 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8927_ _4361_ _4381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4705__I _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6192__I _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8858_ reg_file.reg_storage\[10\]\[19\] _4336_ _4339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7809_ net57 _3614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8789_ _4238_ _4256_ _4295_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_35_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5159__S0 _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6276__A2 _2187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5323__I1 _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7225__B2 _3073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8973__A1 _3911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5331__S0 _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6035__C _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__S1 _1483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__I _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6140_ _2046_ _2053_ _2054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6071_ _1182_ _1904_ _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_127_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _0631_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8492__I _4079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7216__A1 _3058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8964__A1 reg_file.reg_storage\[9\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6973_ _2861_ _2839_ _2862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9692_ _0478_ clknet_leaf_91_clk reg_file.reg_storage\[15\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8712_ _4246_ _4244_ _4247_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5924_ _1838_ _1839_ _1840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8643_ _4199_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ _1769_ _0792_ _1354_ _1770_ _1771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_36_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8192__A2 _3895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4806_ net24 _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_138_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8574_ _4126_ _4152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5786_ _0491_ _1701_ _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_133_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4737_ _0598_ _0589_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7525_ _3317_ _1404_ _3349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4668_ net27 _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__5389__S0 _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7456_ net79 _1568_ _3286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8667__I _3622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6407_ _2240_ _2235_ _2241_ _2278_ _2315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_clkbuf_leaf_61_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9126_ reg_file.reg_storage\[4\]\[29\] _4496_ _4501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7387_ _3220_ _3222_ _3223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4599_ _0523_ net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6338_ _2001_ _2248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9057_ _4459_ _4460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6269_ _2179_ _2180_ _2181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8008_ reg_file.reg_storage\[3\]\[13\] _3598_ _3768_ _3783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_76_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7207__A1 _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8183__A2 _3882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7746__I _3555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A2 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_134_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9132__A1 _3754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5941__A1 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4744__A2 _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8577__I _4132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7694__A1 _3047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6097__I _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9199__A1 _3992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5640_ _1544_ _1555_ _1556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9123__A1 _3999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5571_ _1432_ reg_file.reg_storage\[2\]\[30\] _1486_ _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8290_ _3964_ _3959_ _3965_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7310_ _3149_ _3150_ _3152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7241_ _3058_ net90 net91 _3088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5904__I _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7172_ _3027_ _3028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_55_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6123_ _2034_ _2037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7988__A2 _3766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5999__A1 _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6054_ _0744_ _1951_ _1968_ _1969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5005_ _0920_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_0_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8937__A1 reg_file.reg_storage\[9\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6956_ _2424_ _2638_ _2845_ _2846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_120_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ _1162_ _1720_ _1823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_37_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6887_ _2677_ _2700_ _2778_ _2746_ _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_48_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9675_ _0461_ clknet_leaf_9_clk reg_file.reg_storage\[15\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8626_ reg_file.reg_storage\[8\]\[2\] _4185_ _4187_ _4188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input91_I pc[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6176__A1 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5838_ _1216_ _1753_ _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8557_ reg_file.reg_storage\[12\]\[10\] _3949_ _4138_ _4143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5769_ reg_file.reg_storage\[2\]\[12\] reg_file.reg_storage\[3\]\[12\] _1357_ _1685_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7508_ _3035_ _2855_ _3200_ _3328_ _3333_ net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8488_ _3967_ _4094_ _4098_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_114_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6479__A2 _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output178_I net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7439_ _3060_ _3270_ _3271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4585__S1 _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9109_ _3980_ _4488_ _4491_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6403__A2 _2234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7600__B2 _3403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7600__A1 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8156__A2 _3870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9309__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5773__S0 _1532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7419__A1 _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6810_ _2002_ _2503_ _2705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7790_ _3596_ _3597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6741_ _2324_ _2638_ _2326_ _2639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6672_ _1112_ _2571_ _2572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9460_ _0246_ clknet_leaf_28_clk reg_file.reg_storage\[12\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9391_ _0177_ clknet_leaf_54_clk reg_file.reg_storage\[14\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8411_ reg_file.reg_storage\[14\]\[19\] _4049_ _4052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5623_ _0491_ _1538_ _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_73_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8342_ _4004_ _4001_ _4005_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5554_ _1427_ _1016_ _1467_ _1469_ _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_103_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5485_ _1400_ _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8273_ _3583_ _3953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8010__I _3764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7224_ _3067_ _3069_ _3072_ _3073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6330__A1 _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7155_ _3001_ _3018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4731__I2 reg_file.reg_storage\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6106_ _0833_ _0972_ _2011_ _2020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7086_ _2969_ _2970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4644__A1 _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__I _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6037_ _1175_ _1163_ _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xrebuffer30 _1519_ net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XTAP_TAPCELL_ROW_68_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8680__I _3666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7988_ reg_file.reg_storage\[3\]\[4\] _3766_ _3772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6939_ _2829_ net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_49_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9658_ _0444_ clknet_leaf_99_clk reg_file.reg_storage\[4\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8609_ _4172_ _4173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9589_ _0375_ clknet_leaf_119_clk reg_file.reg_storage\[9\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5124__A2 _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4883__A1 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6308__C _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4730__S1 _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8377__A2 _4025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_72_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_28_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5060__A1 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5655__S _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9281__CLK clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5363__A2 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput106 net106 mem_addr[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_106_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput139 net139 mem_st_dat[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput128 net128 mem_addr[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput117 net117 mem_addr[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5270_ reg_file.reg_storage\[1\]\[11\] _1185_ _1135_ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_81_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5115__A2 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5746__S0 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4874__A1 _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8960_ reg_file.reg_storage\[9\]\[28\] _4396_ _4400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7911_ _3400_ _3705_ _3706_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_90_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8891_ _4170_ _4356_ _4358_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8368__A2 _4026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7842_ _3438_ _3645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4985_ _0765_ _0895_ _0898_ _0900_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5051__A1 _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7773_ _1692_ _3464_ _3466_ _3581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9512_ _0298_ clknet_leaf_53_clk reg_file.reg_storage\[11\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6724_ _2599_ _2621_ _2622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_73_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9443_ _0229_ clknet_leaf_136_clk reg_file.reg_storage\[12\]\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6655_ _2056_ _2545_ _2550_ _2192_ _2555_ _2556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_61_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9374_ _0160_ clknet_leaf_87_clk reg_file.reg_storage\[14\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7894__A4 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _2482_ _2488_ _2489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5606_ _0995_ _1521_ _1522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer27_I _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5537_ reg_file.reg_storage\[12\]\[24\] reg_file.reg_storage\[13\]\[24\] reg_file.reg_storage\[14\]\[24\]
+ reg_file.reg_storage\[15\]\[24\] _1428_ _1451_ _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_103_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8325_ _3709_ _3992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5364__I _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8256_ _3921_ _3941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_42_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input54_I mem_ld_dat[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7207_ _1324_ _3042_ _3057_ net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5468_ _1381_ _1382_ _1383_ _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8187_ _3867_ _3893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5399_ reg_file.reg_storage\[3\]\[3\] _0999_ _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7138_ net156 _3004_ _3008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7069_ _2194_ _1921_ _2108_ _2954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_129_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6128__C _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_138_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5475__S _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 inst[26] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5274__I _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7098__A2 _2972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__S0 _1532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5223__B _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__A1 _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8770__A2 _4275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5033__A1 _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ _0685_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_7_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6533__A1 _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6440_ _2343_ _1827_ _2344_ _2347_ _2348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_43_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6371_ _1938_ _2234_ _2280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7089__A2 _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8110_ reg_file.reg_storage\[2\]\[20\] _3842_ _3846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5322_ _1235_ _1237_ _0738_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9090_ _4480_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8041_ reg_file.reg_storage\[3\]\[27\] _3799_ _3802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5253_ _0813_ reg_file.reg_storage\[2\]\[15\] _0814_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5184_ _1099_ _0875_ _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_110_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4942__S1 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8943_ _4228_ _4388_ _4390_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8874_ _4240_ _4306_ _4347_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7825_ net48 _3404_ _3406_ _3629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8210__A1 _3726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7756_ _3161_ _3402_ _3546_ _3563_ _3564_ _3565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4968_ net226 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4899_ _0813_ reg_file.reg_storage\[2\]\[21\] _0814_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7687_ net125 _3432_ _3495_ _3500_ _3501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_6707_ _2194_ _2604_ _2605_ _2606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5178__I2 reg_file.reg_storage\[14\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9426_ _0212_ clknet_leaf_71_clk reg_file.reg_storage\[13\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6638_ _1731_ _2538_ _2539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_50_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9357_ _0143_ clknet_leaf_12_clk reg_file.reg_storage\[7\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8308_ _3978_ _3975_ _3979_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_76_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6569_ _2193_ _2472_ _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9288_ _0074_ clknet_leaf_45_clk reg_file.reg_storage\[2\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output160_I net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8239_ reg_file.reg_storage\[7\]\[2\] _3926_ _3928_ _3929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5043__B _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7788__B1 _3573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5110__S1 _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7960__B1 _3496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4613__I1 reg_file.reg_storage\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4901__I _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5318__A2 _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4621__S0 _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6818__A2 _1542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6294__A3 _2204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7491__A2 _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5254__A1 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ _1556_ _1855_ _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8991__A2 _4411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7610_ _0600_ _0661_ _0665_ _3429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5871_ _1766_ _1787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8590_ reg_file.reg_storage\[12\]\[25\] _4122_ _4161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4822_ _0592_ _0662_ _0654_ _0656_ _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_29_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4753_ _0668_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_50_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7541_ _3359_ _3360_ _3363_ _3364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_28_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6506__A1 _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7472_ _3286_ _3298_ _3300_ _3301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4811__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9211_ _4009_ _4548_ _4552_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6423_ _2245_ _1797_ _2331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4684_ net29 _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_141_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9142_ _4509_ _4513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6354_ _2071_ _2263_ _2022_ _2264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_112_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5305_ reg_file.reg_storage\[1\]\[8\] _1220_ _1062_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9073_ reg_file.reg_storage\[4\]\[6\] _4463_ _4471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6285_ _2194_ _2195_ _2196_ _2197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5236_ reg_file.reg_storage\[4\]\[14\] reg_file.reg_storage\[5\]\[14\] reg_file.reg_storage\[6\]\[14\]
+ reg_file.reg_storage\[7\]\[14\] _1021_ _1022_ _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_8024_ _3667_ _3791_ _3792_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_71_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5167_ _0754_ _1082_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7569__I net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5245__A1 _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5098_ _0753_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input17_I inst[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8926_ _4380_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8857_ _4316_ _4338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8734__A2 _4262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8788_ reg_file.reg_storage\[11\]\[25\] _4257_ _4295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7808_ net103 _3472_ _3613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_35_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7739_ _3447_ _3481_ _3517_ _3549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9409_ _0195_ clknet_leaf_132_clk reg_file.reg_storage\[13\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5720__A2 _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5159__S1 _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_89_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8422__A1 _3990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7225__A2 net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8973__A2 _4406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5331__S1 _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5787__A2 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7161__A1 net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7161__B2 _1690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7942__I _3733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5462__I _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6070_ _1983_ _1984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input9_I inst[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_127_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ _0621_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_140_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4806__I net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8711_ reg_file.reg_storage\[8\]\[28\] _4241_ _4247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_109_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6972_ _2841_ _2837_ _2861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9691_ _0477_ clknet_leaf_96_clk reg_file.reg_storage\[15\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5923_ _1731_ _1839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8642_ reg_file.reg_storage\[8\]\[7\] _4197_ _4198_ _4199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6727__B2 _2560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5854_ _0690_ _0584_ _0691_ _0692_ _1770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_8573_ _3967_ _4147_ _4151_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4805_ _0713_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5785_ _1696_ _1698_ _1699_ _1700_ _1533_ _1536_ _1701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_17_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7524_ _3309_ _3319_ _3347_ _3348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_29_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4736_ _0609_ _0604_ _0612_ _0607_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__7152__A1 _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4667_ _0585_ net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7455_ _3284_ _3274_ _3285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_142_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7386_ _3173_ _3175_ _3221_ _3168_ _3222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6406_ _1810_ _2277_ _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_9125_ _4003_ _4498_ _4500_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6337_ _2246_ _2032_ _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4598_ _0487_ _0522_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_101_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__S0 _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9056_ _3424_ _4124_ _4459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6268_ _2041_ _1045_ _2180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5219_ _0635_ _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8007_ _3782_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6199_ _2110_ _2111_ _2112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output123_I net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4716__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8909_ reg_file.reg_storage\[9\]\[6\] _4363_ _4371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__S0 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5547__I _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9132__A2 _4015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7694__A2 _3115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8946__A2 _4361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7937__I _3547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_136_clk clknet_4_4_0_clk clknet_leaf_136_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5570_ _1426_ _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4735__A3 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7134__A1 net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9123__A2 _4498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7240_ net92 _3087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7171_ _3026_ _3027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6122_ _2035_ _2036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6053_ _1111_ _1967_ _1968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5004_ _0919_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8937__A2 _4386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6948__A1 _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _2005_ _2843_ _2844_ _2214_ _2845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_49_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_138_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_120_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5906_ _1816_ _1819_ _1821_ _1822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9674_ _0460_ clknet_leaf_8_clk reg_file.reg_storage\[15\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_127_clk clknet_4_5_0_clk clknet_leaf_127_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6886_ _2723_ _2778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8625_ _4186_ _4187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_36_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5837_ _1497_ _0736_ _1402_ net213 _1753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_101_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8556_ _3946_ _4128_ _4142_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5768_ reg_file.reg_storage\[8\]\[12\] reg_file.reg_storage\[9\]\[12\] reg_file.reg_storage\[10\]\[12\]
+ reg_file.reg_storage\[11\]\[12\] _1606_ _1608_ _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_133_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7125__A1 _1717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8487_ reg_file.reg_storage\[13\]\[17\] _4088_ _4098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9114__A2 _4457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4719_ _0634_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input84_I pc[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7507_ _3330_ _3331_ _3332_ _3333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_32_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5699_ _1614_ _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_60_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7438_ _3265_ _3268_ _3264_ _3270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_102_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7369_ _1165_ _3205_ _3206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9108_ reg_file.reg_storage\[4\]\[21\] _4486_ _4491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9039_ reg_file.reg_storage\[1\]\[27\] _4443_ _4448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_110_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8928__A2 _4375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9050__A1 _3388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6661__I _2560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_118_clk clknet_4_1_0_clk clknet_leaf_118_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_15_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7116__A1 _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9105__A2 _4488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5773__S1 _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_109_clk clknet_4_13_0_clk clknet_leaf_109_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6740_ _2524_ _2637_ _2101_ _2638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_60_clk_I clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6671_ _2570_ _2571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6158__A2 _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7355__A1 _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5187__I _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9390_ _0176_ clknet_leaf_56_clk reg_file.reg_storage\[14\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5622_ _1526_ _1528_ _1529_ _1530_ _1534_ _1537_ _1538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_8410_ _4029_ _4051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_61_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8341_ reg_file.reg_storage\[7\]\[28\] _3997_ _4005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5553_ _1432_ reg_file.reg_storage\[2\]\[31\] _1468_ _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_75_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8272_ _3952_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5484_ _1378_ _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5669__A1 _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5213__S0 _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7658__A2 _3080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7223_ _3070_ _3063_ _3071_ _3072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7154_ _1457_ _3012_ _3017_ net212 _2990_ net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__8607__A1 _3760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4731__I3 reg_file.reg_storage\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6105_ _0877_ _1073_ _2018_ _2019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_133_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7085_ _0727_ _2969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_13_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7778__S _3569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6036_ _1786_ _1943_ _1950_ _1119_ _1951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xrebuffer20 _1506_ net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4644__A2 net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5841__A1 _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer31 _2886_ net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XTAP_TAPCELL_ROW_68_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_28_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6481__I _1959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7987_ _3771_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6938_ _2813_ _2815_ _2824_ _2828_ _2829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_64_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9657_ _0443_ clknet_leaf_102_clk reg_file.reg_storage\[4\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6869_ _2742_ _1844_ _2345_ _2761_ _2762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_76_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8608_ _4118_ _4171_ _4172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9588_ _0374_ clknet_leaf_117_clk reg_file.reg_storage\[9\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7897__A2 _3294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8539_ reg_file.reg_storage\[12\]\[2\] _3926_ _4132_ _4133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_output190_I net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8074__A2 _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6605__B _2507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6560__A2 _2187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput107 net107 mem_addr[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_50_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput118 net118 mem_addr[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput129 net129 mem_ld_en vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_121_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5746__S1 _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4874__A2 _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8065__A2 _3819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8982__S _4415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8890_ reg_file.reg_storage\[9\]\[0\] _4357_ _4358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7910_ reg_file.reg_storage\[5\]\[24\] _3422_ _3706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7841_ _3640_ _3643_ _3539_ _3644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7772_ _3537_ _3578_ _3579_ _3580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4984_ _0773_ reg_file.reg_storage\[2\]\[17\] _0899_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9511_ _0297_ clknet_leaf_27_clk reg_file.reg_storage\[11\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6723_ _2593_ _2595_ _2621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_58_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5051__A2 _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6654_ _2551_ _1839_ _2552_ _2554_ _2555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_63_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9442_ _0228_ clknet_leaf_131_clk reg_file.reg_storage\[12\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5605_ _1417_ _1511_ _1520_ _1521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__6000__A1 _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9373_ _0159_ clknet_leaf_91_clk reg_file.reg_storage\[7\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6585_ _2483_ _2487_ _2488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8324_ _3990_ _3915_ _3991_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5536_ reg_file.reg_storage\[1\]\[24\] _1449_ _1451_ _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8255_ _3509_ _3940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5467_ _1355_ _1383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7860__I _3431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7206_ _3051_ _1982_ _3053_ _3056_ _3057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input47_I mem_ld_dat[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8186_ _3649_ _3888_ _3892_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5398_ reg_file.reg_storage\[1\]\[3\] _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7137_ _3006_ net222 _3007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7068_ _1873_ _2951_ _2952_ _2953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7803__A2 _3194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4925__S _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5814__A1 _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6019_ _0980_ _1926_ _1933_ _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_69_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5673__S0 _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9599__CLK clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5555__I _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__S1 _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7645__I2 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4634__I _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6230__A1 _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_clk clknet_4_2_0_clk clknet_leaf_40_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_71_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4792__B2 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5416__S0 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5465__I _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6370_ _2278_ _2279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7730__B2 _1829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7089__A3 _2972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5321_ _1236_ _0618_ _0616_ _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8040_ _3756_ _3801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_121_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ _0811_ reg_file.reg_storage\[3\]\[15\] _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8038__A2 _3799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5183_ _1098_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_143_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8942_ reg_file.reg_storage\[9\]\[20\] _4386_ _4390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8873_ reg_file.reg_storage\[10\]\[26\] _4346_ _4347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7824_ net39 _3023_ _3627_ _3628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7013__A3 _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7855__I _3656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7755_ _3484_ _3156_ _3430_ _3564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_22_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4967_ net145 _0882_ _0679_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_31_clk clknet_4_9_0_clk clknet_leaf_31_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4898_ _0763_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_46_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6706_ _2049_ _2546_ _2605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7686_ _3048_ _3099_ _3497_ _3498_ _3499_ _3500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_117_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9425_ _0211_ clknet_leaf_30_clk reg_file.reg_storage\[13\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6637_ _1720_ _2511_ _2537_ _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_62_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9356_ _0142_ clknet_leaf_55_clk reg_file.reg_storage\[7\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6568_ _2017_ _2200_ _2471_ _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_6_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5519_ reg_file.reg_storage\[12\]\[27\] reg_file.reg_storage\[13\]\[27\] reg_file.reg_storage\[14\]\[27\]
+ reg_file.reg_storage\[15\]\[27\] _1419_ _1423_ _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_104_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8307_ reg_file.reg_storage\[7\]\[20\] _3971_ _3979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_76_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4630__S1 _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9287_ _0073_ clknet_4_3_0_clk reg_file.reg_storage\[2\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6499_ _2397_ _2402_ _2405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6288__A1 _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8238_ _3927_ _3928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_output153_I net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_98_clk clknet_4_15_0_clk clknet_leaf_98_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4719__I _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8029__A2 _3764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8169_ _3543_ _3869_ _3883_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6835__I0 _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7788__B2 _3593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6460__A1 _2110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5646__S0 _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6212__A1 _2117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6763__A2 _2659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7960__B2 _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_22_clk clknet_4_1_0_clk clknet_leaf_22_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7712__A1 _3506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_89_clk clknet_4_14_0_clk clknet_leaf_89_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_18_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5870_ _1103_ _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4821_ net3 _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_34_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7675__I _3489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_13_clk clknet_4_0_0_clk clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_60_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7540_ _3361_ _3354_ _3362_ _3363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4752_ _0666_ _0667_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_141_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4683_ _0599_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7471_ _3284_ _3299_ _3300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5195__I _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9210_ reg_file.reg_storage\[15\]\[30\] _4505_ _4552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6422_ _2325_ _2327_ _2329_ _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9141_ _4511_ _4512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6353_ _2028_ _2195_ _2262_ _2263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_112_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5304_ reg_file.reg_storage\[2\]\[8\] reg_file.reg_storage\[3\]\[8\] _0919_ _1220_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9072_ _4470_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6284_ _2049_ _1311_ _1337_ _2196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6020__S _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9294__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8023_ reg_file.reg_storage\[3\]\[19\] _3789_ _3792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5235_ net70 _0852_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6690__A1 _2463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5166_ _1075_ _1079_ _1080_ _1081_ _0965_ _0929_ _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ net89 _0750_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6442__A1 _2323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8925_ reg_file.reg_storage\[9\]\[13\] _4211_ _4365_ _4380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8856_ _4222_ _4331_ _4337_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7807_ _3600_ _3611_ _3612_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8787_ _4236_ _4256_ _4294_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5999_ _1057_ _0970_ _1914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7738_ net34 net42 _3027_ _3548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_81_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8498__A2 _4101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9408_ _0194_ clknet_leaf_134_clk reg_file.reg_storage\[13\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7669_ _0613_ _3484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5800__S0 _1533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9339_ _0125_ clknet_leaf_94_clk reg_file.reg_storage\[6\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5181__A1 _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6681__A1 _2573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6664__I _2153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6984__A2 _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6105__S _2018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6672__A1 _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5020_ net74 _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_127_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_2_clk clknet_4_4_0_clk clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8413__A2 _4049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7621__B1 _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8710_ _3733_ _4246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_109_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6971_ _1099_ _2859_ _2860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9690_ _0476_ clknet_leaf_96_clk reg_file.reg_storage\[15\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _1175_ _1838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7924__A1 net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8641_ _4180_ _4198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5853_ net20 _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8572_ reg_file.reg_storage\[12\]\[17\] _4141_ _4151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7924__B2 _3714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5784_ reg_file.reg_storage\[4\]\[13\] reg_file.reg_storage\[5\]\[13\] reg_file.reg_storage\[6\]\[13\]
+ reg_file.reg_storage\[7\]\[13\] _0687_ _1695_ _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_8_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4804_ _0704_ _0719_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_90_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4735_ _0620_ _0631_ _0650_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_8_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7523_ _3331_ _3337_ _3347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_138_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4666_ _0493_ _0584_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_44_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7454_ net79 _3284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_141_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5163__A1 _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7385_ _3185_ _3186_ _3215_ _3221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6405_ _2311_ _2312_ _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4597_ _0515_ _0517_ _0519_ _0520_ _0521_ _0485_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_9124_ reg_file.reg_storage\[4\]\[28\] _4496_ _4500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6336_ _2120_ _2246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8101__A1 _3638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9055_ _3911_ _4456_ _4458_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6267_ _2044_ _2179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5010__S1 _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5710__I0 reg_file.reg_storage\[1\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8006_ reg_file.reg_storage\[3\]\[12\] _3585_ _3768_ _3782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6198_ _1931_ _1923_ _2097_ _2111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5218_ net69 _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__8404__A2 _4044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ reg_file.reg_storage\[2\]\[25\] reg_file.reg_storage\[3\]\[25\] _0920_ _1065_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6415__A1 _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output116_I net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8908_ _4370_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8839_ reg_file.reg_storage\[10\]\[11\] _4207_ _4322_ _4328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5077__S1 _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4732__I _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4907__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6957__A2 _2386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6709__A2 _2607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4642__I _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7170_ _3025_ _3026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6121_ _2034_ _2035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_55_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6645__A1 _1955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6052_ _1958_ _1966_ _1103_ _1967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7621__C _3417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5003_ _0755_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7070__A1 _2036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6954_ _2010_ _2729_ _2844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9673_ _0459_ clknet_leaf_50_clk reg_file.reg_storage\[15\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5905_ _1820_ _1815_ _1821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6885_ _2774_ _2775_ _2776_ _2777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8624_ _4179_ _4186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_118_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5836_ _1622_ _0715_ _0692_ _1751_ _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__7373__A2 net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8555_ reg_file.reg_storage\[12\]\[9\] _4141_ _4142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5767_ _1669_ _1682_ _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8486_ _3964_ _4094_ _4097_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5698_ _0577_ _1614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_72_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7506_ _3330_ _3331_ _3044_ _3332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4718_ net8 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4649_ reg_file.reg_storage\[2\]\[6\] reg_file.reg_storage\[3\]\[6\] _0534_ _0569_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input77_I pc[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7437_ _3264_ _3265_ _3268_ _3269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_32_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8873__A2 _4346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5383__I _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7368_ _1722_ _3205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9107_ _3977_ _4488_ _4490_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7299_ _3137_ _3141_ _3142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6319_ net19 _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9038_ _3995_ _4445_ _4447_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__S _1672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9050__A2 _4118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7061__A1 _2046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5375__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8864__A2 _4311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6627__A1 _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_106_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6670_ _2251_ _2258_ _2570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_45_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5621_ _1536_ _1537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_42_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7683__I _3496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8340_ _4003_ _4004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5552_ _1426_ _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8271_ reg_file.reg_storage\[7\]\[11\] _3951_ _3941_ _3952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5118__A1 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8855__A2 _4336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5508__I3 reg_file.reg_storage\[7\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6866__A1 _2742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5483_ _1379_ _1384_ _1398_ _1071_ _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__5213__S1 _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7222_ _3066_ _0977_ _3071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7153_ _2973_ _3017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8607__A2 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5931__I _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7084_ _2967_ _2968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6618__A1 _2135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6104_ _1971_ _2018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6248__B _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6035_ _1269_ _1945_ _1949_ _0980_ _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_68_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer21 _1733_ net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer10 _1752_ net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5841__A2 _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer32 _0739_ net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XTAP_TAPCELL_ROW_81_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7986_ reg_file.reg_storage\[3\]\[3\] _3470_ _3769_ _3771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6937_ _1934_ _2796_ _2827_ _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9656_ _0442_ clknet_leaf_104_clk reg_file.reg_storage\[4\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6868_ _2759_ _2576_ _2760_ _2761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7346__A2 _3184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9587_ _0373_ clknet_leaf_77_clk reg_file.reg_storage\[9\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8607_ _3760_ _1106_ _4171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_9_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5819_ net21 _1411_ _0669_ _1735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_119_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6799_ _2583_ _2694_ _2695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8538_ _4131_ _4132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__9099__A2 _4481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output183_I net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8846__A2 _4325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8469_ _4073_ _4088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_79_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9023__A2 _4435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4920__I _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput108 net108 mem_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput119 net119 mem_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_121_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6848__A1 _1852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9014__A2 _4430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7840_ _2968_ _3641_ _3642_ net41 _3643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_78_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7771_ _3514_ _3579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_4983_ _0774_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5198__I _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9510_ _0296_ clknet_leaf_45_clk reg_file.reg_storage\[11\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6722_ _2616_ _1858_ _2574_ _2619_ _2620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__7328__A2 _1692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6653_ _2073_ _2553_ _2554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_63_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9441_ _0227_ clknet_leaf_133_clk reg_file.reg_storage\[12\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8302__I _3928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6531__B _2435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ _1351_ _1519_ _1520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6000__A2 _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9372_ _0158_ clknet_leaf_90_clk reg_file.reg_storage\[7\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6584_ _2484_ _2486_ _2487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8323_ reg_file.reg_storage\[7\]\[24\] _3916_ _3991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5535_ _1450_ _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8828__A2 _4312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6839__A1 _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8254_ _3938_ _3923_ _3939_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5466_ net18 _1382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7205_ _3054_ _3055_ _3056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8185_ reg_file.reg_storage\[6\]\[17\] _3882_ _3892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5397_ reg_file.reg_storage\[4\]\[3\] reg_file.reg_storage\[5\]\[3\] reg_file.reg_storage\[6\]\[3\]
+ reg_file.reg_storage\[7\]\[3\] _0866_ _0867_ _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7136_ _0494_ _3006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7067_ _1495_ _2928_ _2537_ _2952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5814__A2 _1729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6018_ _0980_ _1932_ _1933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6492__I _2157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_6_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5122__S0 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7969_ _3756_ _3757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5578__A1 _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5673__S1 _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9639_ _0425_ clknet_leaf_30_clk reg_file.reg_storage\[4\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5750__A1 _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7699__S _3492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6302__I0 _2211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7645__I3 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_74_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7007__A1 _2117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5361__S0 _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5569__A1 _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_89_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6230__A2 _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9180__A1 reg_file.reg_storage\[15\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_132_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4650__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5416__S1 _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_12_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__A2 _3136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer1 _1509_ net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5320_ net32 _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XTAP_TAPCELL_ROW_114_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5251_ reg_file.reg_storage\[1\]\[15\] _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_27_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4927__S0 _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8993__S _4421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5182_ _1088_ _0913_ _1097_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6049__A2 _1963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8941_ _4225_ _4388_ _4389_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_143_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8872_ _4304_ _4346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7201__I _3038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7549__A2 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7823_ _3614_ _3022_ _3627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7754_ _3514_ _3562_ _3563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6705_ _2573_ _2107_ _2603_ _2604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_46_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4966_ _0879_ _0881_ _0739_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7685_ _3486_ _3499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4897_ _0771_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_34_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9424_ _0210_ clknet_leaf_33_clk reg_file.reg_storage\[13\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6636_ _2398_ _2537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_50_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6567_ _2288_ _2470_ _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6688__S _2120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9355_ _0141_ clknet_leaf_9_clk reg_file.reg_storage\[7\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5518_ _1427_ _1090_ _1430_ _1433_ _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8306_ _3977_ _3978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_76_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9286_ _0072_ clknet_leaf_41_clk reg_file.reg_storage\[2\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6498_ _2086_ _2404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5449_ reg_file.reg_storage\[4\]\[26\] reg_file.reg_storage\[5\]\[26\] reg_file.reg_storage\[6\]\[26\]
+ reg_file.reg_storage\[7\]\[26\] _1360_ _1364_ _1365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8237_ _3920_ _3927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8168_ reg_file.reg_storage\[6\]\[9\] _3882_ _3883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output146_I net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7119_ _2988_ _2995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8099_ _3839_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7788__A2 _3182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6436__B _2171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7960__A2 _3384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5566__I _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4613__I3 reg_file.reg_storage\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5574__I1 reg_file.reg_storage\[13\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7781__I net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7476__A1 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_69_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4645__I _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8728__A1 _3761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7956__I _3745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4820_ _0735_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__9149__S _4516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7951__A2 _3740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_78_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_60_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8988__S _4415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4751_ _0599_ _0593_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_28_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4682_ _0598_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7470_ _1437_ _3138_ _1414_ _3299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_28_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6421_ _1104_ _2328_ _2329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9140_ _4510_ _4511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6352_ _2104_ _1283_ _1266_ _2262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_110_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5303_ reg_file.reg_storage\[4\]\[8\] reg_file.reg_storage\[5\]\[8\] reg_file.reg_storage\[6\]\[8\]
+ reg_file.reg_storage\[7\]\[8\] _0940_ _1062_ _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_11_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9071_ reg_file.reg_storage\[4\]\[5\] _3490_ _4466_ _4470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6283_ _1296_ _1322_ _2195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8022_ _3769_ _3791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_58_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5234_ _1133_ _1149_ _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5165_ reg_file.reg_storage\[8\]\[26\] reg_file.reg_storage\[9\]\[26\] reg_file.reg_storage\[10\]\[26\]
+ reg_file.reg_storage\[11\]\[26\] _0990_ _0922_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XPHY_EDGE_ROW_87_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_71_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5096_ _0997_ _0851_ _1011_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8924_ _4379_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8855_ reg_file.reg_storage\[10\]\[18\] _4336_ _4337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7806_ reg_file.reg_storage\[5\]\[14\] _3544_ _3612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7866__I _3666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8195__A2 _3893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_96_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8786_ reg_file.reg_storage\[11\]\[24\] _4257_ _4294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5998_ _0973_ _1908_ _1909_ _1912_ _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_35_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7737_ _3546_ _3547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4949_ _0775_ _0859_ _0862_ _0864_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7668_ _3414_ _3482_ _3483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_90_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5705__A1 _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6619_ _2248_ _2253_ _2026_ _2521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9407_ _0193_ clknet_leaf_4_clk reg_file.reg_storage\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7599_ _3409_ _3415_ _3418_ _3419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_105_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5800__S1 _1536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9338_ _0124_ clknet_leaf_95_clk reg_file.reg_storage\[6\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5181__A2 _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9269_ _0055_ clknet_leaf_23_clk reg_file.reg_storage\[3\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6681__A2 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8186__A2 _3888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7776__I _3583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8110__A2 _3842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_127_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5307__S0 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6970_ _2856_ _2858_ _2859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7621__A1 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5921_ _1826_ _1834_ _1836_ _1837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_88_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8640_ _3509_ _4197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5852_ _1293_ _1766_ _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8571_ _3964_ _4147_ _4150_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5935__A1 _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5783_ reg_file.reg_storage\[12\]\[13\] reg_file.reg_storage\[13\]\[13\] reg_file.reg_storage\[14\]\[13\]
+ reg_file.reg_storage\[15\]\[13\] _0687_ _1695_ _1699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4803_ _0713_ _0718_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4734_ _0636_ _0643_ _0646_ _0647_ _0648_ _0649_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_56_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7522_ _1511_ _3346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4665_ _0579_ _0581_ _0582_ _0583_ _0542_ _0563_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_7453_ _3144_ _3277_ _3282_ _3283_ net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_141_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8310__I _3980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7384_ _3203_ _3214_ _3218_ _3219_ _3220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_3_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6404_ _1810_ _2277_ _2312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4596_ net16 _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__4597__S1 _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9123_ _3999_ _4498_ _4499_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6335_ _2183_ _2245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9054_ reg_file.reg_storage\[4\]\[0\] _4457_ _4458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8005_ _3781_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6266_ _0887_ _1102_ _2063_ _2178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9141__I _4511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5217_ _1132_ _1042_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6197_ _2109_ _2110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5148_ reg_file.reg_storage\[4\]\[25\] reg_file.reg_storage\[5\]\[25\] reg_file.reg_storage\[6\]\[25\]
+ reg_file.reg_storage\[7\]\[25\] _1061_ _1063_ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_input22_I inst[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5079_ _0982_ _0994_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8907_ reg_file.reg_storage\[9\]\[5\] _4193_ _4366_ _4370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8168__A2 _3882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output109_I net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8838_ _4327_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8769_ _4218_ _4281_ _4284_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5777__I1 _1692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9117__A1 _3992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7143__A3 _3010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8220__I _3911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5785__S0 _1533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5537__S0 _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7603__A1 reg_file.reg_storage\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6406__A2 _2277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5480__I3 _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4923__I _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6590__A1 _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5393__A2 _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5754__I _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6120_ _1971_ _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7693__I1 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4656__A1 _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6645__A2 _2335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6051_ _0973_ _1961_ _1965_ _1966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5002_ _0893_ reg_file.reg_storage\[1\]\[16\] _0917_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_37_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5700__S0 _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6953_ _2788_ _2842_ _2105_ _2843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9672_ _0458_ clknet_leaf_49_clk reg_file.reg_storage\[15\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6884_ _1838_ _2540_ _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5904_ _1147_ _1820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5835_ _1746_ _1748_ _1749_ _1750_ _1532_ _1535_ _1751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_66_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8623_ _3454_ _4185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8570__A2 _4141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8554_ _4126_ _4141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5766_ _1681_ _1682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8485_ reg_file.reg_storage\[13\]\[16\] _4088_ _4097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5697_ reg_file.reg_storage\[1\]\[18\] _1612_ _1609_ _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4717_ _0632_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5664__I _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7505_ _3326_ _1356_ _3331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_60_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4648_ reg_file.reg_storage\[8\]\[6\] reg_file.reg_storage\[9\]\[6\] reg_file.reg_storage\[10\]\[6\]
+ reg_file.reg_storage\[11\]\[6\] _0566_ _0567_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_4_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7436_ _3256_ _3266_ _3267_ _3268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9106_ reg_file.reg_storage\[4\]\[20\] _4486_ _4490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4579_ reg_file.reg_storage\[1\]\[0\] _0504_ _0500_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7367_ _3196_ _3197_ _3203_ _3204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5519__S0 _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6318_ _2228_ net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7298_ _3139_ _3140_ _3141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7833__B2 _3636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7833__A1 net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9037_ reg_file.reg_storage\[1\]\[26\] _4443_ _4447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6249_ _2160_ _2161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8389__A2 _4025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_24_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5072__A1 _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4743__I _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4899__B _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5375__A2 _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7990__S _3769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6324__A1 _2231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_33_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6627__A2 _2510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7052__A2 _2304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_106_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5620_ _1535_ _1536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6563__A1 _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5551_ _1429_ reg_file.reg_storage\[3\]\[31\] _1467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8270_ _3566_ _3951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8304__A2 _3975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6315__A1 _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5482_ _1386_ _1397_ _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7221_ _3066_ _0977_ _3070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_117_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7152_ _1552_ _3012_ _3016_ net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7083_ _1709_ _2967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6618__A2 _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6103_ _2016_ _2017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4828__I _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6034_ _1269_ _1946_ _1948_ _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4629__A1 _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer11 _2934_ net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer22 _1631_ net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_68_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer33 _1496_ net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_49_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7985_ _3770_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6936_ _2826_ _2827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_81_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4801__A1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9655_ _0441_ clknet_leaf_115_clk reg_file.reg_storage\[4\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6867_ _2759_ _2269_ _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9067__S _4466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8543__A2 _4129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9586_ _0372_ clknet_leaf_67_clk reg_file.reg_storage\[9\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8606_ _3420_ _4170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6798_ _2176_ _2140_ _2200_ _2689_ _2693_ _2694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_8_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5818_ _1227_ _1734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_91_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8537_ _4125_ _4131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5749_ _0670_ _1664_ _1665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5394__I _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4660__S0 _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8468_ _4087_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_79_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8399_ reg_file.reg_storage\[14\]\[14\] _4038_ _4045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6857__A2 _2549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output176_I net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7419_ _0952_ _3251_ _3252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_130_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8059__A1 _3421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6609__A2 _2486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8782__A2 _4261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A2 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput109 net109 mem_addr[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_130_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__B _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5284__A1 _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8773__A2 _4286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5479__I _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7770_ _3574_ _3405_ _3407_ _3577_ _3578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4982_ _0897_ reg_file.reg_storage\[3\]\[17\] _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6784__A1 _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6721_ _2617_ _2577_ _2618_ _2619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6652_ _2551_ _1839_ _2167_ _2553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_63_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9440_ _0226_ clknet_leaf_134_clk reg_file.reg_storage\[12\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9371_ _0157_ clknet_leaf_98_clk reg_file.reg_storage\[7\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5603_ _1445_ _1518_ _1519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_73_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8322_ _3989_ _3990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_119_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6583_ _1666_ _2485_ _1681_ net209 _2486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5534_ _1421_ _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6839__A2 _2265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8253_ reg_file.reg_storage\[7\]\[6\] _3924_ _3939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ _1380_ _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8184_ _3638_ _3888_ _3891_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7204_ _1324_ _1180_ _3055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7135_ net225 _3000_ _3005_ net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_111_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5396_ net90 _0798_ _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7066_ _2926_ _2929_ _2930_ _2934_ _2951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5275__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ _1928_ _1931_ _1178_ _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8764__A2 _4275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5122__S1 _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7968_ _3755_ _3756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5578__A2 _1493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6919_ _1878_ _2809_ _2810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7899_ _3695_ _3696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_25_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9638_ _0424_ clknet_leaf_43_clk reg_file.reg_storage\[4\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6441__C _2348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9569_ _0355_ clknet_4_5_0_clk reg_file.reg_storage\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_107_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6302__I1 _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A1 _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8204__A1 _3710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5361__S1 _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_116_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5018__A1 _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9004__I0 reg_file.reg_storage\[1\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9180__A2 _4525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7715__B1 _3496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__S0 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7191__A1 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_125_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer2 _1509_ net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__S _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5250_ reg_file.reg_storage\[4\]\[15\] reg_file.reg_storage\[5\]\[15\] reg_file.reg_storage\[6\]\[15\]
+ reg_file.reg_storage\[7\]\[15\] _0802_ _0804_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_121_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4927__S1 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5181_ _1014_ _1096_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8443__A1 reg_file.reg_storage\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8940_ reg_file.reg_storage\[9\]\[19\] _4386_ _4389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6593__I _2170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8871_ _4238_ _4306_ _4345_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8746__A2 _4262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7822_ _3010_ _3408_ _3626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7753_ _3461_ _3559_ _3561_ _3522_ _3562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_93_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4965_ _0880_ _0618_ _0616_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4841__I _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6704_ _0908_ _2363_ _2603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9423_ _0209_ clknet_leaf_55_clk reg_file.reg_storage\[13\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4896_ _0811_ reg_file.reg_storage\[3\]\[21\] _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7684_ net19 _3138_ _3498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6635_ _2518_ _2534_ _2535_ _2536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_27_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer25_I _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9354_ _0140_ clknet_leaf_7_clk reg_file.reg_storage\[7\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _2338_ _2469_ _2052_ _2470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5517_ _1432_ reg_file.reg_storage\[2\]\[27\] _1427_ _1433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8305_ _3674_ _3977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_76_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9285_ _0071_ clknet_leaf_38_clk reg_file.reg_storage\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5672__I _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6497_ _2397_ _2402_ _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8236_ _3454_ _3926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input52_I mem_ld_dat[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5448_ _1363_ _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8167_ _3867_ _3882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5379_ _0850_ _1295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7118_ _1664_ _2989_ _2994_ net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8098_ reg_file.reg_storage\[2\]\[15\] _3624_ _3821_ _3839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7237__A2 _3081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output139_I net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7049_ _2930_ net214 _2086_ _2935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5248__A1 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4606__S0 _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6920__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6678__I _2304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5031__S0 _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7476__A2 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8893__I _4359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__C _3472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5239__A1 _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4926__I _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_4_7_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4750_ _0586_ _0661_ _0662_ _0663_ _0665_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_28_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7164__A1 _1475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7164__B2 _1729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4681_ net27 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9165__S _4522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6911__A1 _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6420_ _2065_ _2114_ _2328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6351_ _2214_ _2261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5302_ _0834_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_122_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9070_ _3932_ _4462_ _4469_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6282_ _2121_ _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5425__C _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8021_ _3657_ _3784_ _3790_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_58_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5233_ _1147_ _1148_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5164_ reg_file.reg_storage\[12\]\[26\] reg_file.reg_storage\[13\]\[26\] reg_file.reg_storage\[14\]\[26\]
+ reg_file.reg_storage\[15\]\[26\] _0921_ _0922_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_71_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5095_ _1010_ _0875_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8923_ reg_file.reg_storage\[9\]\[12\] _4209_ _4365_ _4379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8854_ _4310_ _4336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5650__A1 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5089__S0 _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7805_ _3610_ _3611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8785_ _4234_ _4263_ _4293_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5997_ _1268_ _1910_ _1911_ _1912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4571__I _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7736_ _0595_ _3524_ _3546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4948_ _0863_ reg_file.reg_storage\[2\]\[23\] _0764_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7667_ net60 net37 net46 net54 _3481_ _3461_ _3482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_129_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4879_ _0794_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9144__A2 _4512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9406_ _0192_ clknet_leaf_87_clk reg_file.reg_storage\[13\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6618_ _2135_ _2250_ _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7598_ _1901_ _3417_ _3418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6498__I _2086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9337_ _0123_ clknet_leaf_104_clk reg_file.reg_storage\[6\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6549_ _2161_ _2162_ _2205_ _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_30_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9268_ _0054_ clknet_leaf_27_clk reg_file.reg_storage\[3\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_9199_ _3992_ _4506_ _4545_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8219_ _3420_ _3911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_7_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_88_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_131_clk_I clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_11_clk_I clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8154__S _3873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_26_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5944__A2 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7146__A1 net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5180__I0 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_127_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8949__A2 _4363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5307__S1 _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__B2 _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A1 _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ _1194_ _1835_ _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4592__S _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ _1293_ _1766_ _1767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_8570_ reg_file.reg_storage\[12\]\[16\] _4141_ _4150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_122_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ reg_file.reg_storage\[1\]\[13\] _1697_ _1695_ _1698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4802_ _0717_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9126__A2 _4496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7521_ _3344_ _3345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4733_ net10 _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_138_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7452_ _3248_ net110 _3283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6312__S _2105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5243__S0 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4664_ reg_file.reg_storage\[4\]\[7\] reg_file.reg_storage\[5\]\[7\] reg_file.reg_storage\[6\]\[7\]
+ reg_file.reg_storage\[7\]\[7\] _0566_ _0567_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_71_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6403_ _1265_ _2234_ _2311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_101_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6360__A2 _2269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4595_ reg_file.reg_storage\[4\]\[1\] reg_file.reg_storage\[5\]\[1\] reg_file.reg_storage\[6\]\[1\]
+ reg_file.reg_storage\[7\]\[1\] _0480_ _0518_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_7383_ net71 _3205_ _3219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9122_ reg_file.reg_storage\[4\]\[27\] _4496_ _4499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6334_ _2236_ _2243_ _2244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9053_ _4454_ _4457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6265_ _2045_ _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8239__S _3928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8004_ reg_file.reg_storage\[3\]\[11\] _3568_ _3775_ _3781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5216_ _1131_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6196_ _1786_ _2109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5147_ _1062_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4566__I _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5078_ _0754_ _0993_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5623__A1 _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8906_ _4191_ _4362_ _4369_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input15_I inst[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8837_ reg_file.reg_storage\[10\]\[10\] _4205_ _4322_ _4327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7376__A1 _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8768_ reg_file.reg_storage\[11\]\[16\] _4275_ _4284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5926__A2 _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9117__A2 _4456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7719_ _3530_ _3531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_81_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8699_ _3709_ _4238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__S1 _1536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5154__A3 _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5537__S1 _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8800__A1 reg_file.reg_storage\[11\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5917__A2 _1832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5473__S0 _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9108__A2 _4486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6342__A2 _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _0886_ _1964_ _1965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5001_ _0897_ _0915_ _0916_ _0893_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4656__A2 _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input7_I inst[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7697__I _3509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__A1 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5700__S1 _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6952_ _2841_ _2142_ _1072_ _2842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9671_ _0457_ clknet_leaf_35_clk reg_file.reg_storage\[15\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6883_ _1838_ _2539_ _2775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5903_ _1817_ _1818_ _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_49_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ reg_file.reg_storage\[4\]\[9\] reg_file.reg_storage\[5\]\[9\] reg_file.reg_storage\[6\]\[9\]
+ reg_file.reg_storage\[7\]\[9\] _1590_ _1642_ _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_66_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8622_ _4177_ _4182_ _4184_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4967__I0 net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8553_ _4140_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8321__I _3704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5765_ _1670_ _1671_ _1680_ _1681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_45_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5696_ reg_file.reg_storage\[2\]\[18\] reg_file.reg_storage\[3\]\[18\] _1611_ _1612_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8484_ _4096_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7504_ _3329_ _3320_ _3316_ _3330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4716_ net7 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_142_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6869__B1 _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4647_ _0483_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7435_ net75 _3253_ _3267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7366_ _3192_ _1710_ _3203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9105_ _3973_ _4488_ _4489_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4578_ reg_file.reg_storage\[2\]\[0\] reg_file.reg_storage\[3\]\[0\] _0503_ _0504_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6317_ _1997_ _2208_ _2221_ _2227_ _2228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5680__I _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5519__S1 _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8086__A2 _3818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7297_ _3127_ _3129_ _3140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7833__A2 _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_15_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9036_ _3992_ _4445_ _4446_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6248_ _2156_ _2159_ _1292_ _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6179_ _2090_ _2091_ _2092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output121_I net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6217__S _2022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5455__S0 _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__A1 _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_97_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8231__I _3921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8077__A2 _3819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9026__A1 _3980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5694__S0 _1607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6260__A1 _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8001__A2 _3765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_70_clk clknet_4_9_0_clk clknet_leaf_70_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6563__A2 _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5550_ reg_file.reg_storage\[4\]\[31\] reg_file.reg_storage\[5\]\[31\] reg_file.reg_storage\[6\]\[31\]
+ reg_file.reg_storage\[7\]\[31\] _1464_ _1465_ _1466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_14_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5481_ _0492_ _1396_ _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_81_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7220_ _1108_ _3069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6315__A2 _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7151_ net163 _2979_ _3016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7082_ _2966_ net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6102_ _1120_ _2016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7815__A2 _3202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5826__A1 _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6033_ _1947_ _0851_ _1948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5005__I _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer12 _0656_ net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4844__I _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer34 _1648_ net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XTAP_TAPCELL_ROW_68_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7984_ reg_file.reg_storage\[3\]\[2\] _3456_ _3769_ _3770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xrebuffer23 _0883_ net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_95_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6935_ _1878_ _2807_ _2074_ _2825_ _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_81_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_61_clk clknet_4_11_0_clk clknet_leaf_61_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_119_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9654_ _0440_ clknet_leaf_113_clk reg_file.reg_storage\[4\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6866_ _2742_ _1844_ _2759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8605_ _4013_ _4122_ _4169_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9585_ _0371_ clknet_leaf_67_clk reg_file.reg_storage\[9\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6797_ _2585_ _2692_ _2492_ _2693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5817_ _1694_ _1708_ _1721_ _1732_ _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_18_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5748_ _0490_ _1663_ _1664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_91_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8051__I net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8536_ _3919_ _4128_ _4130_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_134_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4660__S1 _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input82_I pc[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5679_ _1531_ _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_114_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9083__S _4472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8467_ reg_file.reg_storage\[13\]\[8\] _3943_ _4085_ _4087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_79_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8398_ _4024_ _4044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7418_ net74 _3233_ _3251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_92_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8059__A2 _3812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7349_ _3165_ _1692_ _3188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7806__A2 _3544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9019_ _3969_ _4430_ _4436_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5132__I3 reg_file.reg_storage\[7\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6242__A1 _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6793__A2 _2470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_52_clk clknet_4_10_0_clk clknet_leaf_52_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_0_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7742__A1 _1671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8896__I _4359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8298__A2 _3971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5600__S0 _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5108__I0 reg_file.reg_storage\[8\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8470__A2 _4088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6365__B _2274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4981_ _0896_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5696__S _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7908__C _3703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_43_clk clknet_4_8_0_clk clknet_leaf_43_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6720_ _2617_ _2578_ _2618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4795__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6651_ _2551_ _1839_ _2496_ _2552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_63_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9370_ _0156_ clknet_leaf_98_clk reg_file.reg_storage\[7\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_119_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5602_ _1512_ _1515_ _1516_ _1517_ _1455_ _1395_ _1518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_73_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6582_ _1693_ _2485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8321_ _3704_ _3989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5533_ reg_file.reg_storage\[2\]\[24\] reg_file.reg_storage\[3\]\[24\] _1360_ _1449_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8289__A2 _3947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8252_ _3937_ _3938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5464_ net25 _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_8183_ reg_file.reg_storage\[6\]\[16\] _3882_ _3891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7203_ net65 _0689_ _3054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5395_ _1310_ _1030_ _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7134_ net145 _3004_ _3005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7065_ _2950_ net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6016_ _1929_ _1930_ _1931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5275__A2 _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4574__I _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5658__S0 _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7967_ _3753_ _3754_ _3755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9078__S _4472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7972__A1 _3421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_34_clk clknet_4_2_0_clk clknet_leaf_34_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_76_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6918_ _2807_ _2808_ _2809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7898_ net112 _3446_ _3692_ _3694_ _3695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_25_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4786__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9637_ _0423_ clknet_leaf_39_clk reg_file.reg_storage\[4\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6849_ _0874_ _2742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5050__I2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5830__S0 _1590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9568_ _0354_ clknet_leaf_127_clk reg_file.reg_storage\[9\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8519_ reg_file.reg_storage\[13\]\[31\] _4068_ _4116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9499_ _0285_ clknet_leaf_100_clk reg_file.reg_storage\[8\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5266__A2 _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7795__I _3472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_25_clk clknet_4_3_0_clk clknet_leaf_25_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__9004__I1 _3584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4777__A1 _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6518__A2 _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4624__S1 _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7191__A2 _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7744__B _3553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_3_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer3 net210 net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8140__A1 reg_file.reg_storage\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4659__I _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8691__A2 _4181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5180_ _1089_ _1093_ _1094_ _1095_ _0870_ _1025_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__7651__B1 _3463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8870_ reg_file.reg_storage\[10\]\[25\] _4307_ _4345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6206__A1 _2117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7821_ _3625_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7752_ _3517_ _3560_ _3561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_125_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_16_clk clknet_4_0_0_clk clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4964_ net31 _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_117_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6703_ _2424_ _2368_ _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_22_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9422_ _0208_ clknet_leaf_55_clk reg_file.reg_storage\[13\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4895_ _0810_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_46_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7683_ _3496_ _3497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_144_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6634_ _2533_ _2514_ _2535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_61_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9353_ _0139_ clknet_leaf_50_clk reg_file.reg_storage\[7\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5812__S0 _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6565_ _2297_ _2381_ _2468_ _2469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5516_ _1431_ _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8304_ _3974_ _3975_ _3976_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9284_ _0070_ clknet_leaf_19_clk reg_file.reg_storage\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6496_ _1669_ _1681_ _2401_ _2402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_5447_ _1362_ _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8131__A1 _3740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8235_ _3919_ _3923_ _3925_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4569__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer18_I _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8682__A2 _4223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input45_I mem_ld_dat[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8166_ _3881_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7890__B1 _3685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5378_ _1293_ _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7117_ net159 _2992_ _2994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8097_ _3611_ _3837_ _3838_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7048_ _2885_ _2890_ _2909_ _2933_ _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8999_ _3945_ _4411_ _4425_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7796__I1 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5420__A2 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__A1 _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__A1 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5031__S1 _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6694__I _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5304__S _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5411__A2 _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4680_ _0596_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_141_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5175__A1 _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6911__A2 _2802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6350_ _2249_ _2252_ _2256_ _2257_ _2259_ _2260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_52_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8113__A1 _3682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5301_ _1216_ _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6281_ _2192_ _2193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8020_ reg_file.reg_storage\[3\]\[18\] _3789_ _3790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6675__A1 _2573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6818__B _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5232_ _0830_ _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_5_clk clknet_4_6_0_clk clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5163_ _0954_ _1076_ _1077_ _1078_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8416__A2 _4051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5094_ _1009_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8922_ _4378_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5013__I _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8853_ _4220_ _4331_ _4335_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5650__A2 _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5089__S1 _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7804_ net102 _3601_ _3606_ _3609_ _3610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_93_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4852__I _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8784_ reg_file.reg_storage\[11\]\[23\] _4261_ _4293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5996_ _0791_ _1148_ _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7735_ _3428_ _3543_ _3545_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4947_ _0771_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7666_ _3026_ _3481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8260__S _3941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4878_ _0793_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_34_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9405_ _0191_ clknet_leaf_88_clk reg_file.reg_storage\[14\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6202__I1 _2113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6617_ _2509_ _2514_ _2518_ _2519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_144_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9336_ _0122_ clknet_leaf_104_clk reg_file.reg_storage\[6\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7597_ _3416_ _3417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_120_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6548_ _2093_ _2091_ _2452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9267_ _0053_ clknet_leaf_25_clk reg_file.reg_storage\[3\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6479_ _2332_ _2384_ _2385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9198_ reg_file.reg_storage\[15\]\[25\] _4507_ _4545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8218_ _3751_ _3863_ _3910_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6666__A1 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output151_I net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_144_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8149_ _3443_ _3869_ _3871_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_89_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7394__A2 _3228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8170__S _3879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7313__I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5880__A2 _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ _1765_ _1766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_122_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9176__S _4515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7983__I _3768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5781_ reg_file.reg_storage\[2\]\[13\] reg_file.reg_storage\[3\]\[13\] _1611_ _1697_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5396__A1 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4801_ _0714_ _0715_ _0716_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_90_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8080__S _3828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7520_ net85 _3344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4732_ _0625_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_32_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4663_ reg_file.reg_storage\[12\]\[7\] reg_file.reg_storage\[13\]\[7\] reg_file.reg_storage\[14\]\[7\]
+ reg_file.reg_storage\[15\]\[7\] _0566_ _0567_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_43_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7451_ _3053_ _3281_ _3282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5243__S1 _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5209__S _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6896__A1 _2742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6402_ _2235_ _2279_ _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7382_ _3215_ _3217_ _3218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4594_ reg_file.reg_storage\[12\]\[1\] reg_file.reg_storage\[13\]\[1\] reg_file.reg_storage\[14\]\[1\]
+ reg_file.reg_storage\[15\]\[1\] _0480_ _0518_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_9121_ _4455_ _4498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6333_ _2238_ _2242_ _2243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9052_ _4455_ _4456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6264_ _2065_ _2176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8003_ _3780_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5215_ _1121_ _1130_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_86_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6195_ _2103_ _2105_ _2107_ _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5146_ net8 _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__9062__A2 _4462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4674__A3 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5077_ _0985_ _0989_ _0991_ _0992_ _0786_ _0929_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_98_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8905_ reg_file.reg_storage\[9\]\[4\] _4363_ _4369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8836_ _4202_ _4312_ _4326_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_11_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8767_ _4283_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ _1873_ _0721_ _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7718_ _3529_ _3530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8698_ _4236_ _4174_ _4237_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8876__A2 _4346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7649_ _3416_ _3466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_132_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9319_ _0105_ clknet_leaf_34_clk reg_file.reg_storage\[6\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7300__A2 net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A2 _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8165__S _3879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6575__B1 _2466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8899__I _4359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5473__S1 _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8867__A2 _4313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4667__I _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _0892_ reg_file.reg_storage\[3\]\[16\] _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7978__I _3764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8075__S _3822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__A2 _1511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_72_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6951_ _1085_ _2841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9670_ _0456_ clknet_leaf_43_clk reg_file.reg_storage\[15\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6882_ _2770_ _2771_ _2772_ _2773_ _2774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_5902_ _1693_ _1818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5833_ reg_file.reg_storage\[12\]\[9\] reg_file.reg_storage\[13\]\[9\] reg_file.reg_storage\[14\]\[9\]
+ reg_file.reg_storage\[15\]\[9\] _0685_ _1623_ _1749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_8621_ reg_file.reg_storage\[8\]\[1\] _4183_ _4184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_87_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8552_ reg_file.reg_storage\[12\]\[8\] _3943_ _4138_ _4140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_66_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5764_ _0670_ _1679_ _1680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7503_ _3318_ _3329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8858__A2 _4336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5695_ _0685_ _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_8483_ reg_file.reg_storage\[13\]\[15\] _3961_ _4078_ _4096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4715_ _0630_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__7218__I net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_130_clk_I clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6869__A1 _2742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4646_ _0503_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7434_ net75 _3253_ _3266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_21_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5541__A1 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7365_ net71 _3201_ _3202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_4_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4577_ _0502_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_97_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9104_ reg_file.reg_storage\[4\]\[19\] _4486_ _4489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6316_ _2192_ _2225_ _2226_ _1345_ _2227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7296_ _3122_ net21 _3138_ _3139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4577__I _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9035_ reg_file.reg_storage\[1\]\[25\] _4443_ _4446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_25_clk_I clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6247_ _0743_ _2157_ _2158_ _2159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6178_ _1777_ _2089_ _2091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5844__A2 _1759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5129_ _1012_ _1044_ _0886_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5152__S0 _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output114_I net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7349__A2 _1692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8819_ reg_file.reg_storage\[10\]\[2\] _4185_ _4316_ _4317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_15_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5455__S1 _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_97_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9026__A2 _4437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__S0 _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5694__S1 _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6260__A2 _2171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4950__I _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5480_ _1389_ _1392_ _1393_ _1394_ _1372_ _1395_ _1396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_41_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7150_ _3014_ _3012_ _3015_ net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_117_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7081_ _2352_ _2953_ _2965_ _2966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6101_ _2005_ _2009_ _2014_ _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__5826__A2 _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6032_ _1310_ _1947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xrebuffer35 net238 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XTAP_TAPCELL_ROW_68_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7983_ _3768_ _3769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xrebuffer24 net226 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer13 _0675_ net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6934_ _2269_ _2080_ _1399_ _2825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5021__I _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9653_ _0439_ clknet_leaf_118_clk reg_file.reg_storage\[4\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8604_ reg_file.reg_storage\[12\]\[31\] _4120_ _4169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _2000_ _2302_ _2750_ _2757_ _2758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_77_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9584_ _0370_ clknet_leaf_68_clk reg_file.reg_storage\[9\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5816_ _1175_ _1731_ _1732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_57_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6796_ _2587_ _2691_ _2183_ _2692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5747_ _1658_ _1660_ _1661_ _1662_ _1595_ _1596_ _1663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8535_ reg_file.reg_storage\[12\]\[1\] _4129_ _4130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8466_ _4086_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5678_ reg_file.reg_storage\[4\]\[16\] reg_file.reg_storage\[5\]\[16\] reg_file.reg_storage\[6\]\[16\]
+ reg_file.reg_storage\[7\]\[16\] _1587_ _1420_ _1594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5514__A1 _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input75_I pc[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7417_ _3041_ _3250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_20_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5691__I _1606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4629_ _0510_ _0550_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8397_ _4043_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7348_ _3185_ _3186_ _3187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7279_ _3122_ _3112_ _3123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__7267__A1 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9018_ reg_file.reg_storage\[1\]\[18\] _4435_ _4436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5373__S0 _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8507__I _4067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9569__CLK clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4971__S _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6242__A2 _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4770__I _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7742__A2 _3402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5087__B _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5753__A1 _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5600__S1 _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5108__I1 reg_file.reg_storage\[9\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5106__I _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5116__S0 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6769__B1 _2651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6233__A2 _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4980_ _0854_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_58_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7981__A2 _3765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6650_ _2532_ _2551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_63_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5601_ reg_file.reg_storage\[8\]\[28\] reg_file.reg_storage\[9\]\[28\] reg_file.reg_storage\[10\]\[28\]
+ reg_file.reg_storage\[11\]\[28\] _1446_ _1447_ _1517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6581_ _2439_ _2484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_119_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5532_ reg_file.reg_storage\[4\]\[24\] reg_file.reg_storage\[5\]\[24\] reg_file.reg_storage\[6\]\[24\]
+ reg_file.reg_storage\[7\]\[24\] _1446_ _1447_ _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8320_ _3987_ _3924_ _3988_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7924__C _3717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8251_ _3501_ _3937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5463_ _1378_ _1379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_8182_ _3890_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7202_ _3052_ _3053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5394_ _1309_ _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7133_ _3001_ _3004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7249__B2 _3095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7064_ _2936_ _2949_ _2950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6472__A2 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _1098_ _0850_ _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4855__I _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5107__S0 _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7421__A1 _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7966_ _0880_ _3396_ _3754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6917_ _2797_ _2767_ _2484_ _2808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6291__B _2202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7897_ _3671_ _3294_ _3499_ _3693_ _3694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_25_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6848_ _1852_ _2722_ _2741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_76_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8062__I _3816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9636_ _0422_ clknet_leaf_17_clk reg_file.reg_storage\[4\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8997__I _4414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9567_ _0353_ clknet_leaf_123_clk reg_file.reg_storage\[9\]\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8518_ _4010_ _4111_ _4115_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6779_ _2672_ _2674_ _2675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9094__S _4465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9498_ _0284_ clknet_leaf_99_clk reg_file.reg_storage\[8\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5830__S1 _1642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8449_ _4072_ _4076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output181_I net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7488__A1 _3144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5346__S0 _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7660__A1 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5797__S _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4777__A2 _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8901__S _4366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7715__A2 _3123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer4 _2400_ net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7479__A1 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_39_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6454__A2 _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7651__A1 _2148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7820_ reg_file.reg_storage\[5\]\[15\] _3624_ _3569_ _3625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7403__A1 _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7954__A2 _3370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7751_ _3518_ _3031_ net52 _3560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_125_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4963_ _0878_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_86_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6702_ _2598_ _2600_ _2601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_58_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7682_ _3429_ _3437_ _3496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_117_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4894_ _0809_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9421_ _0207_ clknet_leaf_12_clk reg_file.reg_storage\[13\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6633_ _2533_ _2514_ _2534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5717__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9352_ _0138_ clknet_leaf_49_clk reg_file.reg_storage\[7\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5812__S1 _1596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6564_ _2011_ _2467_ _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8303_ reg_file.reg_storage\[7\]\[19\] _3971_ _3976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6495_ _2398_ net207 _2401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5515_ _0688_ _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9283_ _0069_ clknet_leaf_0_clk reg_file.reg_storage\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5446_ _1361_ _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_76_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6130__I _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8234_ reg_file.reg_storage\[7\]\[1\] _3924_ _3925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5576__S0 _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8165_ reg_file.reg_storage\[6\]\[8\] _3531_ _3879_ _3881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7890__A1 net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7890__B2 _3687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5377_ _1292_ _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7116_ _1679_ _2989_ _2993_ net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8096_ reg_file.reg_storage\[2\]\[14\] _3831_ _3838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input38_I mem_ld_dat[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5099__I3 reg_file.reg_storage\[7\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ _2905_ _2908_ _2932_ _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_2_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8198__A2 _3895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9089__S _4465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8998_ reg_file.reg_storage\[1\]\[9\] _4424_ _4425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7949_ _3739_ _3740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5956__A1 _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4759__A2 _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9619_ _0405_ clknet_leaf_76_clk reg_file.reg_storage\[1\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7136__I _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__I _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6684__A2 _2339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8189__A2 _3888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9287__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8984__I1 _3469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9138__A1 _3761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8113__A2 _3844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _1215_ _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5558__S0 _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6280_ _1790_ _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_121_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6675__A2 _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5231_ _1146_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5162_ _0957_ reg_file.reg_storage\[2\]\[26\] _0958_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_71_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5093_ _0998_ _1008_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8921_ reg_file.reg_storage\[9\]\[11\] _4207_ _4372_ _4378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_56_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8852_ reg_file.reg_storage\[10\]\[17\] _4325_ _4335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5938__A1 _1852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8783_ _4232_ _4288_ _4292_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7803_ _3607_ _3194_ _3446_ _3608_ _3609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__9129__A1 _4009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7734_ reg_file.reg_storage\[5\]\[9\] _3544_ _3545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5995_ _0968_ _1163_ _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8541__S _4132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _0861_ reg_file.reg_storage\[3\]\[23\] _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_35_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7665_ net124 _3480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4877_ _0792_ _0660_ _0675_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9404_ _0190_ clknet_leaf_96_clk reg_file.reg_storage\[14\]\[30\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8340__I _4003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer30_I _1519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6616_ _2443_ _2461_ _2489_ _2517_ _2518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7596_ _3391_ _3416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9335_ _0121_ clknet_leaf_114_clk reg_file.reg_storage\[6\]\[25\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_65_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6547_ _2444_ _2450_ _2451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9266_ _0052_ clknet_leaf_72_clk reg_file.reg_storage\[3\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7312__B1 _3144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6478_ _2263_ _2383_ _2109_ _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9197_ _3989_ _4506_ _4544_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8217_ reg_file.reg_storage\[6\]\[31\] _3861_ _3910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7863__B2 _3253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5429_ net24 _0704_ _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8148_ reg_file.reg_storage\[6\]\[1\] _3870_ _3871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output144_I net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5477__I0 reg_file.reg_storage\[12\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8079_ _3816_ _3828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_69_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A1 _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7854__A1 net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7854__B2 _3655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7606__A1 _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5114__I _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8626__S _4187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5468__I0 _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5712__S0 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8425__I _4016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8582__A2 _4152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4800_ _0706_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_122_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5780_ reg_file.reg_storage\[8\]\[13\] reg_file.reg_storage\[9\]\[13\] reg_file.reg_storage\[10\]\[13\]
+ reg_file.reg_storage\[11\]\[13\] _0687_ _1695_ _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4731_ reg_file.reg_storage\[8\]\[0\] reg_file.reg_storage\[9\]\[0\] reg_file.reg_storage\[10\]\[0\]
+ reg_file.reg_storage\[11\]\[0\] _0644_ _0645_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_56_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4662_ reg_file.reg_storage\[1\]\[7\] _0580_ _0578_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7450_ _3275_ _3278_ _3280_ _3281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_142_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6401_ _2309_ net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_3_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9120_ _3995_ _4456_ _4497_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7381_ _3188_ _3216_ _3186_ _3217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4593_ _0482_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_141_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7932__C _3724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6332_ _2240_ _2241_ _2242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7845__A1 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7845__B2 _3647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9051_ _4454_ _4455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6263_ _1768_ _2169_ _2172_ _2174_ _2175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_3_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8002_ reg_file.reg_storage\[3\]\[10\] _3557_ _3775_ _3780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5214_ _0912_ _0938_ _1129_ _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6194_ _2106_ _2107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5145_ _0940_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5024__I _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5076_ reg_file.reg_storage\[8\]\[28\] reg_file.reg_storage\[9\]\[28\] reg_file.reg_storage\[10\]\[28\]
+ reg_file.reg_storage\[11\]\[28\] _0990_ _0984_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__8335__I _3999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4863__I _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6820__A2 _1542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8904_ _4368_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8573__A2 _4147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8835_ reg_file.reg_storage\[10\]\[9\] _4325_ _4326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8271__S _3941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8766_ reg_file.reg_storage\[11\]\[15\] _4216_ _4265_ _4283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5978_ _1872_ _1875_ _1893_ _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_19_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7717_ _2350_ _3504_ _3528_ _3529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_8697_ reg_file.reg_storage\[8\]\[24\] _4175_ _4237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4929_ _0838_ _0841_ _0843_ _0844_ _0785_ _0825_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_90_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7648_ _3047_ _3068_ _3465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7579_ _3398_ _3399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9318_ _0104_ clknet_leaf_42_clk reg_file.reg_storage\[6\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7836__A1 _3600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9249_ _0035_ clknet_leaf_130_clk reg_file.reg_storage\[3\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5135__S _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8181__S _3872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6575__B2 _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8316__A2 _3975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__I _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5779__I _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6950_ _2833_ _2838_ _2351_ _2840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5066__A1 net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5901_ _1131_ _1817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6881_ _2533_ _2514_ _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8555__A2 _4141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5832_ reg_file.reg_storage\[1\]\[9\] _1747_ _1642_ _1748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8091__S _3821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8620_ _4179_ _4183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_17_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ _1604_ _1678_ _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_8551_ _4139_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_66_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8307__A2 _3971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7502_ _3326_ _3327_ _3328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4714_ _0624_ _0625_ _0626_ _0629_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_8482_ _3958_ _4094_ _4095_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_127_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5694_ reg_file.reg_storage\[8\]\[18\] reg_file.reg_storage\[9\]\[18\] reg_file.reg_storage\[10\]\[18\]
+ reg_file.reg_storage\[11\]\[18\] _1607_ _1609_ _1610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_16_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4645_ _0565_ net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_112_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7433_ _3240_ _3244_ _3254_ _3238_ _3265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_97_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7364_ _3192_ _3193_ _3201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4576_ net13 _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4858__I _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9103_ _4466_ _4488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6315_ _1281_ _1805_ _0718_ _1764_ _1344_ _2226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_9034_ _4405_ _4445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7295_ _1443_ _3138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7294__A2 _1829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6246_ _1110_ _1240_ _0884_ _0794_ _2158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6177_ _1800_ _2089_ _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5128_ _1029_ _1030_ _1043_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_input20_I inst[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__I _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5152__S1 _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5059_ net32 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_95_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output107_I net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6557__A1 _2458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8818_ _4315_ _4316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_109_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8749_ _4273_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4663__S0 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4768__I _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8176__S _3872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6493__B1 _1829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__S1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8785__A2 _4263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_106_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8703__I _4172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4654__S0 _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_109_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4678__I _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5283__B _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6100_ _2010_ _2013_ _2014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7080_ _2641_ _2960_ _2964_ _2965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7276__A2 _3115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6031_ _1795_ _1295_ _1946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8225__A1 reg_file.reg_storage\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8776__A2 _4286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer25 _1598_ net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer36 net239 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_68_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7982_ _3762_ _3768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xrebuffer14 net232 net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6933_ _2421_ _2370_ _2823_ _2582_ _2824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_89_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6864_ _2324_ _2756_ _2210_ _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9652_ _0438_ clknet_leaf_24_clk reg_file.reg_storage\[4\]\[22\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6539__A1 _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8603_ _4010_ _4164_ _4168_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5815_ _1670_ _1722_ _1730_ _1731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_9_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9583_ _0369_ clknet_leaf_64_clk reg_file.reg_storage\[9\]\[17\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6795_ _2636_ _2690_ _2008_ _2691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__I _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5746_ reg_file.reg_storage\[4\]\[11\] reg_file.reg_storage\[5\]\[11\] reg_file.reg_storage\[6\]\[11\]
+ reg_file.reg_storage\[7\]\[11\] _0686_ _1588_ _1662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8534_ _4125_ _4129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5677_ reg_file.reg_storage\[12\]\[16\] reg_file.reg_storage\[13\]\[16\] reg_file.reg_storage\[14\]\[16\]
+ reg_file.reg_storage\[15\]\[16\] _1587_ _1420_ _1593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8465_ reg_file.reg_storage\[13\]\[7\] _3940_ _4085_ _4086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4628_ reg_file.reg_storage\[4\]\[4\] reg_file.reg_storage\[5\]\[4\] reg_file.reg_storage\[6\]\[4\]
+ reg_file.reg_storage\[7\]\[4\] _0480_ _0518_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7416_ _3248_ net107 _3249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_20_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input68_I pc[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4588__I _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8396_ reg_file.reg_storage\[14\]\[13\] _3955_ _4028_ _4043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4559_ net15 _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7347_ net69 _3183_ _3186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_92_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7278_ net95 _3122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7267__A2 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9017_ _4409_ _4435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6229_ _1924_ _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8216__A1 _3746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5373__S1 _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6778__A1 _1707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6242__A3 _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9192__A2 _4511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5202__A1 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__A2 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_71_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5108__I2 reg_file.reg_storage\[10\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_86_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8207__A1 _3719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5116__S1 _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6769__A1 _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9183__A2 _4536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5600_ reg_file.reg_storage\[12\]\[28\] reg_file.reg_storage\[13\]\[28\] reg_file.reg_storage\[14\]\[28\]
+ reg_file.reg_storage\[15\]\[28\] _1446_ _1447_ _1516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_clkbuf_leaf_24_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6580_ _1707_ _2483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5531_ _1363_ _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_119_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8250_ _3936_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_39_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5462_ _1115_ _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_120_clk clknet_4_7_0_clk clknet_leaf_120_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7201_ _3038_ _3052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8181_ reg_file.reg_storage\[6\]\[15\] _3624_ _3872_ _3890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5393_ _1300_ _0621_ _1218_ _1308_ _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_7132_ net228 _3000_ _3003_ net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7249__A2 net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7063_ _2254_ _2849_ _2940_ _2948_ _2949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_94_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6014_ _0996_ _1163_ _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5107__S1 _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7421__A2 _3253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8343__I _3739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__S0 _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4871__I _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7965_ _0975_ net2 _3753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__9174__A2 _4525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6916_ _1879_ _2807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7896_ _3295_ _3464_ _3693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_25_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6847_ _2740_ net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9635_ _0421_ clknet_leaf_0_clk reg_file.reg_storage\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9566_ _0352_ clknet_leaf_110_clk reg_file.reg_storage\[9\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6778_ _1707_ _2486_ _2563_ _2673_ _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_9_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8517_ reg_file.reg_storage\[13\]\[30\] _4068_ _4115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5729_ _1644_ _1622_ _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_80_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9497_ _0283_ clknet_leaf_101_clk reg_file.reg_storage\[8\]\[27\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8448_ _4074_ _4075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5499__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5207__I _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8379_ _4033_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6999__A1 _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5346__S1 _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8454__S _4079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6482__B _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5974__A2 _1519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7176__A1 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer5 _2400_ net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_102_clk clknet_4_15_0_clk clknet_leaf_102_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7479__A2 _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8629__S _4187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8979__A2 _4411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7100__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5662__A1 _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7750_ net35 net43 _3027_ _3559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_125_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4962_ _0483_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7681_ net129 _3494_ _3495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6701_ _2561_ _2567_ _2599_ _2600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9156__A2 _4512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4893_ _0755_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9420_ _0206_ clknet_leaf_54_clk reg_file.reg_storage\[13\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6632_ _1162_ _2533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5273__S0 _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6914__A1 _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9351_ _0137_ clknet_leaf_34_clk reg_file.reg_storage\[7\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ _2432_ _2142_ _1133_ _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_15_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5514_ _1429_ reg_file.reg_storage\[3\]\[27\] _1430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8302_ _3928_ _3975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9282_ _0068_ clknet_leaf_19_clk reg_file.reg_storage\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6494_ _2154_ _2232_ _2317_ _2399_ _2400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5445_ _0539_ _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_76_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8233_ _3920_ _3924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8539__S _4132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5576__S1 _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8164_ _3880_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7115_ net156 _2992_ _2993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7890__A2 _3661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ _1218_ _1290_ _1291_ _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8095_ _3817_ _3837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7046_ _2883_ _2931_ _2932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8274__S _3927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8997_ _4414_ _4424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5405__A1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7948_ net118 _3728_ _3729_ _3736_ _3738_ _3739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_96_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7879_ _3632_ _3677_ _3652_ _3678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_108_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9618_ _0404_ clknet_leaf_72_clk reg_file.reg_storage\[1\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9549_ _0335_ clknet_leaf_12_clk reg_file.reg_storage\[10\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output99_I net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5192__I0 _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8248__I _3489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8912__S _4372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5947__A2 _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7149__A1 net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5255__S0 _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5007__S0 _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5558__S1 _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5230_ _1134_ _0912_ _1145_ _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7321__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5161_ _0768_ reg_file.reg_storage\[3\]\[26\] _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5092_ _0891_ _1007_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8920_ _4377_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_3_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8851_ _4218_ _4331_ _4334_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9231__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8782_ reg_file.reg_storage\[11\]\[22\] _4261_ _4292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5994_ _0949_ _0951_ _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7802_ _1710_ _3439_ _3608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9129__A2 _4498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7733_ _3457_ _3544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4945_ _0860_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_86_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7664_ _3428_ _3478_ _3479_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4876_ _0668_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_7_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9403_ _0189_ clknet_leaf_96_clk reg_file.reg_storage\[14\]\[29\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7595_ _3410_ _3413_ _3414_ _3415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_90_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6363__A2 _2265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6615_ _2494_ _2488_ _2516_ _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9334_ _0120_ clknet_leaf_114_clk reg_file.reg_storage\[6\]\[24\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6546_ _2396_ _2445_ _2447_ _2448_ _2449_ _2316_ _2450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XANTENNA_rebuffer23_I _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9265_ _0051_ clknet_leaf_72_clk reg_file.reg_storage\[3\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7312__B2 _3146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7312__A1 _3035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6477_ _2037_ _2381_ _2382_ _2383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input50_I mem_ld_dat[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9196_ reg_file.reg_storage\[15\]\[24\] _4507_ _4544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8216_ _3746_ _3905_ _3909_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_7_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7863__A2 _3252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5428_ _0721_ _1344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8147_ _3866_ _3870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8068__I _3821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5359_ reg_file.reg_storage\[12\]\[5\] reg_file.reg_storage\[13\]\[5\] reg_file.reg_storage\[14\]\[5\]
+ reg_file.reg_storage\[15\]\[5\] _0637_ _0634_ _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4596__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5874__A1 _1787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8078_ _3502_ _3818_ _3827_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5477__I1 reg_file.reg_storage\[13\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7029_ _2212_ _2796_ _2915_ _2916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output137_I net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7854__A2 _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9056__A1 _3424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8907__S _4366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__I3 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__S1 _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8706__I _3725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__A1 _1767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8642__S _4198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8031__A2 _3764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5130__I net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6042__A1 _1955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4730_ reg_file.reg_storage\[12\]\[0\] reg_file.reg_storage\[13\]\[0\] reg_file.reg_storage\[14\]\[0\]
+ reg_file.reg_storage\[15\]\[0\] _0644_ _0645_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_44_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4661_ reg_file.reg_storage\[2\]\[7\] reg_file.reg_storage\[3\]\[7\] _0497_ _0580_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6345__A2 _2254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5228__S0 _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6400_ _2087_ _2283_ _2295_ _2296_ _2308_ _2309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7380_ _3180_ _3184_ _3216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_12_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6331_ _1280_ _2239_ _2160_ _2241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4592_ reg_file.reg_storage\[1\]\[1\] _0516_ _0514_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8089__S _3828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7845__A2 _3601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9050_ _3388_ _4118_ _4454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6262_ _2173_ _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9047__A1 _4009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8001_ _3543_ _3765_ _3779_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5213_ _1124_ _1126_ _1127_ _1128_ _0822_ _0871_ _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_6193_ _1253_ _2106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5144_ net82 _0852_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5075_ reg_file.reg_storage\[12\]\[28\] reg_file.reg_storage\[13\]\[28\] reg_file.reg_storage\[14\]\[28\]
+ reg_file.reg_storage\[15\]\[28\] _0990_ _0984_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__7520__I net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8903_ reg_file.reg_storage\[9\]\[3\] _4189_ _4366_ _4368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8552__S _4138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8834_ _4310_ _4325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_91_clk clknet_4_14_0_clk clknet_leaf_91_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6033__A1 _1947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8765_ _4213_ _4281_ _4282_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6584__A2 _2486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5977_ _1888_ _1892_ _1873_ net237 _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8351__I _3750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7716_ _3526_ _3527_ _3528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8696_ _3704_ _4236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4928_ reg_file.reg_storage\[8\]\[22\] reg_file.reg_storage\[9\]\[22\] reg_file.reg_storage\[10\]\[22\]
+ reg_file.reg_storage\[11\]\[22\] _0757_ _0842_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_19_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7647_ _3437_ _3464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4859_ _0774_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7578_ _3388_ _3397_ _3398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9182__I _4510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9317_ _0103_ clknet_leaf_39_clk reg_file.reg_storage\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6529_ _2432_ _1835_ _2080_ _2433_ _2434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__7836__A2 _3638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9248_ _0034_ clknet_leaf_132_clk reg_file.reg_storage\[3\]\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9038__A1 _3995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9179_ _3963_ _4531_ _4534_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__I _4119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_82_clk clknet_4_12_0_clk clknet_leaf_82_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6024__A1 _1938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4586__A1 _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5138__I0 _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_55_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5838__A1 _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__I3 _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4964__I net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6263__A1 _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5900_ _1147_ _1815_ _1816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8372__S _4029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5449__S0 _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_93_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6880_ _2533_ _2513_ _2772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6015__A1 _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5831_ reg_file.reg_storage\[2\]\[9\] reg_file.reg_storage\[3\]\[9\] _1605_ _1747_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7763__A1 _2479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5762_ _1673_ _1675_ _1676_ _1677_ _1595_ _1596_ _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_8550_ reg_file.reg_storage\[12\]\[7\] _3940_ _4138_ _4139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_66_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7501_ _3317_ _3322_ _3327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4713_ net10 _0628_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8481_ reg_file.reg_storage\[13\]\[14\] _4088_ _4095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5693_ _1608_ _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ _0494_ net221 _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_44_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7432_ net77 _3263_ _3264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_141_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4575_ reg_file.reg_storage\[4\]\[0\] reg_file.reg_storage\[5\]\[0\] reg_file.reg_storage\[6\]\[0\]
+ reg_file.reg_storage\[7\]\[0\] _0497_ _0500_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_7363_ _3075_ _3200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_4_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9102_ _3969_ _4481_ _4487_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7294_ _3134_ _1829_ _3137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6314_ _2046_ _2224_ _2225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9033_ _3989_ _4406_ _4444_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6245_ _1903_ _0731_ _2157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5829__A1 _1734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8491__A2 _4094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6176_ _1110_ net203 _2089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_5127_ _1041_ _1042_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5058_ _0935_ _0972_ _0973_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input13_I inst[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_64_clk clknet_4_11_0_clk clknet_leaf_64_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8817_ _4309_ _4315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_48_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8748_ reg_file.reg_storage\[11\]\[7\] _4197_ _4272_ _4273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4663__S1 _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8679_ _4222_ _4214_ _4224_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6309__A2 _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6714__C1 _1636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8482__A2 _4094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6493__B2 _1586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8256__I _3921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8234__A2 _3924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_55_clk clknet_4_10_0_clk clknet_leaf_55_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_106_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7745__A1 net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4654__S1 _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6020__I1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6030_ _1800_ _1924_ _1944_ _1945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input5_I inst[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6787__A2 _2682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7981_ _3443_ _3765_ _3767_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xrebuffer26 _0498_ net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xrebuffer15 _0522_ net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_46_clk clknet_4_8_0_clk clknet_leaf_46_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6932_ _2585_ _2821_ _2822_ _2326_ _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_9651_ _0437_ clknet_leaf_78_clk reg_file.reg_storage\[4\]\[21\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6863_ _2360_ _2754_ _2755_ _2756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_49_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8602_ reg_file.reg_storage\[12\]\[30\] _4120_ _4168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7736__A1 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8830__S _4322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5814_ _0735_ _1729_ _1730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9582_ _0368_ clknet_leaf_66_clk reg_file.reg_storage\[9\]\[16\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6794_ _0797_ _0971_ _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5745_ reg_file.reg_storage\[12\]\[11\] reg_file.reg_storage\[13\]\[11\] reg_file.reg_storage\[14\]\[11\]
+ reg_file.reg_storage\[15\]\[11\] _0686_ _1588_ _1661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8533_ _4127_ _4128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5676_ reg_file.reg_storage\[1\]\[16\] _1591_ _1420_ _1592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8464_ _4073_ _4085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_44_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4869__I _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4627_ _0546_ _0548_ _0528_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7415_ _3208_ _3248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8395_ _4042_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5770__I0 reg_file.reg_storage\[1\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7346_ _3180_ _3184_ _3185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4558_ _0481_ _0483_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_130_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8277__S _3927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7277_ _3076_ _3121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9016_ _3966_ _4430_ _4434_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6228_ _2075_ _2136_ _2138_ _2140_ _2134_ _2141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__6475__A1 _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6159_ _1347_ _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4581__S0 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_142_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6778__A2 _2486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7975__A1 _3760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6242__A4 _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5833__S0 _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4961__A1 _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__I _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7750__I1 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4713__A1 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5108__I3 reg_file.reg_storage\[11\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6218__A1 _2046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6769__A2 _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7966__A1 _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_28_clk clknet_4_3_0_clk clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_47_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5824__S0 _1605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5530_ _1390_ _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_5_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8143__A1 _3424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5461_ _1084_ _1376_ _1377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8694__A2 _4181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7200_ _3050_ _3051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8180_ _3611_ _3888_ _3889_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5392_ _1307_ _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7131_ net134 _3002_ _3003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7062_ _2492_ _2526_ _2947_ _2582_ _2948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_1_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A1 _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6013_ _1071_ _1086_ _1927_ _1928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8825__S _4316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7964_ _3422_ _3751_ _3752_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_19_clk clknet_4_7_0_clk clknet_leaf_19_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8624__I _4179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__S1 _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ _2769_ _2786_ _2806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7895_ _3632_ _3691_ _3573_ _3692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_119_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6846_ _2724_ _2727_ _2739_ _2740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9634_ _0420_ clknet_leaf_18_clk reg_file.reg_storage\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_9565_ _0351_ clknet_leaf_105_clk reg_file.reg_storage\[10\]\[31\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6777_ _1620_ _1648_ _2626_ _2673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_8516_ _4007_ _4111_ _4114_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5728_ _1638_ _1640_ _1641_ _1643_ _1532_ _1535_ _1644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_91_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9496_ _0282_ clknet_leaf_106_clk reg_file.reg_storage\[8\]\[26\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input80_I pc[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8685__A2 _4223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8447_ _4073_ _4074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5659_ _1570_ _1572_ _1573_ _1574_ _1534_ _1537_ _1575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_21_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8378_ reg_file.reg_storage\[14\]\[5\] _3935_ _4029_ _4033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7329_ _3150_ _3162_ _3169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5120__A1 _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6319__I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7948__A1 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7948__B2 _3736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6620__A1 _2254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5893__I _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer6 _2400_ net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7613__I _3431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7636__B1 _3450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6439__A1 _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8645__S _4198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5133__I _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5111__A1 _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7939__A1 _3346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6611__A1 _2510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4961_ _0849_ _0851_ _0876_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8739__I0 reg_file.reg_storage\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7680_ net61 net38 net47 net56 _3433_ _3434_ _3494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_125_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6700_ _2573_ _2566_ _2599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4892_ reg_file.reg_storage\[1\]\[21\] _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6631_ _1838_ _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_22_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5568__I3 reg_file.reg_storage\[7\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5273__S1 _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9350_ _0136_ clknet_leaf_44_clk reg_file.reg_storage\[7\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8301_ _3973_ _3974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8116__A1 reg_file.reg_storage\[2\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6562_ _2180_ _2463_ _2465_ _2257_ _2466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_42_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5513_ _1428_ _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_89_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9281_ _0067_ clknet_4_5_0_clk reg_file.reg_storage\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6493_ _1735_ _1743_ _1829_ _1586_ _1752_ _2399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_140_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5444_ _1359_ _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_76_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8232_ _3922_ _3923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_8_clk clknet_4_6_0_clk clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8163_ reg_file.reg_storage\[6\]\[7\] _3511_ _3879_ _3880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8419__A2 _4024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8619__I _4181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7114_ _2987_ _2992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5375_ net91 _0888_ _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9092__A2 _4475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8094_ _3836_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5102__A1 _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7045_ _2905_ _2908_ _2931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8996_ _4423_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_70_clk_I clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7947_ _3715_ _3366_ _3737_ _3738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7878_ _2967_ _3641_ _3642_ net46 _3677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_65_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8355__A1 _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9617_ _0403_ clknet_leaf_71_clk reg_file.reg_storage\[1\]\[19\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6829_ _1852_ _2722_ _2723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_65_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9185__I _4516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4916__A1 _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6905__A2 _1881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9548_ _0334_ clknet_leaf_65_clk reg_file.reg_storage\[10\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_85_clk_I clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9479_ _0265_ clknet_leaf_27_clk reg_file.reg_storage\[8\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_129_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8465__S _4085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_23_clk_I clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8264__I _3921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8594__A1 _3996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_38_clk_I clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7608__I _3426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5329__S _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5255__S1 _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8897__A2 _4363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8649__A2 _4203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5007__S1 _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6668__B _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7321__A2 _3161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5160_ reg_file.reg_storage\[1\]\[26\] _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__9074__A2 _4462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5091_ _1000_ _1004_ _1005_ _1006_ _0786_ _0788_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_71_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8850_ reg_file.reg_storage\[10\]\[16\] _4325_ _4334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8781_ _4230_ _4288_ _4291_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5993_ _1862_ _0910_ _1908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7801_ _3572_ _3607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_87_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7732_ _3542_ _3543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _0756_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6623__S _2052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8337__A1 reg_file.reg_storage\[7\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_9402_ _0188_ clknet_leaf_96_clk reg_file.reg_storage\[14\]\[28\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4875_ _0751_ _0790_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7663_ reg_file.reg_storage\[5\]\[4\] _3444_ _3479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7594_ _0595_ _3414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_131_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6614_ _1817_ _2442_ _2515_ _2482_ _2516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_46_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5038__I _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_104_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_9333_ _0119_ clknet_leaf_23_clk reg_file.reg_storage\[6\]\[23\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6545_ _2391_ _2445_ _2449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_6_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9264_ _0050_ clknet_leaf_46_clk reg_file.reg_storage\[3\]\[18\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer16_I _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8215_ reg_file.reg_storage\[6\]\[30\] _3861_ _3909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7312__A2 _2413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _2121_ _2336_ _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9195_ _3986_ _4513_ _4543_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_7_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5427_ _0745_ _1112_ _1113_ _1342_ _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_input43_I mem_ld_dat[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8146_ _3868_ _3869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5358_ reg_file.reg_storage\[1\]\[5\] _1273_ _1271_ _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5874__A2 _1789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8285__S _3927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8077_ reg_file.reg_storage\[2\]\[6\] _3819_ _3827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7076__A1 _2103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5477__I2 reg_file.reg_storage\[14\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7028_ _2906_ _2912_ _2174_ _2914_ _2915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5289_ _1195_ _1204_ _0970_ _1205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_EDGE_ROW_113_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8084__I _3816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8979_ _3918_ _4411_ _4413_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8812__I _4310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5149__S _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7000__A1 _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7428__I net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_122_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5562__A1 _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7551__A2 _3360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4787__I _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6488__B _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8259__I _3529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__A2 _1780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_131_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7606__A3 _3394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6814__A1 _2038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__S0 _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8923__S _4365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6042__A2 _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8319__A1 reg_file.reg_storage\[7\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_140_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4660_ reg_file.reg_storage\[8\]\[7\] reg_file.reg_storage\[9\]\[7\] reg_file.reg_storage\[10\]\[7\]
+ reg_file.reg_storage\[11\]\[7\] _0577_ _0578_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_44_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5228__S1 _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7542__A2 _3356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _1281_ _2239_ _2240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4591_ reg_file.reg_storage\[2\]\[1\] reg_file.reg_storage\[3\]\[1\] _0502_ _0516_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6261_ _1344_ _1346_ _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__9047__A2 _4407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8000_ reg_file.reg_storage\[3\]\[9\] _3778_ _3779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5212_ reg_file.reg_storage\[8\]\[12\] reg_file.reg_storage\[9\]\[12\] reg_file.reg_storage\[10\]\[12\]
+ reg_file.reg_storage\[11\]\[12\] _1122_ _1123_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6192_ _2104_ _2105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5143_ _1057_ _1058_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_43_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5164__S0 _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5074_ _0779_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_79_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8902_ _4367_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8833_ _4324_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_84_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6033__A2 _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8764_ reg_file.reg_storage\[11\]\[14\] _4275_ _4282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5976_ _1010_ _1508_ _1891_ _1892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4927_ reg_file.reg_storage\[12\]\[22\] reg_file.reg_storage\[13\]\[22\] reg_file.reg_storage\[14\]\[22\]
+ reg_file.reg_storage\[15\]\[22\] _0757_ _0842_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_63_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8695_ _4234_ _4183_ _4235_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7715_ _3485_ _3123_ _3496_ _3128_ _3486_ _3527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_19_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7646_ _3414_ _3462_ _3463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_117_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4858_ _0763_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_62_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7533__A2 _3356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4789_ net4 _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__4978__S0 _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7577_ _3389_ _3396_ _3397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_9316_ _0102_ clknet_leaf_17_clk reg_file.reg_storage\[6\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4601__S _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6528_ _2432_ _1835_ _2076_ _2433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8079__I _3816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9247_ _0033_ clknet_leaf_19_clk reg_file.reg_storage\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6459_ _2035_ _2364_ _2365_ _2366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9178_ reg_file.reg_storage\[15\]\[16\] _4525_ _4534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8129_ _3734_ _3854_ _3856_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_126_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8743__S _4266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4980__I _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7212__A1 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5449__S1 _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ reg_file.reg_storage\[8\]\[9\] reg_file.reg_storage\[9\]\[9\] reg_file.reg_storage\[10\]\[9\]
+ reg_file.reg_storage\[11\]\[9\] _1590_ _1642_ _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_76_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5761_ reg_file.reg_storage\[4\]\[10\] reg_file.reg_storage\[5\]\[10\] reg_file.reg_storage\[6\]\[10\]
+ reg_file.reg_storage\[7\]\[10\] _1358_ _1657_ _1677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_56_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5774__A1 _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8480_ _4074_ _4094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7500_ net83 _3326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4712_ _0627_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_126_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7431_ _1557_ _3263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5692_ _0518_ _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_142_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5526__A1 _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4643_ _0558_ _0560_ _0561_ _0562_ _0542_ _0563_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_114_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4574_ _0499_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7362_ _3179_ _3194_ _3199_ net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9101_ reg_file.reg_storage\[4\]\[18\] _4486_ _4487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7293_ _3133_ _3135_ _3136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_12_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6313_ _1978_ _2223_ _2198_ _2224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9032_ reg_file.reg_storage\[1\]\[24\] _4443_ _4444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6244_ _2153_ _2155_ _1766_ _2156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_0_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6175_ _1239_ _0884_ _0793_ _0729_ _0725_ _0713_ _2088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XANTENNA__5137__S0 _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5126_ _0795_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5057_ _0884_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8563__S _4131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7203__A1 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8816_ _4177_ _4312_ _4314_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8747_ _4260_ _4272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5959_ _1873_ _1031_ _1040_ _1874_ _1875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_36_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8678_ reg_file.reg_storage\[8\]\[18\] _4223_ _4224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7629_ net51 _3447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__7706__I _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7690__A1 _3428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7993__A2 _3765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7745__A2 _3504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7681__A1 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8447__I _4073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6484__A2 _1832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8383__S _4035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4590__S1 _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer16 _1439_ net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7980_ reg_file.reg_storage\[3\]\[1\] _3766_ _3767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xrebuffer27 _0610_ net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6931_ _2137_ _2607_ _2822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5995__A1 _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9650_ _0436_ clknet_leaf_79_clk reg_file.reg_storage\[4\]\[20\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6862_ _2217_ _2658_ _2755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8601_ _4007_ _4164_ _4167_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5813_ _1604_ _1728_ _1729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_9581_ _0367_ clknet_leaf_14_clk reg_file.reg_storage\[9\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8532_ _4126_ _4127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6793_ _2289_ _2470_ _2689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6795__I0 _2636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5744_ reg_file.reg_storage\[1\]\[11\] _1659_ _1657_ _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ reg_file.reg_storage\[2\]\[16\] reg_file.reg_storage\[3\]\[16\] _1590_ _1591_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8463_ _3938_ _4075_ _4084_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8161__A2 _3869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8394_ reg_file.reg_storage\[14\]\[12\] _3953_ _4028_ _4042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4626_ reg_file.reg_storage\[1\]\[4\] _0547_ _0499_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7414_ _3200_ _3237_ _3246_ _3046_ _3247_ net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_103_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7345_ _3183_ _3184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4557_ _0482_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_92_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7276_ _3077_ _3115_ _3120_ net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9015_ reg_file.reg_storage\[1\]\[17\] _4424_ _4434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8357__I _4016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4885__I _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6227_ _2139_ _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6158_ _2069_ _2071_ _2072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ _0824_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4581__S1 _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5710__S _1623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6089_ _1241_ _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output112_I net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5738__A1 _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5589__I1 _1502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_101_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5833__S1 _1623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4961__A2 _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5210__I0 reg_file.reg_storage\[1\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4713__A2 _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8267__I _3555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4744__B _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5824__S1 _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8730__I _4260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6451__S _2137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8143__A2 _3865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5460_ _1351_ _1356_ _1375_ _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5588__S0 _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8378__S _4029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _1302_ _1304_ _1305_ _1306_ _0914_ net9 _1307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7130_ _3001_ _3002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7061_ _2046_ _2945_ _2946_ _1999_ _2947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6012_ _1084_ _1058_ _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
.ends

