VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tinyrv
  CLASS BLOCK ;
  FOREIGN tinyrv ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 600.000 ;
  PIN alu_out_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 282.240 500.000 282.800 ;
    END
  END alu_out_out[0]
  PIN alu_out_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 596.000 413.840 600.000 ;
    END
  END alu_out_out[10]
  PIN alu_out_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 596.000 427.280 600.000 ;
    END
  END alu_out_out[11]
  PIN alu_out_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 596.000 444.080 600.000 ;
    END
  END alu_out_out[12]
  PIN alu_out_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 596.000 450.800 600.000 ;
    END
  END alu_out_out[13]
  PIN alu_out_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 596.000 440.720 600.000 ;
    END
  END alu_out_out[14]
  PIN alu_out_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 596.000 360.080 600.000 ;
    END
  END alu_out_out[15]
  PIN alu_out_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 329.280 500.000 329.840 ;
    END
  END alu_out_out[16]
  PIN alu_out_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 252.000 500.000 252.560 ;
    END
  END alu_out_out[17]
  PIN alu_out_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 245.280 500.000 245.840 ;
    END
  END alu_out_out[18]
  PIN alu_out_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 215.040 500.000 215.600 ;
    END
  END alu_out_out[19]
  PIN alu_out_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 366.240 500.000 366.800 ;
    END
  END alu_out_out[1]
  PIN alu_out_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 198.240 500.000 198.800 ;
    END
  END alu_out_out[20]
  PIN alu_out_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 178.080 500.000 178.640 ;
    END
  END alu_out_out[21]
  PIN alu_out_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 0.000 360.080 4.000 ;
    END
  END alu_out_out[22]
  PIN alu_out_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 0.000 363.440 4.000 ;
    END
  END alu_out_out[23]
  PIN alu_out_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 0.000 376.880 4.000 ;
    END
  END alu_out_out[24]
  PIN alu_out_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 0.000 417.200 4.000 ;
    END
  END alu_out_out[25]
  PIN alu_out_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 0.000 403.760 4.000 ;
    END
  END alu_out_out[26]
  PIN alu_out_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 0.000 410.480 4.000 ;
    END
  END alu_out_out[27]
  PIN alu_out_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 0.000 413.840 4.000 ;
    END
  END alu_out_out[28]
  PIN alu_out_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 0.000 400.400 4.000 ;
    END
  END alu_out_out[29]
  PIN alu_out_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 376.320 500.000 376.880 ;
    END
  END alu_out_out[2]
  PIN alu_out_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 0.000 407.120 4.000 ;
    END
  END alu_out_out[30]
  PIN alu_out_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 0.000 373.520 4.000 ;
    END
  END alu_out_out[31]
  PIN alu_out_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 399.840 500.000 400.400 ;
    END
  END alu_out_out[3]
  PIN alu_out_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 596.000 373.520 600.000 ;
    END
  END alu_out_out[4]
  PIN alu_out_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 596.000 363.440 600.000 ;
    END
  END alu_out_out[5]
  PIN alu_out_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 596.000 386.960 600.000 ;
    END
  END alu_out_out[6]
  PIN alu_out_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 596.000 383.600 600.000 ;
    END
  END alu_out_out[7]
  PIN alu_out_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 596.000 423.920 600.000 ;
    END
  END alu_out_out[8]
  PIN alu_out_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 596.000 390.320 600.000 ;
    END
  END alu_out_out[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.560 4.000 575.120 ;
    END
  END clk
  PIN inst_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 262.080 500.000 262.640 ;
    END
  END inst_in[0]
  PIN inst_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 312.480 4.000 313.040 ;
    END
  END inst_in[10]
  PIN inst_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 309.120 500.000 309.680 ;
    END
  END inst_in[11]
  PIN inst_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 285.600 500.000 286.160 ;
    END
  END inst_in[12]
  PIN inst_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 295.680 500.000 296.240 ;
    END
  END inst_in[13]
  PIN inst_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 299.040 500.000 299.600 ;
    END
  END inst_in[14]
  PIN inst_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.080 4.000 262.640 ;
    END
  END inst_in[15]
  PIN inst_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 255.360 4.000 255.920 ;
    END
  END inst_in[16]
  PIN inst_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 0.000 229.040 4.000 ;
    END
  END inst_in[17]
  PIN inst_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 218.400 500.000 218.960 ;
    END
  END inst_in[18]
  PIN inst_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 235.200 500.000 235.760 ;
    END
  END inst_in[19]
  PIN inst_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 265.440 500.000 266.000 ;
    END
  END inst_in[1]
  PIN inst_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.400 4.000 386.960 ;
    END
  END inst_in[20]
  PIN inst_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 359.520 4.000 360.080 ;
    END
  END inst_in[21]
  PIN inst_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 349.440 4.000 350.000 ;
    END
  END inst_in[22]
  PIN inst_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 336.000 4.000 336.560 ;
    END
  END inst_in[23]
  PIN inst_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 315.840 500.000 316.400 ;
    END
  END inst_in[24]
  PIN inst_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 332.640 500.000 333.200 ;
    END
  END inst_in[25]
  PIN inst_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 336.000 500.000 336.560 ;
    END
  END inst_in[26]
  PIN inst_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 386.400 500.000 386.960 ;
    END
  END inst_in[27]
  PIN inst_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 339.360 500.000 339.920 ;
    END
  END inst_in[28]
  PIN inst_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 342.720 500.000 343.280 ;
    END
  END inst_in[29]
  PIN inst_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 272.160 500.000 272.720 ;
    END
  END inst_in[2]
  PIN inst_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 278.880 500.000 279.440 ;
    END
  END inst_in[30]
  PIN inst_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 201.600 500.000 202.160 ;
    END
  END inst_in[31]
  PIN inst_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 268.800 500.000 269.360 ;
    END
  END inst_in[3]
  PIN inst_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 275.520 500.000 276.080 ;
    END
  END inst_in[4]
  PIN inst_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 288.960 500.000 289.520 ;
    END
  END inst_in[5]
  PIN inst_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 292.320 500.000 292.880 ;
    END
  END inst_in[6]
  PIN inst_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.880 4.000 279.440 ;
    END
  END inst_in[7]
  PIN inst_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 309.120 4.000 309.680 ;
    END
  END inst_in[8]
  PIN inst_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 295.680 4.000 296.240 ;
    END
  END inst_in[9]
  PIN mem_load_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 349.440 500.000 350.000 ;
    END
  END mem_load_out[0]
  PIN mem_load_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 596.000 376.880 600.000 ;
    END
  END mem_load_out[10]
  PIN mem_load_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 596.000 380.240 600.000 ;
    END
  END mem_load_out[11]
  PIN mem_load_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 596.000 370.160 600.000 ;
    END
  END mem_load_out[12]
  PIN mem_load_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 596.000 366.800 600.000 ;
    END
  END mem_load_out[13]
  PIN mem_load_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 596.000 356.720 600.000 ;
    END
  END mem_load_out[14]
  PIN mem_load_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 596.000 353.360 600.000 ;
    END
  END mem_load_out[15]
  PIN mem_load_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 302.400 500.000 302.960 ;
    END
  END mem_load_out[16]
  PIN mem_load_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 305.760 500.000 306.320 ;
    END
  END mem_load_out[17]
  PIN mem_load_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 231.840 500.000 232.400 ;
    END
  END mem_load_out[18]
  PIN mem_load_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 228.480 500.000 229.040 ;
    END
  END mem_load_out[19]
  PIN mem_load_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 362.880 500.000 363.440 ;
    END
  END mem_load_out[1]
  PIN mem_load_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 194.880 500.000 195.440 ;
    END
  END mem_load_out[20]
  PIN mem_load_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 0.000 350.000 4.000 ;
    END
  END mem_load_out[21]
  PIN mem_load_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 0.000 356.720 4.000 ;
    END
  END mem_load_out[22]
  PIN mem_load_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 0.000 353.360 4.000 ;
    END
  END mem_load_out[23]
  PIN mem_load_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 0.000 366.800 4.000 ;
    END
  END mem_load_out[24]
  PIN mem_load_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 0.000 370.160 4.000 ;
    END
  END mem_load_out[25]
  PIN mem_load_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 0.000 380.240 4.000 ;
    END
  END mem_load_out[26]
  PIN mem_load_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 0.000 383.600 4.000 ;
    END
  END mem_load_out[27]
  PIN mem_load_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 0.000 397.040 4.000 ;
    END
  END mem_load_out[28]
  PIN mem_load_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 0.000 393.680 4.000 ;
    END
  END mem_load_out[29]
  PIN mem_load_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 379.680 500.000 380.240 ;
    END
  END mem_load_out[2]
  PIN mem_load_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 0.000 386.960 4.000 ;
    END
  END mem_load_out[30]
  PIN mem_load_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 0.000 390.320 4.000 ;
    END
  END mem_load_out[31]
  PIN mem_load_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 393.120 500.000 393.680 ;
    END
  END mem_load_out[3]
  PIN mem_load_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 596.000 336.560 600.000 ;
    END
  END mem_load_out[4]
  PIN mem_load_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 596.000 350.000 600.000 ;
    END
  END mem_load_out[5]
  PIN mem_load_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 596.000 343.280 600.000 ;
    END
  END mem_load_out[6]
  PIN mem_load_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 413.280 500.000 413.840 ;
    END
  END mem_load_out[7]
  PIN mem_load_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 596.000 346.640 600.000 ;
    END
  END mem_load_out[8]
  PIN mem_load_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 596.000 339.920 600.000 ;
    END
  END mem_load_out[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 492.800 585.610 ;
      LAYER Metal2 ;
        RECT 0.140 595.700 335.700 596.000 ;
        RECT 336.860 595.700 339.060 596.000 ;
        RECT 340.220 595.700 342.420 596.000 ;
        RECT 343.580 595.700 345.780 596.000 ;
        RECT 346.940 595.700 349.140 596.000 ;
        RECT 350.300 595.700 352.500 596.000 ;
        RECT 353.660 595.700 355.860 596.000 ;
        RECT 357.020 595.700 359.220 596.000 ;
        RECT 360.380 595.700 362.580 596.000 ;
        RECT 363.740 595.700 365.940 596.000 ;
        RECT 367.100 595.700 369.300 596.000 ;
        RECT 370.460 595.700 372.660 596.000 ;
        RECT 373.820 595.700 376.020 596.000 ;
        RECT 377.180 595.700 379.380 596.000 ;
        RECT 380.540 595.700 382.740 596.000 ;
        RECT 383.900 595.700 386.100 596.000 ;
        RECT 387.260 595.700 389.460 596.000 ;
        RECT 390.620 595.700 412.980 596.000 ;
        RECT 414.140 595.700 423.060 596.000 ;
        RECT 424.220 595.700 426.420 596.000 ;
        RECT 427.580 595.700 439.860 596.000 ;
        RECT 441.020 595.700 443.220 596.000 ;
        RECT 444.380 595.700 449.940 596.000 ;
        RECT 451.100 595.700 497.700 596.000 ;
        RECT 0.140 4.300 497.700 595.700 ;
        RECT 0.140 4.000 228.180 4.300 ;
        RECT 229.340 4.000 349.140 4.300 ;
        RECT 350.300 4.000 352.500 4.300 ;
        RECT 353.660 4.000 355.860 4.300 ;
        RECT 357.020 4.000 359.220 4.300 ;
        RECT 360.380 4.000 362.580 4.300 ;
        RECT 363.740 4.000 365.940 4.300 ;
        RECT 367.100 4.000 369.300 4.300 ;
        RECT 370.460 4.000 372.660 4.300 ;
        RECT 373.820 4.000 376.020 4.300 ;
        RECT 377.180 4.000 379.380 4.300 ;
        RECT 380.540 4.000 382.740 4.300 ;
        RECT 383.900 4.000 386.100 4.300 ;
        RECT 387.260 4.000 389.460 4.300 ;
        RECT 390.620 4.000 392.820 4.300 ;
        RECT 393.980 4.000 396.180 4.300 ;
        RECT 397.340 4.000 399.540 4.300 ;
        RECT 400.700 4.000 402.900 4.300 ;
        RECT 404.060 4.000 406.260 4.300 ;
        RECT 407.420 4.000 409.620 4.300 ;
        RECT 410.780 4.000 412.980 4.300 ;
        RECT 414.140 4.000 416.340 4.300 ;
        RECT 417.500 4.000 497.700 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 575.420 497.750 587.860 ;
        RECT 4.300 574.260 497.750 575.420 ;
        RECT 0.090 414.140 497.750 574.260 ;
        RECT 0.090 412.980 495.700 414.140 ;
        RECT 0.090 400.700 497.750 412.980 ;
        RECT 0.090 399.540 495.700 400.700 ;
        RECT 0.090 393.980 497.750 399.540 ;
        RECT 0.090 392.820 495.700 393.980 ;
        RECT 0.090 387.260 497.750 392.820 ;
        RECT 4.300 386.100 495.700 387.260 ;
        RECT 0.090 380.540 497.750 386.100 ;
        RECT 0.090 379.380 495.700 380.540 ;
        RECT 0.090 377.180 497.750 379.380 ;
        RECT 0.090 376.020 495.700 377.180 ;
        RECT 0.090 367.100 497.750 376.020 ;
        RECT 0.090 365.940 495.700 367.100 ;
        RECT 0.090 363.740 497.750 365.940 ;
        RECT 0.090 362.580 495.700 363.740 ;
        RECT 0.090 360.380 497.750 362.580 ;
        RECT 4.300 359.220 497.750 360.380 ;
        RECT 0.090 350.300 497.750 359.220 ;
        RECT 4.300 349.140 495.700 350.300 ;
        RECT 0.090 343.580 497.750 349.140 ;
        RECT 0.090 342.420 495.700 343.580 ;
        RECT 0.090 340.220 497.750 342.420 ;
        RECT 0.090 339.060 495.700 340.220 ;
        RECT 0.090 336.860 497.750 339.060 ;
        RECT 4.300 335.700 495.700 336.860 ;
        RECT 0.090 333.500 497.750 335.700 ;
        RECT 0.090 332.340 495.700 333.500 ;
        RECT 0.090 330.140 497.750 332.340 ;
        RECT 0.090 328.980 495.700 330.140 ;
        RECT 0.090 316.700 497.750 328.980 ;
        RECT 0.090 315.540 495.700 316.700 ;
        RECT 0.090 313.340 497.750 315.540 ;
        RECT 4.300 312.180 497.750 313.340 ;
        RECT 0.090 309.980 497.750 312.180 ;
        RECT 4.300 308.820 495.700 309.980 ;
        RECT 0.090 306.620 497.750 308.820 ;
        RECT 0.090 305.460 495.700 306.620 ;
        RECT 0.090 303.260 497.750 305.460 ;
        RECT 0.090 302.100 495.700 303.260 ;
        RECT 0.090 299.900 497.750 302.100 ;
        RECT 0.090 298.740 495.700 299.900 ;
        RECT 0.090 296.540 497.750 298.740 ;
        RECT 4.300 295.380 495.700 296.540 ;
        RECT 0.090 293.180 497.750 295.380 ;
        RECT 0.090 292.020 495.700 293.180 ;
        RECT 0.090 289.820 497.750 292.020 ;
        RECT 0.090 288.660 495.700 289.820 ;
        RECT 0.090 286.460 497.750 288.660 ;
        RECT 0.090 285.300 495.700 286.460 ;
        RECT 0.090 283.100 497.750 285.300 ;
        RECT 0.090 281.940 495.700 283.100 ;
        RECT 0.090 279.740 497.750 281.940 ;
        RECT 4.300 278.580 495.700 279.740 ;
        RECT 0.090 276.380 497.750 278.580 ;
        RECT 0.090 275.220 495.700 276.380 ;
        RECT 0.090 273.020 497.750 275.220 ;
        RECT 0.090 271.860 495.700 273.020 ;
        RECT 0.090 269.660 497.750 271.860 ;
        RECT 0.090 268.500 495.700 269.660 ;
        RECT 0.090 266.300 497.750 268.500 ;
        RECT 0.090 265.140 495.700 266.300 ;
        RECT 0.090 262.940 497.750 265.140 ;
        RECT 4.300 261.780 495.700 262.940 ;
        RECT 0.090 256.220 497.750 261.780 ;
        RECT 4.300 255.060 497.750 256.220 ;
        RECT 0.090 252.860 497.750 255.060 ;
        RECT 0.090 251.700 495.700 252.860 ;
        RECT 0.090 246.140 497.750 251.700 ;
        RECT 0.090 244.980 495.700 246.140 ;
        RECT 0.090 236.060 497.750 244.980 ;
        RECT 0.090 234.900 495.700 236.060 ;
        RECT 0.090 232.700 497.750 234.900 ;
        RECT 0.090 231.540 495.700 232.700 ;
        RECT 0.090 229.340 497.750 231.540 ;
        RECT 0.090 228.180 495.700 229.340 ;
        RECT 0.090 219.260 497.750 228.180 ;
        RECT 0.090 218.100 495.700 219.260 ;
        RECT 0.090 215.900 497.750 218.100 ;
        RECT 0.090 214.740 495.700 215.900 ;
        RECT 0.090 202.460 497.750 214.740 ;
        RECT 0.090 201.300 495.700 202.460 ;
        RECT 0.090 199.100 497.750 201.300 ;
        RECT 0.090 197.940 495.700 199.100 ;
        RECT 0.090 195.740 497.750 197.940 ;
        RECT 0.090 194.580 495.700 195.740 ;
        RECT 0.090 178.940 497.750 194.580 ;
        RECT 0.090 177.780 495.700 178.940 ;
        RECT 0.090 10.220 497.750 177.780 ;
      LAYER Metal4 ;
        RECT 20.860 16.890 21.940 582.310 ;
        RECT 24.140 16.890 98.740 582.310 ;
        RECT 100.940 16.890 175.540 582.310 ;
        RECT 177.740 16.890 252.340 582.310 ;
        RECT 254.540 16.890 329.140 582.310 ;
        RECT 331.340 16.890 405.940 582.310 ;
        RECT 408.140 16.890 482.740 582.310 ;
        RECT 484.940 16.890 493.220 582.310 ;
  END
END tinyrv
END LIBRARY

