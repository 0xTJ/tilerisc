magic
tech gf180mcuD
magscale 1 10
timestamp 1700139236
<< metal2 >>
rect 3744 48104 3856 48776
rect 3724 47976 3856 48104
rect 4444 48104 4556 48776
rect 5344 48104 5456 48776
rect 4444 47976 4564 48104
rect 5344 47976 5460 48104
rect 13444 47976 13556 48776
rect 14144 48104 14256 48776
rect 14140 47976 14256 48104
rect 14544 47976 14656 48776
rect 14994 47976 15106 48776
rect 15444 47976 15556 48776
rect 16044 47976 16156 48776
rect 24244 48104 24356 48776
rect 24220 47976 24356 48104
rect 25044 48104 25156 48776
rect 25044 47976 25172 48104
rect 25744 47976 25856 48776
rect 30944 48104 31056 48776
rect 30940 47976 31056 48104
rect 31944 47976 32056 48776
rect 32744 48104 32856 48776
rect 32732 47976 32856 48104
rect 36844 47976 36956 48776
rect 46568 47976 46680 48776
rect 52944 48104 53056 48776
rect 52944 47976 53060 48104
rect 54644 47976 54756 48776
rect 56344 47976 56456 48776
rect 59244 47976 59356 48776
rect 63344 48104 63456 48776
rect 63344 47976 63476 48104
rect 63744 47976 63856 48776
rect 64944 47976 65056 48776
rect 73044 47976 73156 48776
rect 73744 48104 73856 48776
rect 73724 47976 73856 48104
rect 74144 47976 74256 48776
rect 74544 48104 74656 48776
rect 74544 47976 74676 48104
rect 74944 47976 75056 48776
rect 75644 48104 75756 48776
rect 75628 47976 75756 48104
rect 83844 48104 83956 48776
rect 83844 47976 83972 48104
rect 84644 47976 84756 48776
rect 85344 47976 85456 48776
rect 3724 47796 3780 47976
rect 3724 47740 3836 47796
rect 3780 47544 3836 47740
rect 4508 47544 4564 47976
rect 5404 47544 5460 47976
rect 13468 47544 13524 47976
rect 14140 47544 14196 47976
rect 14588 47544 14644 47976
rect 15036 47544 15092 47976
rect 15484 47544 15540 47976
rect 16044 47544 16100 47976
rect 24220 47544 24276 47976
rect 25116 47544 25172 47976
rect 25788 47544 25844 47976
rect 30940 47544 30996 47976
rect 31948 47796 32004 47976
rect 31948 47740 32060 47796
rect 32004 47544 32060 47740
rect 32732 47544 32788 47976
rect 36876 47544 36932 47976
rect 46620 47544 46676 47976
rect 53004 47544 53060 47976
rect 54684 47544 54740 47976
rect 56364 47544 56420 47976
rect 59276 47544 59332 47976
rect 63420 47544 63476 47976
rect 63756 47544 63812 47976
rect 64988 47544 65044 47976
rect 73052 47544 73108 47976
rect 73724 47544 73780 47976
rect 74172 47544 74228 47976
rect 74620 47544 74676 47976
rect 74956 47544 75012 47976
rect 75628 47544 75684 47976
rect 83916 47544 83972 47976
rect 84700 47544 84756 47976
rect 85372 47544 85428 47976
<< metal3 >>
rect 1106 45436 1582 45472
rect 1106 45380 1130 45436
rect 1186 45380 1254 45436
rect 1310 45380 1378 45436
rect 1434 45380 1502 45436
rect 1558 45380 1582 45436
rect 1106 45344 1582 45380
rect 85788 45436 86264 45472
rect 85788 45380 85812 45436
rect 85868 45380 85936 45436
rect 85992 45380 86060 45436
rect 86116 45380 86184 45436
rect 86240 45380 86264 45436
rect 85788 45344 86264 45380
rect 1844 45025 2014 45074
rect 1844 44969 1901 45025
rect 1957 44969 2014 45025
rect 1844 44901 2014 44969
rect 1844 44845 1901 44901
rect 1957 44845 2014 44901
rect 1844 44777 2014 44845
rect 1844 44721 1901 44777
rect 1957 44721 2014 44777
rect 1844 44653 2014 44721
rect 1844 44597 1901 44653
rect 1957 44597 2014 44653
rect 1844 44529 2014 44597
rect 1844 44473 1901 44529
rect 1957 44473 2014 44529
rect 1844 44405 2014 44473
rect 1844 44349 1901 44405
rect 1957 44349 2014 44405
rect 1844 44281 2014 44349
rect 1844 44225 1901 44281
rect 1957 44225 2014 44281
rect 1844 44157 2014 44225
rect 1844 44101 1901 44157
rect 1957 44101 2014 44157
rect 1844 44033 2014 44101
rect 1844 43977 1901 44033
rect 1957 43977 2014 44033
rect 1844 43909 2014 43977
rect 1844 43853 1901 43909
rect 1957 43853 2014 43909
rect 1844 43804 2014 43853
rect 86526 45025 86630 45074
rect 86526 44969 86550 45025
rect 86606 44969 86630 45025
rect 86526 44901 86630 44969
rect 86526 44845 86550 44901
rect 86606 44845 86630 44901
rect 86526 44777 86630 44845
rect 86526 44721 86550 44777
rect 86606 44721 86630 44777
rect 86526 44653 86630 44721
rect 86526 44597 86550 44653
rect 86606 44597 86630 44653
rect 86526 44529 86630 44597
rect 86526 44473 86550 44529
rect 86606 44473 86630 44529
rect 86526 44405 86630 44473
rect 86526 44349 86550 44405
rect 86606 44349 86630 44405
rect 86526 44281 86630 44349
rect 86526 44225 86550 44281
rect 86606 44225 86630 44281
rect 86526 44157 86630 44225
rect 86526 44101 86550 44157
rect 86606 44101 86630 44157
rect 86526 44033 86630 44101
rect 86526 43977 86550 44033
rect 86606 43977 86630 44033
rect 86526 43909 86630 43977
rect 86526 43853 86550 43909
rect 86606 43853 86630 43909
rect 86526 43804 86630 43853
rect 86650 45025 87126 45074
rect 86650 44969 86674 45025
rect 86730 44969 86798 45025
rect 86854 44969 86922 45025
rect 86978 44969 87046 45025
rect 87102 44969 87126 45025
rect 86650 44901 87126 44969
rect 86650 44845 86674 44901
rect 86730 44845 86798 44901
rect 86854 44845 86922 44901
rect 86978 44845 87046 44901
rect 87102 44845 87126 44901
rect 86650 44777 87126 44845
rect 86650 44721 86674 44777
rect 86730 44721 86798 44777
rect 86854 44721 86922 44777
rect 86978 44721 87046 44777
rect 87102 44721 87126 44777
rect 86650 44653 87126 44721
rect 86650 44597 86674 44653
rect 86730 44597 86798 44653
rect 86854 44597 86922 44653
rect 86978 44597 87046 44653
rect 87102 44597 87126 44653
rect 86650 44529 87126 44597
rect 86650 44473 86674 44529
rect 86730 44473 86798 44529
rect 86854 44473 86922 44529
rect 86978 44473 87046 44529
rect 87102 44473 87126 44529
rect 86650 44405 87126 44473
rect 86650 44349 86674 44405
rect 86730 44349 86798 44405
rect 86854 44349 86922 44405
rect 86978 44349 87046 44405
rect 87102 44349 87126 44405
rect 86650 44281 87126 44349
rect 86650 44225 86674 44281
rect 86730 44225 86798 44281
rect 86854 44225 86922 44281
rect 86978 44225 87046 44281
rect 87102 44225 87126 44281
rect 86650 44157 87126 44225
rect 86650 44101 86674 44157
rect 86730 44101 86798 44157
rect 86854 44101 86922 44157
rect 86978 44101 87046 44157
rect 87102 44101 87126 44157
rect 86650 44033 87126 44101
rect 86650 43977 86674 44033
rect 86730 43977 86798 44033
rect 86854 43977 86922 44033
rect 86978 43977 87046 44033
rect 87102 43977 87126 44033
rect 86650 43909 87126 43977
rect 86650 43853 86674 43909
rect 86730 43853 86798 43909
rect 86854 43853 86922 43909
rect 86978 43853 87046 43909
rect 87102 43853 87126 43909
rect 86650 43804 87126 43853
rect 86526 41791 86630 41810
rect 86526 41735 86550 41791
rect 86606 41735 86630 41791
rect 86526 41667 86630 41735
rect 86526 41611 86550 41667
rect 86606 41611 86630 41667
rect 86526 41543 86630 41611
rect 86526 41487 86550 41543
rect 86606 41487 86630 41543
rect 86526 41419 86630 41487
rect 86526 41363 86550 41419
rect 86606 41363 86630 41419
rect 86526 41344 86630 41363
rect 86650 41791 87126 41810
rect 86650 41735 86674 41791
rect 86730 41735 86798 41791
rect 86854 41735 86922 41791
rect 86978 41735 87046 41791
rect 87102 41735 87126 41791
rect 86650 41667 87126 41735
rect 86650 41611 86674 41667
rect 86730 41611 86798 41667
rect 86854 41611 86922 41667
rect 86978 41611 87046 41667
rect 87102 41611 87126 41667
rect 86650 41543 87126 41611
rect 86650 41487 86674 41543
rect 86730 41487 86798 41543
rect 86854 41487 86922 41543
rect 86978 41487 87046 41543
rect 87102 41487 87126 41543
rect 86650 41419 87126 41487
rect 86650 41363 86674 41419
rect 86730 41363 86798 41419
rect 86854 41363 86922 41419
rect 86978 41363 87046 41419
rect 87102 41363 87126 41419
rect 86650 41344 87126 41363
rect 86526 41295 86630 41314
rect 86526 41239 86550 41295
rect 86606 41239 86630 41295
rect 86526 41171 86630 41239
rect 86526 41115 86550 41171
rect 86606 41115 86630 41171
rect 86526 41047 86630 41115
rect 86526 40991 86550 41047
rect 86606 40991 86630 41047
rect 86526 40923 86630 40991
rect 86526 40867 86550 40923
rect 86606 40867 86630 40923
rect 86526 40848 86630 40867
rect 86650 41295 87126 41314
rect 86650 41239 86674 41295
rect 86730 41239 86798 41295
rect 86854 41239 86922 41295
rect 86978 41239 87046 41295
rect 87102 41239 87126 41295
rect 86650 41171 87126 41239
rect 86650 41115 86674 41171
rect 86730 41115 86798 41171
rect 86854 41115 86922 41171
rect 86978 41115 87046 41171
rect 87102 41115 87126 41171
rect 86650 41047 87126 41115
rect 86650 40991 86674 41047
rect 86730 40991 86798 41047
rect 86854 40991 86922 41047
rect 86978 40991 87046 41047
rect 87102 40991 87126 41047
rect 86650 40923 87126 40991
rect 86650 40867 86674 40923
rect 86730 40867 86798 40923
rect 86854 40867 86922 40923
rect 86978 40867 87046 40923
rect 87102 40867 87126 40923
rect 86650 40848 87126 40867
rect 86526 40799 86630 40818
rect 86526 40743 86550 40799
rect 86606 40743 86630 40799
rect 86526 40675 86630 40743
rect 86526 40619 86550 40675
rect 86606 40619 86630 40675
rect 86526 40551 86630 40619
rect 1906 40501 2382 40532
rect 1906 40445 1930 40501
rect 1986 40445 2054 40501
rect 2110 40445 2178 40501
rect 2234 40445 2302 40501
rect 2358 40445 2382 40501
rect 1906 40377 2382 40445
rect 1906 40321 1930 40377
rect 1986 40321 2054 40377
rect 2110 40321 2178 40377
rect 2234 40321 2302 40377
rect 2358 40321 2382 40377
rect 86526 40495 86550 40551
rect 86606 40495 86630 40551
rect 86526 40427 86630 40495
rect 86526 40371 86550 40427
rect 86606 40371 86630 40427
rect 86526 40352 86630 40371
rect 86650 40799 87126 40818
rect 86650 40743 86674 40799
rect 86730 40743 86798 40799
rect 86854 40743 86922 40799
rect 86978 40743 87046 40799
rect 87102 40743 87126 40799
rect 86650 40675 87126 40743
rect 86650 40619 86674 40675
rect 86730 40619 86798 40675
rect 86854 40619 86922 40675
rect 86978 40619 87046 40675
rect 87102 40619 87126 40675
rect 86650 40551 87126 40619
rect 86650 40495 86674 40551
rect 86730 40495 86798 40551
rect 86854 40495 86922 40551
rect 86978 40495 87046 40551
rect 87102 40495 87126 40551
rect 86650 40427 87126 40495
rect 86650 40371 86674 40427
rect 86730 40371 86798 40427
rect 86854 40371 86922 40427
rect 86978 40371 87046 40427
rect 87102 40371 87126 40427
rect 86650 40352 87126 40371
rect 1906 40253 2382 40321
rect 1906 40197 1930 40253
rect 1986 40197 2054 40253
rect 2110 40197 2178 40253
rect 2234 40197 2302 40253
rect 2358 40197 2382 40253
rect 1906 40129 2382 40197
rect 1906 40073 1930 40129
rect 1986 40073 2054 40129
rect 2110 40073 2178 40129
rect 2234 40073 2302 40129
rect 2358 40073 2382 40129
rect 1906 40042 2382 40073
rect 86526 40303 86630 40322
rect 86526 40247 86550 40303
rect 86606 40247 86630 40303
rect 86526 40179 86630 40247
rect 86526 40123 86550 40179
rect 86606 40123 86630 40179
rect 86526 40055 86630 40123
rect 86526 39999 86550 40055
rect 86606 39999 86630 40055
rect 86526 39980 86630 39999
rect 86650 40303 87126 40322
rect 86650 40247 86674 40303
rect 86730 40247 86798 40303
rect 86854 40247 86922 40303
rect 86978 40247 87046 40303
rect 87102 40247 87126 40303
rect 86650 40179 87126 40247
rect 86650 40123 86674 40179
rect 86730 40123 86798 40179
rect 86854 40123 86922 40179
rect 86978 40123 87046 40179
rect 87102 40123 87126 40179
rect 86650 40055 87126 40123
rect 86650 39999 86674 40055
rect 86730 39999 86798 40055
rect 86854 39999 86922 40055
rect 86978 39999 87046 40055
rect 87102 39999 87126 40055
rect 86650 39980 87126 39999
rect 85726 39391 85830 39424
rect 85726 39335 85750 39391
rect 85806 39335 85830 39391
rect 85726 39267 85830 39335
rect 85726 39211 85750 39267
rect 85806 39211 85830 39267
rect 85726 39143 85830 39211
rect 85726 39087 85750 39143
rect 85806 39087 85830 39143
rect 85726 39019 85830 39087
rect 85726 38963 85750 39019
rect 85806 38963 85830 39019
rect 85726 38930 85830 38963
rect 85850 39391 86326 39424
rect 85850 39335 85874 39391
rect 85930 39335 85998 39391
rect 86054 39335 86122 39391
rect 86178 39335 86246 39391
rect 86302 39335 86326 39391
rect 85850 39267 86326 39335
rect 85850 39211 85874 39267
rect 85930 39211 85998 39267
rect 86054 39211 86122 39267
rect 86178 39211 86246 39267
rect 86302 39211 86326 39267
rect 85850 39143 86326 39211
rect 85850 39087 85874 39143
rect 85930 39087 85998 39143
rect 86054 39087 86122 39143
rect 86178 39087 86246 39143
rect 86302 39087 86326 39143
rect 85850 39019 86326 39087
rect 85850 38963 85874 39019
rect 85930 38963 85998 39019
rect 86054 38963 86122 39019
rect 86178 38963 86246 39019
rect 86302 38963 86326 39019
rect 85850 38930 86326 38963
rect 85726 38895 85830 38928
rect 85726 38839 85750 38895
rect 85806 38839 85830 38895
rect 85726 38771 85830 38839
rect 85726 38715 85750 38771
rect 85806 38715 85830 38771
rect 85726 38647 85830 38715
rect 85726 38591 85750 38647
rect 85806 38591 85830 38647
rect 85726 38523 85830 38591
rect 85726 38467 85750 38523
rect 85806 38467 85830 38523
rect 85726 38434 85830 38467
rect 85850 38895 86326 38928
rect 85850 38839 85874 38895
rect 85930 38839 85998 38895
rect 86054 38839 86122 38895
rect 86178 38839 86246 38895
rect 86302 38839 86326 38895
rect 85850 38771 86326 38839
rect 85850 38715 85874 38771
rect 85930 38715 85998 38771
rect 86054 38715 86122 38771
rect 86178 38715 86246 38771
rect 86302 38715 86326 38771
rect 85850 38647 86326 38715
rect 85850 38591 85874 38647
rect 85930 38591 85998 38647
rect 86054 38591 86122 38647
rect 86178 38591 86246 38647
rect 86302 38591 86326 38647
rect 85850 38523 86326 38591
rect 85850 38467 85874 38523
rect 85930 38467 85998 38523
rect 86054 38467 86122 38523
rect 86178 38467 86246 38523
rect 86302 38467 86326 38523
rect 85850 38434 86326 38467
rect 85726 38399 85830 38432
rect 85726 38343 85750 38399
rect 85806 38343 85830 38399
rect 85726 38275 85830 38343
rect 85726 38219 85750 38275
rect 85806 38219 85830 38275
rect 85726 38151 85830 38219
rect 85726 38095 85750 38151
rect 85806 38095 85830 38151
rect 85726 38062 85830 38095
rect 85850 38399 86326 38432
rect 85850 38343 85874 38399
rect 85930 38343 85998 38399
rect 86054 38343 86122 38399
rect 86178 38343 86246 38399
rect 86302 38343 86326 38399
rect 85850 38275 86326 38343
rect 85850 38219 85874 38275
rect 85930 38219 85998 38275
rect 86054 38219 86122 38275
rect 86178 38219 86246 38275
rect 86302 38219 86326 38275
rect 85850 38151 86326 38219
rect 85850 38095 85874 38151
rect 85930 38095 85998 38151
rect 86054 38095 86122 38151
rect 86178 38095 86246 38151
rect 86302 38095 86326 38151
rect 85850 38062 86326 38095
rect 1044 35489 1148 35540
rect 1044 35433 1068 35489
rect 1124 35433 1148 35489
rect 1044 35365 1148 35433
rect 1044 35309 1068 35365
rect 1124 35309 1148 35365
rect 1044 35241 1148 35309
rect 1044 35185 1068 35241
rect 1124 35185 1148 35241
rect 1044 35117 1148 35185
rect 1044 35061 1068 35117
rect 1124 35061 1148 35117
rect 1044 34993 1148 35061
rect 1044 34937 1068 34993
rect 1124 34937 1148 34993
rect 1044 34869 1148 34937
rect 1044 34813 1068 34869
rect 1124 34813 1148 34869
rect 1044 34745 1148 34813
rect 1044 34689 1068 34745
rect 1124 34689 1148 34745
rect 1044 34621 1148 34689
rect 1044 34565 1068 34621
rect 1124 34565 1148 34621
rect 1044 34497 1148 34565
rect 1044 34441 1068 34497
rect 1124 34441 1148 34497
rect 1044 34373 1148 34441
rect 1044 34317 1068 34373
rect 1124 34317 1148 34373
rect 1044 34249 1148 34317
rect 1044 34193 1068 34249
rect 1124 34193 1148 34249
rect 1044 34125 1148 34193
rect 1044 34069 1068 34125
rect 1124 34069 1148 34125
rect 1044 34001 1148 34069
rect 1044 33945 1068 34001
rect 1124 33945 1148 34001
rect 1044 33877 1148 33945
rect 1044 33821 1068 33877
rect 1124 33821 1148 33877
rect 1044 33753 1148 33821
rect 1044 33697 1068 33753
rect 1124 33697 1148 33753
rect 1044 33629 1148 33697
rect 1044 33573 1068 33629
rect 1124 33573 1148 33629
rect 1044 33505 1148 33573
rect 1044 33449 1068 33505
rect 1124 33449 1148 33505
rect 1044 33398 1148 33449
rect 1168 35489 1644 35540
rect 1168 35433 1192 35489
rect 1248 35433 1316 35489
rect 1372 35433 1440 35489
rect 1496 35433 1564 35489
rect 1620 35433 1644 35489
rect 1168 35365 1644 35433
rect 1168 35309 1192 35365
rect 1248 35309 1316 35365
rect 1372 35309 1440 35365
rect 1496 35309 1564 35365
rect 1620 35309 1644 35365
rect 1168 35241 1644 35309
rect 1168 35185 1192 35241
rect 1248 35185 1316 35241
rect 1372 35185 1440 35241
rect 1496 35185 1564 35241
rect 1620 35185 1644 35241
rect 1168 35117 1644 35185
rect 1168 35061 1192 35117
rect 1248 35061 1316 35117
rect 1372 35061 1440 35117
rect 1496 35061 1564 35117
rect 1620 35061 1644 35117
rect 1168 34993 1644 35061
rect 1168 34937 1192 34993
rect 1248 34937 1316 34993
rect 1372 34937 1440 34993
rect 1496 34937 1564 34993
rect 1620 34937 1644 34993
rect 1168 34869 1644 34937
rect 1168 34813 1192 34869
rect 1248 34813 1316 34869
rect 1372 34813 1440 34869
rect 1496 34813 1564 34869
rect 1620 34813 1644 34869
rect 1168 34745 1644 34813
rect 1168 34689 1192 34745
rect 1248 34689 1316 34745
rect 1372 34689 1440 34745
rect 1496 34689 1564 34745
rect 1620 34689 1644 34745
rect 1168 34621 1644 34689
rect 1168 34565 1192 34621
rect 1248 34565 1316 34621
rect 1372 34565 1440 34621
rect 1496 34565 1564 34621
rect 1620 34565 1644 34621
rect 1168 34497 1644 34565
rect 1168 34441 1192 34497
rect 1248 34441 1316 34497
rect 1372 34441 1440 34497
rect 1496 34441 1564 34497
rect 1620 34441 1644 34497
rect 1168 34373 1644 34441
rect 1168 34317 1192 34373
rect 1248 34317 1316 34373
rect 1372 34317 1440 34373
rect 1496 34317 1564 34373
rect 1620 34317 1644 34373
rect 1168 34249 1644 34317
rect 1168 34193 1192 34249
rect 1248 34193 1316 34249
rect 1372 34193 1440 34249
rect 1496 34193 1564 34249
rect 1620 34193 1644 34249
rect 1168 34125 1644 34193
rect 1168 34069 1192 34125
rect 1248 34069 1316 34125
rect 1372 34069 1440 34125
rect 1496 34069 1564 34125
rect 1620 34069 1644 34125
rect 1168 34001 1644 34069
rect 1168 33945 1192 34001
rect 1248 33945 1316 34001
rect 1372 33945 1440 34001
rect 1496 33945 1564 34001
rect 1620 33945 1644 34001
rect 1168 33877 1644 33945
rect 1168 33821 1192 33877
rect 1248 33821 1316 33877
rect 1372 33821 1440 33877
rect 1496 33821 1564 33877
rect 1620 33821 1644 33877
rect 1168 33753 1644 33821
rect 1168 33697 1192 33753
rect 1248 33697 1316 33753
rect 1372 33697 1440 33753
rect 1496 33697 1564 33753
rect 1620 33697 1644 33753
rect 1168 33629 1644 33697
rect 1168 33573 1192 33629
rect 1248 33573 1316 33629
rect 1372 33573 1440 33629
rect 1496 33573 1564 33629
rect 1620 33573 1644 33629
rect 1168 33505 1644 33573
rect 1168 33449 1192 33505
rect 1248 33449 1316 33505
rect 1372 33449 1440 33505
rect 1496 33449 1564 33505
rect 1620 33449 1644 33505
rect 1168 33398 1644 33449
rect 85726 35489 85830 35540
rect 85726 35433 85750 35489
rect 85806 35433 85830 35489
rect 85726 35365 85830 35433
rect 85726 35309 85750 35365
rect 85806 35309 85830 35365
rect 85726 35241 85830 35309
rect 85726 35185 85750 35241
rect 85806 35185 85830 35241
rect 85726 35117 85830 35185
rect 85726 35061 85750 35117
rect 85806 35061 85830 35117
rect 85726 34993 85830 35061
rect 85726 34937 85750 34993
rect 85806 34937 85830 34993
rect 85726 34869 85830 34937
rect 85726 34813 85750 34869
rect 85806 34813 85830 34869
rect 85726 34745 85830 34813
rect 85726 34689 85750 34745
rect 85806 34689 85830 34745
rect 85726 34621 85830 34689
rect 85726 34565 85750 34621
rect 85806 34565 85830 34621
rect 85726 34497 85830 34565
rect 85726 34441 85750 34497
rect 85806 34441 85830 34497
rect 85726 34373 85830 34441
rect 85726 34317 85750 34373
rect 85806 34317 85830 34373
rect 85726 34249 85830 34317
rect 85726 34193 85750 34249
rect 85806 34193 85830 34249
rect 85726 34125 85830 34193
rect 85726 34069 85750 34125
rect 85806 34069 85830 34125
rect 85726 34001 85830 34069
rect 85726 33945 85750 34001
rect 85806 33945 85830 34001
rect 85726 33877 85830 33945
rect 85726 33821 85750 33877
rect 85806 33821 85830 33877
rect 85726 33753 85830 33821
rect 85726 33697 85750 33753
rect 85806 33697 85830 33753
rect 85726 33629 85830 33697
rect 85726 33573 85750 33629
rect 85806 33573 85830 33629
rect 85726 33505 85830 33573
rect 85726 33449 85750 33505
rect 85806 33449 85830 33505
rect 85726 33398 85830 33449
rect 85850 35489 86326 35540
rect 85850 35433 85874 35489
rect 85930 35433 85998 35489
rect 86054 35433 86122 35489
rect 86178 35433 86246 35489
rect 86302 35433 86326 35489
rect 85850 35365 86326 35433
rect 85850 35309 85874 35365
rect 85930 35309 85998 35365
rect 86054 35309 86122 35365
rect 86178 35309 86246 35365
rect 86302 35309 86326 35365
rect 85850 35241 86326 35309
rect 85850 35185 85874 35241
rect 85930 35185 85998 35241
rect 86054 35185 86122 35241
rect 86178 35185 86246 35241
rect 86302 35185 86326 35241
rect 85850 35117 86326 35185
rect 85850 35061 85874 35117
rect 85930 35061 85998 35117
rect 86054 35061 86122 35117
rect 86178 35061 86246 35117
rect 86302 35061 86326 35117
rect 85850 34993 86326 35061
rect 85850 34937 85874 34993
rect 85930 34937 85998 34993
rect 86054 34937 86122 34993
rect 86178 34937 86246 34993
rect 86302 34937 86326 34993
rect 85850 34869 86326 34937
rect 85850 34813 85874 34869
rect 85930 34813 85998 34869
rect 86054 34813 86122 34869
rect 86178 34813 86246 34869
rect 86302 34813 86326 34869
rect 85850 34745 86326 34813
rect 85850 34689 85874 34745
rect 85930 34689 85998 34745
rect 86054 34689 86122 34745
rect 86178 34689 86246 34745
rect 86302 34689 86326 34745
rect 85850 34621 86326 34689
rect 85850 34565 85874 34621
rect 85930 34565 85998 34621
rect 86054 34565 86122 34621
rect 86178 34565 86246 34621
rect 86302 34565 86326 34621
rect 85850 34497 86326 34565
rect 85850 34441 85874 34497
rect 85930 34441 85998 34497
rect 86054 34441 86122 34497
rect 86178 34441 86246 34497
rect 86302 34441 86326 34497
rect 85850 34373 86326 34441
rect 85850 34317 85874 34373
rect 85930 34317 85998 34373
rect 86054 34317 86122 34373
rect 86178 34317 86246 34373
rect 86302 34317 86326 34373
rect 85850 34249 86326 34317
rect 85850 34193 85874 34249
rect 85930 34193 85998 34249
rect 86054 34193 86122 34249
rect 86178 34193 86246 34249
rect 86302 34193 86326 34249
rect 85850 34125 86326 34193
rect 85850 34069 85874 34125
rect 85930 34069 85998 34125
rect 86054 34069 86122 34125
rect 86178 34069 86246 34125
rect 86302 34069 86326 34125
rect 85850 34001 86326 34069
rect 85850 33945 85874 34001
rect 85930 33945 85998 34001
rect 86054 33945 86122 34001
rect 86178 33945 86246 34001
rect 86302 33945 86326 34001
rect 85850 33877 86326 33945
rect 85850 33821 85874 33877
rect 85930 33821 85998 33877
rect 86054 33821 86122 33877
rect 86178 33821 86246 33877
rect 86302 33821 86326 33877
rect 85850 33753 86326 33821
rect 85850 33697 85874 33753
rect 85930 33697 85998 33753
rect 86054 33697 86122 33753
rect 86178 33697 86246 33753
rect 86302 33697 86326 33753
rect 85850 33629 86326 33697
rect 85850 33573 85874 33629
rect 85930 33573 85998 33629
rect 86054 33573 86122 33629
rect 86178 33573 86246 33629
rect 86302 33573 86326 33629
rect 85850 33505 86326 33573
rect 85850 33449 85874 33505
rect 85930 33449 85998 33505
rect 86054 33449 86122 33505
rect 86178 33449 86246 33505
rect 86302 33449 86326 33505
rect 85850 33398 86326 33449
rect 1844 33187 1948 33248
rect 1844 33131 1868 33187
rect 1924 33131 1948 33187
rect 1844 33063 1948 33131
rect 1844 33007 1868 33063
rect 1924 33007 1948 33063
rect 1844 32939 1948 33007
rect 1844 32883 1868 32939
rect 1924 32883 1948 32939
rect 1844 32815 1948 32883
rect 1844 32759 1868 32815
rect 1924 32759 1948 32815
rect 1844 32691 1948 32759
rect 1844 32635 1868 32691
rect 1924 32635 1948 32691
rect 1844 32567 1948 32635
rect 1844 32511 1868 32567
rect 1924 32511 1948 32567
rect 1844 32443 1948 32511
rect 1844 32387 1868 32443
rect 1924 32387 1948 32443
rect 1844 32319 1948 32387
rect 1844 32263 1868 32319
rect 1924 32263 1948 32319
rect 1844 32195 1948 32263
rect 1844 32139 1868 32195
rect 1924 32139 1948 32195
rect 1844 32071 1948 32139
rect 1844 32015 1868 32071
rect 1924 32015 1948 32071
rect 1844 31947 1948 32015
rect 1844 31891 1868 31947
rect 1924 31891 1948 31947
rect 1844 31823 1948 31891
rect 1844 31767 1868 31823
rect 1924 31767 1948 31823
rect 1844 31699 1948 31767
rect 1844 31643 1868 31699
rect 1924 31643 1948 31699
rect 1844 31575 1948 31643
rect 1844 31519 1868 31575
rect 1924 31519 1948 31575
rect 1844 31451 1948 31519
rect 1844 31395 1868 31451
rect 1924 31395 1948 31451
rect 1844 31327 1948 31395
rect 1844 31271 1868 31327
rect 1924 31271 1948 31327
rect 1844 31203 1948 31271
rect 1844 31147 1868 31203
rect 1924 31147 1948 31203
rect 1844 31079 1948 31147
rect 1844 31023 1868 31079
rect 1924 31023 1948 31079
rect 1844 30955 1948 31023
rect 1844 30899 1868 30955
rect 1924 30899 1948 30955
rect 1844 30831 1948 30899
rect 1844 30775 1868 30831
rect 1924 30775 1948 30831
rect 1844 30707 1948 30775
rect 1844 30651 1868 30707
rect 1924 30651 1948 30707
rect 1844 30583 1948 30651
rect 1844 30527 1868 30583
rect 1924 30527 1948 30583
rect 1844 30459 1948 30527
rect 1844 30403 1868 30459
rect 1924 30403 1948 30459
rect 1844 30335 1948 30403
rect 1844 30279 1868 30335
rect 1924 30279 1948 30335
rect 1844 30211 1948 30279
rect 1844 30155 1868 30211
rect 1924 30155 1948 30211
rect 1844 30087 1948 30155
rect 1844 30031 1868 30087
rect 1924 30031 1948 30087
rect 1844 29963 1948 30031
rect 1844 29907 1868 29963
rect 1924 29907 1948 29963
rect 1844 29846 1948 29907
rect 1968 33187 2444 33248
rect 1968 33131 1992 33187
rect 2048 33131 2116 33187
rect 2172 33131 2240 33187
rect 2296 33131 2364 33187
rect 2420 33131 2444 33187
rect 1968 33063 2444 33131
rect 1968 33007 1992 33063
rect 2048 33007 2116 33063
rect 2172 33007 2240 33063
rect 2296 33007 2364 33063
rect 2420 33007 2444 33063
rect 1968 32939 2444 33007
rect 1968 32883 1992 32939
rect 2048 32883 2116 32939
rect 2172 32883 2240 32939
rect 2296 32883 2364 32939
rect 2420 32883 2444 32939
rect 1968 32815 2444 32883
rect 1968 32759 1992 32815
rect 2048 32759 2116 32815
rect 2172 32759 2240 32815
rect 2296 32759 2364 32815
rect 2420 32759 2444 32815
rect 1968 32691 2444 32759
rect 1968 32635 1992 32691
rect 2048 32635 2116 32691
rect 2172 32635 2240 32691
rect 2296 32635 2364 32691
rect 2420 32635 2444 32691
rect 1968 32567 2444 32635
rect 1968 32511 1992 32567
rect 2048 32511 2116 32567
rect 2172 32511 2240 32567
rect 2296 32511 2364 32567
rect 2420 32511 2444 32567
rect 1968 32443 2444 32511
rect 1968 32387 1992 32443
rect 2048 32387 2116 32443
rect 2172 32387 2240 32443
rect 2296 32387 2364 32443
rect 2420 32387 2444 32443
rect 1968 32319 2444 32387
rect 1968 32263 1992 32319
rect 2048 32263 2116 32319
rect 2172 32263 2240 32319
rect 2296 32263 2364 32319
rect 2420 32263 2444 32319
rect 1968 32195 2444 32263
rect 1968 32139 1992 32195
rect 2048 32139 2116 32195
rect 2172 32139 2240 32195
rect 2296 32139 2364 32195
rect 2420 32139 2444 32195
rect 1968 32071 2444 32139
rect 1968 32015 1992 32071
rect 2048 32015 2116 32071
rect 2172 32015 2240 32071
rect 2296 32015 2364 32071
rect 2420 32015 2444 32071
rect 1968 31947 2444 32015
rect 1968 31891 1992 31947
rect 2048 31891 2116 31947
rect 2172 31891 2240 31947
rect 2296 31891 2364 31947
rect 2420 31891 2444 31947
rect 1968 31823 2444 31891
rect 1968 31767 1992 31823
rect 2048 31767 2116 31823
rect 2172 31767 2240 31823
rect 2296 31767 2364 31823
rect 2420 31767 2444 31823
rect 1968 31699 2444 31767
rect 1968 31643 1992 31699
rect 2048 31643 2116 31699
rect 2172 31643 2240 31699
rect 2296 31643 2364 31699
rect 2420 31643 2444 31699
rect 1968 31575 2444 31643
rect 1968 31519 1992 31575
rect 2048 31519 2116 31575
rect 2172 31519 2240 31575
rect 2296 31519 2364 31575
rect 2420 31519 2444 31575
rect 1968 31451 2444 31519
rect 1968 31395 1992 31451
rect 2048 31395 2116 31451
rect 2172 31395 2240 31451
rect 2296 31395 2364 31451
rect 2420 31395 2444 31451
rect 1968 31327 2444 31395
rect 1968 31271 1992 31327
rect 2048 31271 2116 31327
rect 2172 31271 2240 31327
rect 2296 31271 2364 31327
rect 2420 31271 2444 31327
rect 1968 31203 2444 31271
rect 1968 31147 1992 31203
rect 2048 31147 2116 31203
rect 2172 31147 2240 31203
rect 2296 31147 2364 31203
rect 2420 31147 2444 31203
rect 1968 31079 2444 31147
rect 1968 31023 1992 31079
rect 2048 31023 2116 31079
rect 2172 31023 2240 31079
rect 2296 31023 2364 31079
rect 2420 31023 2444 31079
rect 1968 30955 2444 31023
rect 1968 30899 1992 30955
rect 2048 30899 2116 30955
rect 2172 30899 2240 30955
rect 2296 30899 2364 30955
rect 2420 30899 2444 30955
rect 1968 30831 2444 30899
rect 1968 30775 1992 30831
rect 2048 30775 2116 30831
rect 2172 30775 2240 30831
rect 2296 30775 2364 30831
rect 2420 30775 2444 30831
rect 1968 30707 2444 30775
rect 1968 30651 1992 30707
rect 2048 30651 2116 30707
rect 2172 30651 2240 30707
rect 2296 30651 2364 30707
rect 2420 30651 2444 30707
rect 1968 30583 2444 30651
rect 1968 30527 1992 30583
rect 2048 30527 2116 30583
rect 2172 30527 2240 30583
rect 2296 30527 2364 30583
rect 2420 30527 2444 30583
rect 1968 30459 2444 30527
rect 1968 30403 1992 30459
rect 2048 30403 2116 30459
rect 2172 30403 2240 30459
rect 2296 30403 2364 30459
rect 2420 30403 2444 30459
rect 1968 30335 2444 30403
rect 1968 30279 1992 30335
rect 2048 30279 2116 30335
rect 2172 30279 2240 30335
rect 2296 30279 2364 30335
rect 2420 30279 2444 30335
rect 1968 30211 2444 30279
rect 1968 30155 1992 30211
rect 2048 30155 2116 30211
rect 2172 30155 2240 30211
rect 2296 30155 2364 30211
rect 2420 30155 2444 30211
rect 1968 30087 2444 30155
rect 1968 30031 1992 30087
rect 2048 30031 2116 30087
rect 2172 30031 2240 30087
rect 2296 30031 2364 30087
rect 2420 30031 2444 30087
rect 1968 29963 2444 30031
rect 1968 29907 1992 29963
rect 2048 29907 2116 29963
rect 2172 29907 2240 29963
rect 2296 29907 2364 29963
rect 2420 29907 2444 29963
rect 1968 29846 2444 29907
rect 86526 33187 86630 33248
rect 86526 33131 86550 33187
rect 86606 33131 86630 33187
rect 86526 33063 86630 33131
rect 86526 33007 86550 33063
rect 86606 33007 86630 33063
rect 86526 32939 86630 33007
rect 86526 32883 86550 32939
rect 86606 32883 86630 32939
rect 86526 32815 86630 32883
rect 86526 32759 86550 32815
rect 86606 32759 86630 32815
rect 86526 32691 86630 32759
rect 86526 32635 86550 32691
rect 86606 32635 86630 32691
rect 86526 32567 86630 32635
rect 86526 32511 86550 32567
rect 86606 32511 86630 32567
rect 86526 32443 86630 32511
rect 86526 32387 86550 32443
rect 86606 32387 86630 32443
rect 86526 32319 86630 32387
rect 86526 32263 86550 32319
rect 86606 32263 86630 32319
rect 86526 32195 86630 32263
rect 86526 32139 86550 32195
rect 86606 32139 86630 32195
rect 86526 32071 86630 32139
rect 86526 32015 86550 32071
rect 86606 32015 86630 32071
rect 86526 31947 86630 32015
rect 86526 31891 86550 31947
rect 86606 31891 86630 31947
rect 86526 31823 86630 31891
rect 86526 31767 86550 31823
rect 86606 31767 86630 31823
rect 86526 31699 86630 31767
rect 86526 31643 86550 31699
rect 86606 31643 86630 31699
rect 86526 31575 86630 31643
rect 86526 31519 86550 31575
rect 86606 31519 86630 31575
rect 86526 31451 86630 31519
rect 86526 31395 86550 31451
rect 86606 31395 86630 31451
rect 86526 31327 86630 31395
rect 86526 31271 86550 31327
rect 86606 31271 86630 31327
rect 86526 31203 86630 31271
rect 86526 31147 86550 31203
rect 86606 31147 86630 31203
rect 86526 31079 86630 31147
rect 86526 31023 86550 31079
rect 86606 31023 86630 31079
rect 86526 30955 86630 31023
rect 86526 30899 86550 30955
rect 86606 30899 86630 30955
rect 86526 30831 86630 30899
rect 86526 30775 86550 30831
rect 86606 30775 86630 30831
rect 86526 30707 86630 30775
rect 86526 30651 86550 30707
rect 86606 30651 86630 30707
rect 86526 30583 86630 30651
rect 86526 30527 86550 30583
rect 86606 30527 86630 30583
rect 86526 30459 86630 30527
rect 86526 30403 86550 30459
rect 86606 30403 86630 30459
rect 86526 30335 86630 30403
rect 86526 30279 86550 30335
rect 86606 30279 86630 30335
rect 86526 30211 86630 30279
rect 86526 30155 86550 30211
rect 86606 30155 86630 30211
rect 86526 30087 86630 30155
rect 86526 30031 86550 30087
rect 86606 30031 86630 30087
rect 86526 29963 86630 30031
rect 86526 29907 86550 29963
rect 86606 29907 86630 29963
rect 86526 29846 86630 29907
rect 86650 33187 87126 33248
rect 86650 33131 86674 33187
rect 86730 33131 86798 33187
rect 86854 33131 86922 33187
rect 86978 33131 87046 33187
rect 87102 33131 87126 33187
rect 86650 33063 87126 33131
rect 86650 33007 86674 33063
rect 86730 33007 86798 33063
rect 86854 33007 86922 33063
rect 86978 33007 87046 33063
rect 87102 33007 87126 33063
rect 86650 32939 87126 33007
rect 86650 32883 86674 32939
rect 86730 32883 86798 32939
rect 86854 32883 86922 32939
rect 86978 32883 87046 32939
rect 87102 32883 87126 32939
rect 86650 32815 87126 32883
rect 86650 32759 86674 32815
rect 86730 32759 86798 32815
rect 86854 32759 86922 32815
rect 86978 32759 87046 32815
rect 87102 32759 87126 32815
rect 86650 32691 87126 32759
rect 86650 32635 86674 32691
rect 86730 32635 86798 32691
rect 86854 32635 86922 32691
rect 86978 32635 87046 32691
rect 87102 32635 87126 32691
rect 86650 32567 87126 32635
rect 86650 32511 86674 32567
rect 86730 32511 86798 32567
rect 86854 32511 86922 32567
rect 86978 32511 87046 32567
rect 87102 32511 87126 32567
rect 86650 32443 87126 32511
rect 86650 32387 86674 32443
rect 86730 32387 86798 32443
rect 86854 32387 86922 32443
rect 86978 32387 87046 32443
rect 87102 32387 87126 32443
rect 86650 32319 87126 32387
rect 86650 32263 86674 32319
rect 86730 32263 86798 32319
rect 86854 32263 86922 32319
rect 86978 32263 87046 32319
rect 87102 32263 87126 32319
rect 86650 32195 87126 32263
rect 86650 32139 86674 32195
rect 86730 32139 86798 32195
rect 86854 32139 86922 32195
rect 86978 32139 87046 32195
rect 87102 32139 87126 32195
rect 86650 32071 87126 32139
rect 86650 32015 86674 32071
rect 86730 32015 86798 32071
rect 86854 32015 86922 32071
rect 86978 32015 87046 32071
rect 87102 32015 87126 32071
rect 86650 31947 87126 32015
rect 86650 31891 86674 31947
rect 86730 31891 86798 31947
rect 86854 31891 86922 31947
rect 86978 31891 87046 31947
rect 87102 31891 87126 31947
rect 86650 31823 87126 31891
rect 86650 31767 86674 31823
rect 86730 31767 86798 31823
rect 86854 31767 86922 31823
rect 86978 31767 87046 31823
rect 87102 31767 87126 31823
rect 86650 31699 87126 31767
rect 86650 31643 86674 31699
rect 86730 31643 86798 31699
rect 86854 31643 86922 31699
rect 86978 31643 87046 31699
rect 87102 31643 87126 31699
rect 86650 31575 87126 31643
rect 86650 31519 86674 31575
rect 86730 31519 86798 31575
rect 86854 31519 86922 31575
rect 86978 31519 87046 31575
rect 87102 31519 87126 31575
rect 86650 31451 87126 31519
rect 86650 31395 86674 31451
rect 86730 31395 86798 31451
rect 86854 31395 86922 31451
rect 86978 31395 87046 31451
rect 87102 31395 87126 31451
rect 86650 31327 87126 31395
rect 86650 31271 86674 31327
rect 86730 31271 86798 31327
rect 86854 31271 86922 31327
rect 86978 31271 87046 31327
rect 87102 31271 87126 31327
rect 86650 31203 87126 31271
rect 86650 31147 86674 31203
rect 86730 31147 86798 31203
rect 86854 31147 86922 31203
rect 86978 31147 87046 31203
rect 87102 31147 87126 31203
rect 86650 31079 87126 31147
rect 86650 31023 86674 31079
rect 86730 31023 86798 31079
rect 86854 31023 86922 31079
rect 86978 31023 87046 31079
rect 87102 31023 87126 31079
rect 86650 30955 87126 31023
rect 86650 30899 86674 30955
rect 86730 30899 86798 30955
rect 86854 30899 86922 30955
rect 86978 30899 87046 30955
rect 87102 30899 87126 30955
rect 86650 30831 87126 30899
rect 86650 30775 86674 30831
rect 86730 30775 86798 30831
rect 86854 30775 86922 30831
rect 86978 30775 87046 30831
rect 87102 30775 87126 30831
rect 86650 30707 87126 30775
rect 86650 30651 86674 30707
rect 86730 30651 86798 30707
rect 86854 30651 86922 30707
rect 86978 30651 87046 30707
rect 87102 30651 87126 30707
rect 86650 30583 87126 30651
rect 86650 30527 86674 30583
rect 86730 30527 86798 30583
rect 86854 30527 86922 30583
rect 86978 30527 87046 30583
rect 87102 30527 87126 30583
rect 86650 30459 87126 30527
rect 86650 30403 86674 30459
rect 86730 30403 86798 30459
rect 86854 30403 86922 30459
rect 86978 30403 87046 30459
rect 87102 30403 87126 30459
rect 86650 30335 87126 30403
rect 86650 30279 86674 30335
rect 86730 30279 86798 30335
rect 86854 30279 86922 30335
rect 86978 30279 87046 30335
rect 87102 30279 87126 30335
rect 86650 30211 87126 30279
rect 86650 30155 86674 30211
rect 86730 30155 86798 30211
rect 86854 30155 86922 30211
rect 86978 30155 87046 30211
rect 87102 30155 87126 30211
rect 86650 30087 87126 30155
rect 86650 30031 86674 30087
rect 86730 30031 86798 30087
rect 86854 30031 86922 30087
rect 86978 30031 87046 30087
rect 87102 30031 87126 30087
rect 86650 29963 87126 30031
rect 86650 29907 86674 29963
rect 86730 29907 86798 29963
rect 86854 29907 86922 29963
rect 86978 29907 87046 29963
rect 87102 29907 87126 29963
rect 86650 29846 87126 29907
rect 86526 26256 86630 26294
rect 86526 26200 86550 26256
rect 86606 26200 86630 26256
rect 86526 26132 86630 26200
rect 86526 26076 86550 26132
rect 86606 26076 86630 26132
rect 86526 26008 86630 26076
rect 86526 25952 86550 26008
rect 86606 25952 86630 26008
rect 86526 25884 86630 25952
rect 86526 25828 86550 25884
rect 86606 25828 86630 25884
rect 86526 25760 86630 25828
rect 86526 25704 86550 25760
rect 86606 25704 86630 25760
rect 86526 25636 86630 25704
rect 86526 25580 86550 25636
rect 86606 25580 86630 25636
rect 86526 25512 86630 25580
rect 86526 25456 86550 25512
rect 86606 25456 86630 25512
rect 86526 25388 86630 25456
rect 86526 25332 86550 25388
rect 86606 25332 86630 25388
rect 86526 25294 86630 25332
rect 86650 26256 87126 26294
rect 86650 26200 86674 26256
rect 86730 26200 86798 26256
rect 86854 26200 86922 26256
rect 86978 26200 87046 26256
rect 87102 26200 87126 26256
rect 86650 26132 87126 26200
rect 86650 26076 86674 26132
rect 86730 26076 86798 26132
rect 86854 26076 86922 26132
rect 86978 26076 87046 26132
rect 87102 26076 87126 26132
rect 86650 26008 87126 26076
rect 86650 25952 86674 26008
rect 86730 25952 86798 26008
rect 86854 25952 86922 26008
rect 86978 25952 87046 26008
rect 87102 25952 87126 26008
rect 86650 25884 87126 25952
rect 86650 25828 86674 25884
rect 86730 25828 86798 25884
rect 86854 25828 86922 25884
rect 86978 25828 87046 25884
rect 87102 25828 87126 25884
rect 86650 25760 87126 25828
rect 86650 25704 86674 25760
rect 86730 25704 86798 25760
rect 86854 25704 86922 25760
rect 86978 25704 87046 25760
rect 87102 25704 87126 25760
rect 86650 25636 87126 25704
rect 86650 25580 86674 25636
rect 86730 25580 86798 25636
rect 86854 25580 86922 25636
rect 86978 25580 87046 25636
rect 87102 25580 87126 25636
rect 86650 25512 87126 25580
rect 86650 25456 86674 25512
rect 86730 25456 86798 25512
rect 86854 25456 86922 25512
rect 86978 25456 87046 25512
rect 87102 25456 87126 25512
rect 86650 25388 87126 25456
rect 86650 25332 86674 25388
rect 86730 25332 86798 25388
rect 86854 25332 86922 25388
rect 86978 25332 87046 25388
rect 87102 25332 87126 25388
rect 86650 25294 87126 25332
rect 1044 24600 1148 24638
rect 1044 24544 1068 24600
rect 1124 24544 1148 24600
rect 1044 24476 1148 24544
rect 1044 24420 1068 24476
rect 1124 24420 1148 24476
rect 1044 24352 1148 24420
rect 1044 24296 1068 24352
rect 1124 24296 1148 24352
rect 1044 24228 1148 24296
rect 1044 24172 1068 24228
rect 1124 24172 1148 24228
rect 1044 24104 1148 24172
rect 1044 24048 1068 24104
rect 1124 24048 1148 24104
rect 1044 23980 1148 24048
rect 1044 23924 1068 23980
rect 1124 23924 1148 23980
rect 1044 23856 1148 23924
rect 1044 23800 1068 23856
rect 1124 23800 1148 23856
rect 1044 23732 1148 23800
rect 1044 23676 1068 23732
rect 1124 23676 1148 23732
rect 1044 23638 1148 23676
rect 1168 24600 1644 24638
rect 1168 24544 1192 24600
rect 1248 24544 1316 24600
rect 1372 24544 1440 24600
rect 1496 24544 1564 24600
rect 1620 24544 1644 24600
rect 1168 24476 1644 24544
rect 1168 24420 1192 24476
rect 1248 24420 1316 24476
rect 1372 24420 1440 24476
rect 1496 24420 1564 24476
rect 1620 24420 1644 24476
rect 1168 24352 1644 24420
rect 1168 24296 1192 24352
rect 1248 24296 1316 24352
rect 1372 24296 1440 24352
rect 1496 24296 1564 24352
rect 1620 24296 1644 24352
rect 1168 24228 1644 24296
rect 1168 24172 1192 24228
rect 1248 24172 1316 24228
rect 1372 24172 1440 24228
rect 1496 24172 1564 24228
rect 1620 24172 1644 24228
rect 1168 24104 1644 24172
rect 1168 24048 1192 24104
rect 1248 24048 1316 24104
rect 1372 24048 1440 24104
rect 1496 24048 1564 24104
rect 1620 24048 1644 24104
rect 1168 23980 1644 24048
rect 1168 23924 1192 23980
rect 1248 23924 1316 23980
rect 1372 23924 1440 23980
rect 1496 23924 1564 23980
rect 1620 23924 1644 23980
rect 1168 23856 1644 23924
rect 1168 23800 1192 23856
rect 1248 23800 1316 23856
rect 1372 23800 1440 23856
rect 1496 23800 1564 23856
rect 1620 23800 1644 23856
rect 1168 23732 1644 23800
rect 1168 23676 1192 23732
rect 1248 23676 1316 23732
rect 1372 23676 1440 23732
rect 1496 23676 1564 23732
rect 1620 23676 1644 23732
rect 1168 23638 1644 23676
rect 85726 24600 85830 24638
rect 85726 24544 85750 24600
rect 85806 24544 85830 24600
rect 85726 24476 85830 24544
rect 85726 24420 85750 24476
rect 85806 24420 85830 24476
rect 85726 24352 85830 24420
rect 85726 24296 85750 24352
rect 85806 24296 85830 24352
rect 85726 24228 85830 24296
rect 85726 24172 85750 24228
rect 85806 24172 85830 24228
rect 85726 24104 85830 24172
rect 85726 24048 85750 24104
rect 85806 24048 85830 24104
rect 85726 23980 85830 24048
rect 85726 23924 85750 23980
rect 85806 23924 85830 23980
rect 85726 23856 85830 23924
rect 85726 23800 85750 23856
rect 85806 23800 85830 23856
rect 85726 23732 85830 23800
rect 85726 23676 85750 23732
rect 85806 23676 85830 23732
rect 85726 23638 85830 23676
rect 85850 24600 86326 24638
rect 85850 24544 85874 24600
rect 85930 24544 85998 24600
rect 86054 24544 86122 24600
rect 86178 24544 86246 24600
rect 86302 24544 86326 24600
rect 85850 24476 86326 24544
rect 85850 24420 85874 24476
rect 85930 24420 85998 24476
rect 86054 24420 86122 24476
rect 86178 24420 86246 24476
rect 86302 24420 86326 24476
rect 85850 24352 86326 24420
rect 85850 24296 85874 24352
rect 85930 24296 85998 24352
rect 86054 24296 86122 24352
rect 86178 24296 86246 24352
rect 86302 24296 86326 24352
rect 85850 24228 86326 24296
rect 85850 24172 85874 24228
rect 85930 24172 85998 24228
rect 86054 24172 86122 24228
rect 86178 24172 86246 24228
rect 86302 24172 86326 24228
rect 85850 24104 86326 24172
rect 85850 24048 85874 24104
rect 85930 24048 85998 24104
rect 86054 24048 86122 24104
rect 86178 24048 86246 24104
rect 86302 24048 86326 24104
rect 85850 23980 86326 24048
rect 85850 23924 85874 23980
rect 85930 23924 85998 23980
rect 86054 23924 86122 23980
rect 86178 23924 86246 23980
rect 86302 23924 86326 23980
rect 85850 23856 86326 23924
rect 85850 23800 85874 23856
rect 85930 23800 85998 23856
rect 86054 23800 86122 23856
rect 86178 23800 86246 23856
rect 86302 23800 86326 23856
rect 85850 23732 86326 23800
rect 85850 23676 85874 23732
rect 85930 23676 85998 23732
rect 86054 23676 86122 23732
rect 86178 23676 86246 23732
rect 86302 23676 86326 23732
rect 85850 23638 86326 23676
rect 1906 13014 2382 13040
rect 1906 12958 1930 13014
rect 1986 12958 2054 13014
rect 2110 12958 2178 13014
rect 2234 12958 2302 13014
rect 2358 12958 2382 13014
rect 1906 12890 2382 12958
rect 1906 12834 1930 12890
rect 1986 12834 2054 12890
rect 2110 12834 2178 12890
rect 2234 12834 2302 12890
rect 2358 12834 2382 12890
rect 1906 12766 2382 12834
rect 1906 12710 1930 12766
rect 1986 12710 2054 12766
rect 2110 12710 2178 12766
rect 2234 12710 2302 12766
rect 2358 12710 2382 12766
rect 1906 12642 2382 12710
rect 1906 12586 1930 12642
rect 1986 12586 2054 12642
rect 2110 12586 2178 12642
rect 2234 12586 2302 12642
rect 2358 12586 2382 12642
rect 1906 12560 2382 12586
rect 86588 12859 87064 12916
rect 86588 12803 86612 12859
rect 86668 12803 86736 12859
rect 86792 12803 86860 12859
rect 86916 12803 86984 12859
rect 87040 12803 87064 12859
rect 86588 12735 87064 12803
rect 86588 12679 86612 12735
rect 86668 12679 86736 12735
rect 86792 12679 86860 12735
rect 86916 12679 86984 12735
rect 87040 12679 87064 12735
rect 86588 12611 87064 12679
rect 86588 12555 86612 12611
rect 86668 12555 86736 12611
rect 86792 12555 86860 12611
rect 86916 12555 86984 12611
rect 87040 12555 87064 12611
rect 86588 12487 87064 12555
rect 86588 12431 86612 12487
rect 86668 12431 86736 12487
rect 86792 12431 86860 12487
rect 86916 12431 86984 12487
rect 87040 12431 87064 12487
rect 86588 12374 87064 12431
rect 1106 11664 1582 11676
rect 1106 11608 1130 11664
rect 1186 11608 1254 11664
rect 1310 11608 1378 11664
rect 1434 11608 1502 11664
rect 1558 11608 1582 11664
rect 1106 11540 1582 11608
rect 1106 11484 1130 11540
rect 1186 11484 1254 11540
rect 1310 11484 1378 11540
rect 1434 11484 1502 11540
rect 1558 11484 1582 11540
rect 1106 11416 1582 11484
rect 1106 11360 1130 11416
rect 1186 11360 1254 11416
rect 1310 11360 1378 11416
rect 1434 11360 1502 11416
rect 1558 11360 1582 11416
rect 1106 11292 1582 11360
rect 1106 11236 1130 11292
rect 1186 11236 1254 11292
rect 1310 11236 1378 11292
rect 1434 11236 1502 11292
rect 1558 11236 1582 11292
rect 1106 11224 1582 11236
rect 85788 11664 86264 11676
rect 85788 11608 85812 11664
rect 85868 11608 85936 11664
rect 85992 11608 86060 11664
rect 86116 11608 86184 11664
rect 86240 11608 86264 11664
rect 85788 11540 86264 11608
rect 85788 11484 85812 11540
rect 85868 11484 85936 11540
rect 85992 11484 86060 11540
rect 86116 11484 86184 11540
rect 86240 11484 86264 11540
rect 85788 11416 86264 11484
rect 85788 11360 85812 11416
rect 85868 11360 85936 11416
rect 85992 11360 86060 11416
rect 86116 11360 86184 11416
rect 86240 11360 86264 11416
rect 85788 11292 86264 11360
rect 85788 11236 85812 11292
rect 85868 11236 85936 11292
rect 85992 11236 86060 11292
rect 86116 11236 86184 11292
rect 86240 11236 86264 11292
rect 85788 11224 86264 11236
rect 86588 10764 87064 10776
rect 86588 10708 86612 10764
rect 86668 10708 86736 10764
rect 86792 10708 86860 10764
rect 86916 10708 86984 10764
rect 87040 10708 87064 10764
rect 1906 10640 2382 10700
rect 1906 10584 1930 10640
rect 1986 10584 2054 10640
rect 2110 10584 2178 10640
rect 2234 10584 2302 10640
rect 2358 10584 2382 10640
rect 1906 10516 2382 10584
rect 1906 10460 1930 10516
rect 1986 10460 2054 10516
rect 2110 10460 2178 10516
rect 2234 10460 2302 10516
rect 2358 10460 2382 10516
rect 1906 10400 2382 10460
rect 86588 10640 87064 10708
rect 86588 10584 86612 10640
rect 86668 10584 86736 10640
rect 86792 10584 86860 10640
rect 86916 10584 86984 10640
rect 87040 10584 87064 10640
rect 86588 10516 87064 10584
rect 86588 10460 86612 10516
rect 86668 10460 86736 10516
rect 86792 10460 86860 10516
rect 86916 10460 86984 10516
rect 87040 10460 87064 10516
rect 86588 10392 87064 10460
rect 86588 10336 86612 10392
rect 86668 10336 86736 10392
rect 86792 10336 86860 10392
rect 86916 10336 86984 10392
rect 87040 10336 87064 10392
rect 86588 10324 87064 10336
rect 1106 9864 1582 9876
rect 1106 9808 1130 9864
rect 1186 9808 1254 9864
rect 1310 9808 1378 9864
rect 1434 9808 1502 9864
rect 1558 9808 1582 9864
rect 1106 9740 1582 9808
rect 1106 9684 1130 9740
rect 1186 9684 1254 9740
rect 1310 9684 1378 9740
rect 1434 9684 1502 9740
rect 1558 9684 1582 9740
rect 1106 9616 1582 9684
rect 1106 9560 1130 9616
rect 1186 9560 1254 9616
rect 1310 9560 1378 9616
rect 1434 9560 1502 9616
rect 1558 9560 1582 9616
rect 1106 9492 1582 9560
rect 1106 9436 1130 9492
rect 1186 9436 1254 9492
rect 1310 9436 1378 9492
rect 1434 9436 1502 9492
rect 1558 9436 1582 9492
rect 1106 9424 1582 9436
rect 85788 9864 86264 9876
rect 85788 9808 85812 9864
rect 85868 9808 85936 9864
rect 85992 9808 86060 9864
rect 86116 9808 86184 9864
rect 86240 9808 86264 9864
rect 85788 9740 86264 9808
rect 85788 9684 85812 9740
rect 85868 9684 85936 9740
rect 85992 9684 86060 9740
rect 86116 9684 86184 9740
rect 86240 9684 86264 9740
rect 85788 9616 86264 9684
rect 85788 9560 85812 9616
rect 85868 9560 85936 9616
rect 85992 9560 86060 9616
rect 86116 9560 86184 9616
rect 86240 9560 86264 9616
rect 85788 9492 86264 9560
rect 85788 9436 85812 9492
rect 85868 9436 85936 9492
rect 85992 9436 86060 9492
rect 86116 9436 86184 9492
rect 86240 9436 86264 9492
rect 85788 9424 86264 9436
rect 86588 8964 87064 8976
rect 86588 8908 86612 8964
rect 86668 8908 86736 8964
rect 86792 8908 86860 8964
rect 86916 8908 86984 8964
rect 87040 8908 87064 8964
rect 1906 8840 2382 8900
rect 1906 8784 1930 8840
rect 1986 8784 2054 8840
rect 2110 8784 2178 8840
rect 2234 8784 2302 8840
rect 2358 8784 2382 8840
rect 1906 8716 2382 8784
rect 1906 8660 1930 8716
rect 1986 8660 2054 8716
rect 2110 8660 2178 8716
rect 2234 8660 2302 8716
rect 2358 8660 2382 8716
rect 1906 8600 2382 8660
rect 86588 8840 87064 8908
rect 86588 8784 86612 8840
rect 86668 8784 86736 8840
rect 86792 8784 86860 8840
rect 86916 8784 86984 8840
rect 87040 8784 87064 8840
rect 86588 8716 87064 8784
rect 86588 8660 86612 8716
rect 86668 8660 86736 8716
rect 86792 8660 86860 8716
rect 86916 8660 86984 8716
rect 87040 8660 87064 8716
rect 86588 8592 87064 8660
rect 86588 8536 86612 8592
rect 86668 8536 86736 8592
rect 86792 8536 86860 8592
rect 86916 8536 86984 8592
rect 87040 8536 87064 8592
rect 86588 8524 87064 8536
rect 1106 8064 1582 8076
rect 1106 8008 1130 8064
rect 1186 8008 1254 8064
rect 1310 8008 1378 8064
rect 1434 8008 1502 8064
rect 1558 8008 1582 8064
rect 1106 7940 1582 8008
rect 1106 7884 1130 7940
rect 1186 7884 1254 7940
rect 1310 7884 1378 7940
rect 1434 7884 1502 7940
rect 1558 7884 1582 7940
rect 1106 7816 1582 7884
rect 1106 7760 1130 7816
rect 1186 7760 1254 7816
rect 1310 7760 1378 7816
rect 1434 7760 1502 7816
rect 1558 7760 1582 7816
rect 1106 7692 1582 7760
rect 1106 7636 1130 7692
rect 1186 7636 1254 7692
rect 1310 7636 1378 7692
rect 1434 7636 1502 7692
rect 1558 7636 1582 7692
rect 1106 7624 1582 7636
rect 85788 8064 86264 8076
rect 85788 8008 85812 8064
rect 85868 8008 85936 8064
rect 85992 8008 86060 8064
rect 86116 8008 86184 8064
rect 86240 8008 86264 8064
rect 85788 7940 86264 8008
rect 85788 7884 85812 7940
rect 85868 7884 85936 7940
rect 85992 7884 86060 7940
rect 86116 7884 86184 7940
rect 86240 7884 86264 7940
rect 85788 7816 86264 7884
rect 85788 7760 85812 7816
rect 85868 7760 85936 7816
rect 85992 7760 86060 7816
rect 86116 7760 86184 7816
rect 86240 7760 86264 7816
rect 85788 7692 86264 7760
rect 85788 7636 85812 7692
rect 85868 7636 85936 7692
rect 85992 7636 86060 7692
rect 86116 7636 86184 7692
rect 86240 7636 86264 7692
rect 85788 7624 86264 7636
rect 86588 7164 87064 7176
rect 86588 7108 86612 7164
rect 86668 7108 86736 7164
rect 86792 7108 86860 7164
rect 86916 7108 86984 7164
rect 87040 7108 87064 7164
rect 1906 7040 2382 7100
rect 1906 6984 1930 7040
rect 1986 6984 2054 7040
rect 2110 6984 2178 7040
rect 2234 6984 2302 7040
rect 2358 6984 2382 7040
rect 1906 6916 2382 6984
rect 1906 6860 1930 6916
rect 1986 6860 2054 6916
rect 2110 6860 2178 6916
rect 2234 6860 2302 6916
rect 2358 6860 2382 6916
rect 1906 6800 2382 6860
rect 86588 7040 87064 7108
rect 86588 6984 86612 7040
rect 86668 6984 86736 7040
rect 86792 6984 86860 7040
rect 86916 6984 86984 7040
rect 87040 6984 87064 7040
rect 86588 6916 87064 6984
rect 86588 6860 86612 6916
rect 86668 6860 86736 6916
rect 86792 6860 86860 6916
rect 86916 6860 86984 6916
rect 87040 6860 87064 6916
rect 86588 6792 87064 6860
rect 86588 6736 86612 6792
rect 86668 6736 86736 6792
rect 86792 6736 86860 6792
rect 86916 6736 86984 6792
rect 87040 6736 87064 6792
rect 86588 6724 87064 6736
rect 1106 6264 1582 6276
rect 1106 6208 1130 6264
rect 1186 6208 1254 6264
rect 1310 6208 1378 6264
rect 1434 6208 1502 6264
rect 1558 6208 1582 6264
rect 1106 6140 1582 6208
rect 1106 6084 1130 6140
rect 1186 6084 1254 6140
rect 1310 6084 1378 6140
rect 1434 6084 1502 6140
rect 1558 6084 1582 6140
rect 1106 6016 1582 6084
rect 1106 5960 1130 6016
rect 1186 5960 1254 6016
rect 1310 5960 1378 6016
rect 1434 5960 1502 6016
rect 1558 5960 1582 6016
rect 1106 5892 1582 5960
rect 1106 5836 1130 5892
rect 1186 5836 1254 5892
rect 1310 5836 1378 5892
rect 1434 5836 1502 5892
rect 1558 5836 1582 5892
rect 1106 5824 1582 5836
rect 85788 6264 86264 6276
rect 85788 6208 85812 6264
rect 85868 6208 85936 6264
rect 85992 6208 86060 6264
rect 86116 6208 86184 6264
rect 86240 6208 86264 6264
rect 85788 6140 86264 6208
rect 85788 6084 85812 6140
rect 85868 6084 85936 6140
rect 85992 6084 86060 6140
rect 86116 6084 86184 6140
rect 86240 6084 86264 6140
rect 85788 6016 86264 6084
rect 85788 5960 85812 6016
rect 85868 5960 85936 6016
rect 85992 5960 86060 6016
rect 86116 5960 86184 6016
rect 86240 5960 86264 6016
rect 85788 5892 86264 5960
rect 85788 5836 85812 5892
rect 85868 5836 85936 5892
rect 85992 5836 86060 5892
rect 86116 5836 86184 5892
rect 86240 5836 86264 5892
rect 85788 5824 86264 5836
rect 86588 5364 87064 5376
rect 86588 5308 86612 5364
rect 86668 5308 86736 5364
rect 86792 5308 86860 5364
rect 86916 5308 86984 5364
rect 87040 5308 87064 5364
rect 1906 5240 2382 5300
rect 1906 5184 1930 5240
rect 1986 5184 2054 5240
rect 2110 5184 2178 5240
rect 2234 5184 2302 5240
rect 2358 5184 2382 5240
rect 1906 5116 2382 5184
rect 1906 5060 1930 5116
rect 1986 5060 2054 5116
rect 2110 5060 2178 5116
rect 2234 5060 2302 5116
rect 2358 5060 2382 5116
rect 1906 5000 2382 5060
rect 86588 5240 87064 5308
rect 86588 5184 86612 5240
rect 86668 5184 86736 5240
rect 86792 5184 86860 5240
rect 86916 5184 86984 5240
rect 87040 5184 87064 5240
rect 86588 5116 87064 5184
rect 86588 5060 86612 5116
rect 86668 5060 86736 5116
rect 86792 5060 86860 5116
rect 86916 5060 86984 5116
rect 87040 5060 87064 5116
rect 86588 4992 87064 5060
rect 86588 4936 86612 4992
rect 86668 4936 86736 4992
rect 86792 4936 86860 4992
rect 86916 4936 86984 4992
rect 87040 4936 87064 4992
rect 86588 4924 87064 4936
rect 1106 4464 1582 4476
rect 1106 4408 1130 4464
rect 1186 4408 1254 4464
rect 1310 4408 1378 4464
rect 1434 4408 1502 4464
rect 1558 4408 1582 4464
rect 1106 4340 1582 4408
rect 1106 4284 1130 4340
rect 1186 4284 1254 4340
rect 1310 4284 1378 4340
rect 1434 4284 1502 4340
rect 1558 4284 1582 4340
rect 1106 4216 1582 4284
rect 1106 4160 1130 4216
rect 1186 4160 1254 4216
rect 1310 4160 1378 4216
rect 1434 4160 1502 4216
rect 1558 4160 1582 4216
rect 1106 4092 1582 4160
rect 1106 4036 1130 4092
rect 1186 4036 1254 4092
rect 1310 4036 1378 4092
rect 1434 4036 1502 4092
rect 1558 4036 1582 4092
rect 1106 4024 1582 4036
rect 85788 4464 86264 4476
rect 85788 4408 85812 4464
rect 85868 4408 85936 4464
rect 85992 4408 86060 4464
rect 86116 4408 86184 4464
rect 86240 4408 86264 4464
rect 85788 4340 86264 4408
rect 85788 4284 85812 4340
rect 85868 4284 85936 4340
rect 85992 4284 86060 4340
rect 86116 4284 86184 4340
rect 86240 4284 86264 4340
rect 85788 4216 86264 4284
rect 85788 4160 85812 4216
rect 85868 4160 85936 4216
rect 85992 4160 86060 4216
rect 86116 4160 86184 4216
rect 86240 4160 86264 4216
rect 85788 4092 86264 4160
rect 85788 4036 85812 4092
rect 85868 4036 85936 4092
rect 85992 4036 86060 4092
rect 86116 4036 86184 4092
rect 86240 4036 86264 4092
rect 85788 4024 86264 4036
rect 86588 3632 87064 3700
rect 86588 3576 86612 3632
rect 86668 3576 86736 3632
rect 86792 3576 86860 3632
rect 86916 3576 86984 3632
rect 87040 3576 87064 3632
rect 86588 3508 87064 3576
rect 1906 3440 2382 3500
rect 1906 3384 1930 3440
rect 1986 3384 2054 3440
rect 2110 3384 2178 3440
rect 2234 3384 2302 3440
rect 2358 3384 2382 3440
rect 1906 3316 2382 3384
rect 1906 3260 1930 3316
rect 1986 3260 2054 3316
rect 2110 3260 2178 3316
rect 2234 3260 2302 3316
rect 2358 3260 2382 3316
rect 1906 3200 2382 3260
rect 86588 3452 86612 3508
rect 86668 3452 86736 3508
rect 86792 3452 86860 3508
rect 86916 3452 86984 3508
rect 87040 3452 87064 3508
rect 86588 3384 87064 3452
rect 86588 3328 86612 3384
rect 86668 3328 86736 3384
rect 86792 3328 86860 3384
rect 86916 3328 86984 3384
rect 87040 3328 87064 3384
rect 86588 3260 87064 3328
rect 86588 3204 86612 3260
rect 86668 3204 86736 3260
rect 86792 3204 86860 3260
rect 86916 3204 86984 3260
rect 87040 3204 87064 3260
rect 86588 3136 87064 3204
<< via3 >>
rect 1130 45380 1186 45436
rect 1254 45380 1310 45436
rect 1378 45380 1434 45436
rect 1502 45380 1558 45436
rect 85812 45380 85868 45436
rect 85936 45380 85992 45436
rect 86060 45380 86116 45436
rect 86184 45380 86240 45436
rect 1901 44969 1957 45025
rect 1901 44845 1957 44901
rect 1901 44721 1957 44777
rect 1901 44597 1957 44653
rect 1901 44473 1957 44529
rect 1901 44349 1957 44405
rect 1901 44225 1957 44281
rect 1901 44101 1957 44157
rect 1901 43977 1957 44033
rect 1901 43853 1957 43909
rect 86550 44969 86606 45025
rect 86550 44845 86606 44901
rect 86550 44721 86606 44777
rect 86550 44597 86606 44653
rect 86550 44473 86606 44529
rect 86550 44349 86606 44405
rect 86550 44225 86606 44281
rect 86550 44101 86606 44157
rect 86550 43977 86606 44033
rect 86550 43853 86606 43909
rect 86674 44969 86730 45025
rect 86798 44969 86854 45025
rect 86922 44969 86978 45025
rect 87046 44969 87102 45025
rect 86674 44845 86730 44901
rect 86798 44845 86854 44901
rect 86922 44845 86978 44901
rect 87046 44845 87102 44901
rect 86674 44721 86730 44777
rect 86798 44721 86854 44777
rect 86922 44721 86978 44777
rect 87046 44721 87102 44777
rect 86674 44597 86730 44653
rect 86798 44597 86854 44653
rect 86922 44597 86978 44653
rect 87046 44597 87102 44653
rect 86674 44473 86730 44529
rect 86798 44473 86854 44529
rect 86922 44473 86978 44529
rect 87046 44473 87102 44529
rect 86674 44349 86730 44405
rect 86798 44349 86854 44405
rect 86922 44349 86978 44405
rect 87046 44349 87102 44405
rect 86674 44225 86730 44281
rect 86798 44225 86854 44281
rect 86922 44225 86978 44281
rect 87046 44225 87102 44281
rect 86674 44101 86730 44157
rect 86798 44101 86854 44157
rect 86922 44101 86978 44157
rect 87046 44101 87102 44157
rect 86674 43977 86730 44033
rect 86798 43977 86854 44033
rect 86922 43977 86978 44033
rect 87046 43977 87102 44033
rect 86674 43853 86730 43909
rect 86798 43853 86854 43909
rect 86922 43853 86978 43909
rect 87046 43853 87102 43909
rect 86550 41735 86606 41791
rect 86550 41611 86606 41667
rect 86550 41487 86606 41543
rect 86550 41363 86606 41419
rect 86674 41735 86730 41791
rect 86798 41735 86854 41791
rect 86922 41735 86978 41791
rect 87046 41735 87102 41791
rect 86674 41611 86730 41667
rect 86798 41611 86854 41667
rect 86922 41611 86978 41667
rect 87046 41611 87102 41667
rect 86674 41487 86730 41543
rect 86798 41487 86854 41543
rect 86922 41487 86978 41543
rect 87046 41487 87102 41543
rect 86674 41363 86730 41419
rect 86798 41363 86854 41419
rect 86922 41363 86978 41419
rect 87046 41363 87102 41419
rect 86550 41239 86606 41295
rect 86550 41115 86606 41171
rect 86550 40991 86606 41047
rect 86550 40867 86606 40923
rect 86674 41239 86730 41295
rect 86798 41239 86854 41295
rect 86922 41239 86978 41295
rect 87046 41239 87102 41295
rect 86674 41115 86730 41171
rect 86798 41115 86854 41171
rect 86922 41115 86978 41171
rect 87046 41115 87102 41171
rect 86674 40991 86730 41047
rect 86798 40991 86854 41047
rect 86922 40991 86978 41047
rect 87046 40991 87102 41047
rect 86674 40867 86730 40923
rect 86798 40867 86854 40923
rect 86922 40867 86978 40923
rect 87046 40867 87102 40923
rect 86550 40743 86606 40799
rect 86550 40619 86606 40675
rect 1930 40445 1986 40501
rect 2054 40445 2110 40501
rect 2178 40445 2234 40501
rect 2302 40445 2358 40501
rect 1930 40321 1986 40377
rect 2054 40321 2110 40377
rect 2178 40321 2234 40377
rect 2302 40321 2358 40377
rect 86550 40495 86606 40551
rect 86550 40371 86606 40427
rect 86674 40743 86730 40799
rect 86798 40743 86854 40799
rect 86922 40743 86978 40799
rect 87046 40743 87102 40799
rect 86674 40619 86730 40675
rect 86798 40619 86854 40675
rect 86922 40619 86978 40675
rect 87046 40619 87102 40675
rect 86674 40495 86730 40551
rect 86798 40495 86854 40551
rect 86922 40495 86978 40551
rect 87046 40495 87102 40551
rect 86674 40371 86730 40427
rect 86798 40371 86854 40427
rect 86922 40371 86978 40427
rect 87046 40371 87102 40427
rect 1930 40197 1986 40253
rect 2054 40197 2110 40253
rect 2178 40197 2234 40253
rect 2302 40197 2358 40253
rect 1930 40073 1986 40129
rect 2054 40073 2110 40129
rect 2178 40073 2234 40129
rect 2302 40073 2358 40129
rect 86550 40247 86606 40303
rect 86550 40123 86606 40179
rect 86550 39999 86606 40055
rect 86674 40247 86730 40303
rect 86798 40247 86854 40303
rect 86922 40247 86978 40303
rect 87046 40247 87102 40303
rect 86674 40123 86730 40179
rect 86798 40123 86854 40179
rect 86922 40123 86978 40179
rect 87046 40123 87102 40179
rect 86674 39999 86730 40055
rect 86798 39999 86854 40055
rect 86922 39999 86978 40055
rect 87046 39999 87102 40055
rect 85750 39335 85806 39391
rect 85750 39211 85806 39267
rect 85750 39087 85806 39143
rect 85750 38963 85806 39019
rect 85874 39335 85930 39391
rect 85998 39335 86054 39391
rect 86122 39335 86178 39391
rect 86246 39335 86302 39391
rect 85874 39211 85930 39267
rect 85998 39211 86054 39267
rect 86122 39211 86178 39267
rect 86246 39211 86302 39267
rect 85874 39087 85930 39143
rect 85998 39087 86054 39143
rect 86122 39087 86178 39143
rect 86246 39087 86302 39143
rect 85874 38963 85930 39019
rect 85998 38963 86054 39019
rect 86122 38963 86178 39019
rect 86246 38963 86302 39019
rect 85750 38839 85806 38895
rect 85750 38715 85806 38771
rect 85750 38591 85806 38647
rect 85750 38467 85806 38523
rect 85874 38839 85930 38895
rect 85998 38839 86054 38895
rect 86122 38839 86178 38895
rect 86246 38839 86302 38895
rect 85874 38715 85930 38771
rect 85998 38715 86054 38771
rect 86122 38715 86178 38771
rect 86246 38715 86302 38771
rect 85874 38591 85930 38647
rect 85998 38591 86054 38647
rect 86122 38591 86178 38647
rect 86246 38591 86302 38647
rect 85874 38467 85930 38523
rect 85998 38467 86054 38523
rect 86122 38467 86178 38523
rect 86246 38467 86302 38523
rect 85750 38343 85806 38399
rect 85750 38219 85806 38275
rect 85750 38095 85806 38151
rect 85874 38343 85930 38399
rect 85998 38343 86054 38399
rect 86122 38343 86178 38399
rect 86246 38343 86302 38399
rect 85874 38219 85930 38275
rect 85998 38219 86054 38275
rect 86122 38219 86178 38275
rect 86246 38219 86302 38275
rect 85874 38095 85930 38151
rect 85998 38095 86054 38151
rect 86122 38095 86178 38151
rect 86246 38095 86302 38151
rect 1068 35433 1124 35489
rect 1068 35309 1124 35365
rect 1068 35185 1124 35241
rect 1068 35061 1124 35117
rect 1068 34937 1124 34993
rect 1068 34813 1124 34869
rect 1068 34689 1124 34745
rect 1068 34565 1124 34621
rect 1068 34441 1124 34497
rect 1068 34317 1124 34373
rect 1068 34193 1124 34249
rect 1068 34069 1124 34125
rect 1068 33945 1124 34001
rect 1068 33821 1124 33877
rect 1068 33697 1124 33753
rect 1068 33573 1124 33629
rect 1068 33449 1124 33505
rect 1192 35433 1248 35489
rect 1316 35433 1372 35489
rect 1440 35433 1496 35489
rect 1564 35433 1620 35489
rect 1192 35309 1248 35365
rect 1316 35309 1372 35365
rect 1440 35309 1496 35365
rect 1564 35309 1620 35365
rect 1192 35185 1248 35241
rect 1316 35185 1372 35241
rect 1440 35185 1496 35241
rect 1564 35185 1620 35241
rect 1192 35061 1248 35117
rect 1316 35061 1372 35117
rect 1440 35061 1496 35117
rect 1564 35061 1620 35117
rect 1192 34937 1248 34993
rect 1316 34937 1372 34993
rect 1440 34937 1496 34993
rect 1564 34937 1620 34993
rect 1192 34813 1248 34869
rect 1316 34813 1372 34869
rect 1440 34813 1496 34869
rect 1564 34813 1620 34869
rect 1192 34689 1248 34745
rect 1316 34689 1372 34745
rect 1440 34689 1496 34745
rect 1564 34689 1620 34745
rect 1192 34565 1248 34621
rect 1316 34565 1372 34621
rect 1440 34565 1496 34621
rect 1564 34565 1620 34621
rect 1192 34441 1248 34497
rect 1316 34441 1372 34497
rect 1440 34441 1496 34497
rect 1564 34441 1620 34497
rect 1192 34317 1248 34373
rect 1316 34317 1372 34373
rect 1440 34317 1496 34373
rect 1564 34317 1620 34373
rect 1192 34193 1248 34249
rect 1316 34193 1372 34249
rect 1440 34193 1496 34249
rect 1564 34193 1620 34249
rect 1192 34069 1248 34125
rect 1316 34069 1372 34125
rect 1440 34069 1496 34125
rect 1564 34069 1620 34125
rect 1192 33945 1248 34001
rect 1316 33945 1372 34001
rect 1440 33945 1496 34001
rect 1564 33945 1620 34001
rect 1192 33821 1248 33877
rect 1316 33821 1372 33877
rect 1440 33821 1496 33877
rect 1564 33821 1620 33877
rect 1192 33697 1248 33753
rect 1316 33697 1372 33753
rect 1440 33697 1496 33753
rect 1564 33697 1620 33753
rect 1192 33573 1248 33629
rect 1316 33573 1372 33629
rect 1440 33573 1496 33629
rect 1564 33573 1620 33629
rect 1192 33449 1248 33505
rect 1316 33449 1372 33505
rect 1440 33449 1496 33505
rect 1564 33449 1620 33505
rect 85750 35433 85806 35489
rect 85750 35309 85806 35365
rect 85750 35185 85806 35241
rect 85750 35061 85806 35117
rect 85750 34937 85806 34993
rect 85750 34813 85806 34869
rect 85750 34689 85806 34745
rect 85750 34565 85806 34621
rect 85750 34441 85806 34497
rect 85750 34317 85806 34373
rect 85750 34193 85806 34249
rect 85750 34069 85806 34125
rect 85750 33945 85806 34001
rect 85750 33821 85806 33877
rect 85750 33697 85806 33753
rect 85750 33573 85806 33629
rect 85750 33449 85806 33505
rect 85874 35433 85930 35489
rect 85998 35433 86054 35489
rect 86122 35433 86178 35489
rect 86246 35433 86302 35489
rect 85874 35309 85930 35365
rect 85998 35309 86054 35365
rect 86122 35309 86178 35365
rect 86246 35309 86302 35365
rect 85874 35185 85930 35241
rect 85998 35185 86054 35241
rect 86122 35185 86178 35241
rect 86246 35185 86302 35241
rect 85874 35061 85930 35117
rect 85998 35061 86054 35117
rect 86122 35061 86178 35117
rect 86246 35061 86302 35117
rect 85874 34937 85930 34993
rect 85998 34937 86054 34993
rect 86122 34937 86178 34993
rect 86246 34937 86302 34993
rect 85874 34813 85930 34869
rect 85998 34813 86054 34869
rect 86122 34813 86178 34869
rect 86246 34813 86302 34869
rect 85874 34689 85930 34745
rect 85998 34689 86054 34745
rect 86122 34689 86178 34745
rect 86246 34689 86302 34745
rect 85874 34565 85930 34621
rect 85998 34565 86054 34621
rect 86122 34565 86178 34621
rect 86246 34565 86302 34621
rect 85874 34441 85930 34497
rect 85998 34441 86054 34497
rect 86122 34441 86178 34497
rect 86246 34441 86302 34497
rect 85874 34317 85930 34373
rect 85998 34317 86054 34373
rect 86122 34317 86178 34373
rect 86246 34317 86302 34373
rect 85874 34193 85930 34249
rect 85998 34193 86054 34249
rect 86122 34193 86178 34249
rect 86246 34193 86302 34249
rect 85874 34069 85930 34125
rect 85998 34069 86054 34125
rect 86122 34069 86178 34125
rect 86246 34069 86302 34125
rect 85874 33945 85930 34001
rect 85998 33945 86054 34001
rect 86122 33945 86178 34001
rect 86246 33945 86302 34001
rect 85874 33821 85930 33877
rect 85998 33821 86054 33877
rect 86122 33821 86178 33877
rect 86246 33821 86302 33877
rect 85874 33697 85930 33753
rect 85998 33697 86054 33753
rect 86122 33697 86178 33753
rect 86246 33697 86302 33753
rect 85874 33573 85930 33629
rect 85998 33573 86054 33629
rect 86122 33573 86178 33629
rect 86246 33573 86302 33629
rect 85874 33449 85930 33505
rect 85998 33449 86054 33505
rect 86122 33449 86178 33505
rect 86246 33449 86302 33505
rect 1868 33131 1924 33187
rect 1868 33007 1924 33063
rect 1868 32883 1924 32939
rect 1868 32759 1924 32815
rect 1868 32635 1924 32691
rect 1868 32511 1924 32567
rect 1868 32387 1924 32443
rect 1868 32263 1924 32319
rect 1868 32139 1924 32195
rect 1868 32015 1924 32071
rect 1868 31891 1924 31947
rect 1868 31767 1924 31823
rect 1868 31643 1924 31699
rect 1868 31519 1924 31575
rect 1868 31395 1924 31451
rect 1868 31271 1924 31327
rect 1868 31147 1924 31203
rect 1868 31023 1924 31079
rect 1868 30899 1924 30955
rect 1868 30775 1924 30831
rect 1868 30651 1924 30707
rect 1868 30527 1924 30583
rect 1868 30403 1924 30459
rect 1868 30279 1924 30335
rect 1868 30155 1924 30211
rect 1868 30031 1924 30087
rect 1868 29907 1924 29963
rect 1992 33131 2048 33187
rect 2116 33131 2172 33187
rect 2240 33131 2296 33187
rect 2364 33131 2420 33187
rect 1992 33007 2048 33063
rect 2116 33007 2172 33063
rect 2240 33007 2296 33063
rect 2364 33007 2420 33063
rect 1992 32883 2048 32939
rect 2116 32883 2172 32939
rect 2240 32883 2296 32939
rect 2364 32883 2420 32939
rect 1992 32759 2048 32815
rect 2116 32759 2172 32815
rect 2240 32759 2296 32815
rect 2364 32759 2420 32815
rect 1992 32635 2048 32691
rect 2116 32635 2172 32691
rect 2240 32635 2296 32691
rect 2364 32635 2420 32691
rect 1992 32511 2048 32567
rect 2116 32511 2172 32567
rect 2240 32511 2296 32567
rect 2364 32511 2420 32567
rect 1992 32387 2048 32443
rect 2116 32387 2172 32443
rect 2240 32387 2296 32443
rect 2364 32387 2420 32443
rect 1992 32263 2048 32319
rect 2116 32263 2172 32319
rect 2240 32263 2296 32319
rect 2364 32263 2420 32319
rect 1992 32139 2048 32195
rect 2116 32139 2172 32195
rect 2240 32139 2296 32195
rect 2364 32139 2420 32195
rect 1992 32015 2048 32071
rect 2116 32015 2172 32071
rect 2240 32015 2296 32071
rect 2364 32015 2420 32071
rect 1992 31891 2048 31947
rect 2116 31891 2172 31947
rect 2240 31891 2296 31947
rect 2364 31891 2420 31947
rect 1992 31767 2048 31823
rect 2116 31767 2172 31823
rect 2240 31767 2296 31823
rect 2364 31767 2420 31823
rect 1992 31643 2048 31699
rect 2116 31643 2172 31699
rect 2240 31643 2296 31699
rect 2364 31643 2420 31699
rect 1992 31519 2048 31575
rect 2116 31519 2172 31575
rect 2240 31519 2296 31575
rect 2364 31519 2420 31575
rect 1992 31395 2048 31451
rect 2116 31395 2172 31451
rect 2240 31395 2296 31451
rect 2364 31395 2420 31451
rect 1992 31271 2048 31327
rect 2116 31271 2172 31327
rect 2240 31271 2296 31327
rect 2364 31271 2420 31327
rect 1992 31147 2048 31203
rect 2116 31147 2172 31203
rect 2240 31147 2296 31203
rect 2364 31147 2420 31203
rect 1992 31023 2048 31079
rect 2116 31023 2172 31079
rect 2240 31023 2296 31079
rect 2364 31023 2420 31079
rect 1992 30899 2048 30955
rect 2116 30899 2172 30955
rect 2240 30899 2296 30955
rect 2364 30899 2420 30955
rect 1992 30775 2048 30831
rect 2116 30775 2172 30831
rect 2240 30775 2296 30831
rect 2364 30775 2420 30831
rect 1992 30651 2048 30707
rect 2116 30651 2172 30707
rect 2240 30651 2296 30707
rect 2364 30651 2420 30707
rect 1992 30527 2048 30583
rect 2116 30527 2172 30583
rect 2240 30527 2296 30583
rect 2364 30527 2420 30583
rect 1992 30403 2048 30459
rect 2116 30403 2172 30459
rect 2240 30403 2296 30459
rect 2364 30403 2420 30459
rect 1992 30279 2048 30335
rect 2116 30279 2172 30335
rect 2240 30279 2296 30335
rect 2364 30279 2420 30335
rect 1992 30155 2048 30211
rect 2116 30155 2172 30211
rect 2240 30155 2296 30211
rect 2364 30155 2420 30211
rect 1992 30031 2048 30087
rect 2116 30031 2172 30087
rect 2240 30031 2296 30087
rect 2364 30031 2420 30087
rect 1992 29907 2048 29963
rect 2116 29907 2172 29963
rect 2240 29907 2296 29963
rect 2364 29907 2420 29963
rect 86550 33131 86606 33187
rect 86550 33007 86606 33063
rect 86550 32883 86606 32939
rect 86550 32759 86606 32815
rect 86550 32635 86606 32691
rect 86550 32511 86606 32567
rect 86550 32387 86606 32443
rect 86550 32263 86606 32319
rect 86550 32139 86606 32195
rect 86550 32015 86606 32071
rect 86550 31891 86606 31947
rect 86550 31767 86606 31823
rect 86550 31643 86606 31699
rect 86550 31519 86606 31575
rect 86550 31395 86606 31451
rect 86550 31271 86606 31327
rect 86550 31147 86606 31203
rect 86550 31023 86606 31079
rect 86550 30899 86606 30955
rect 86550 30775 86606 30831
rect 86550 30651 86606 30707
rect 86550 30527 86606 30583
rect 86550 30403 86606 30459
rect 86550 30279 86606 30335
rect 86550 30155 86606 30211
rect 86550 30031 86606 30087
rect 86550 29907 86606 29963
rect 86674 33131 86730 33187
rect 86798 33131 86854 33187
rect 86922 33131 86978 33187
rect 87046 33131 87102 33187
rect 86674 33007 86730 33063
rect 86798 33007 86854 33063
rect 86922 33007 86978 33063
rect 87046 33007 87102 33063
rect 86674 32883 86730 32939
rect 86798 32883 86854 32939
rect 86922 32883 86978 32939
rect 87046 32883 87102 32939
rect 86674 32759 86730 32815
rect 86798 32759 86854 32815
rect 86922 32759 86978 32815
rect 87046 32759 87102 32815
rect 86674 32635 86730 32691
rect 86798 32635 86854 32691
rect 86922 32635 86978 32691
rect 87046 32635 87102 32691
rect 86674 32511 86730 32567
rect 86798 32511 86854 32567
rect 86922 32511 86978 32567
rect 87046 32511 87102 32567
rect 86674 32387 86730 32443
rect 86798 32387 86854 32443
rect 86922 32387 86978 32443
rect 87046 32387 87102 32443
rect 86674 32263 86730 32319
rect 86798 32263 86854 32319
rect 86922 32263 86978 32319
rect 87046 32263 87102 32319
rect 86674 32139 86730 32195
rect 86798 32139 86854 32195
rect 86922 32139 86978 32195
rect 87046 32139 87102 32195
rect 86674 32015 86730 32071
rect 86798 32015 86854 32071
rect 86922 32015 86978 32071
rect 87046 32015 87102 32071
rect 86674 31891 86730 31947
rect 86798 31891 86854 31947
rect 86922 31891 86978 31947
rect 87046 31891 87102 31947
rect 86674 31767 86730 31823
rect 86798 31767 86854 31823
rect 86922 31767 86978 31823
rect 87046 31767 87102 31823
rect 86674 31643 86730 31699
rect 86798 31643 86854 31699
rect 86922 31643 86978 31699
rect 87046 31643 87102 31699
rect 86674 31519 86730 31575
rect 86798 31519 86854 31575
rect 86922 31519 86978 31575
rect 87046 31519 87102 31575
rect 86674 31395 86730 31451
rect 86798 31395 86854 31451
rect 86922 31395 86978 31451
rect 87046 31395 87102 31451
rect 86674 31271 86730 31327
rect 86798 31271 86854 31327
rect 86922 31271 86978 31327
rect 87046 31271 87102 31327
rect 86674 31147 86730 31203
rect 86798 31147 86854 31203
rect 86922 31147 86978 31203
rect 87046 31147 87102 31203
rect 86674 31023 86730 31079
rect 86798 31023 86854 31079
rect 86922 31023 86978 31079
rect 87046 31023 87102 31079
rect 86674 30899 86730 30955
rect 86798 30899 86854 30955
rect 86922 30899 86978 30955
rect 87046 30899 87102 30955
rect 86674 30775 86730 30831
rect 86798 30775 86854 30831
rect 86922 30775 86978 30831
rect 87046 30775 87102 30831
rect 86674 30651 86730 30707
rect 86798 30651 86854 30707
rect 86922 30651 86978 30707
rect 87046 30651 87102 30707
rect 86674 30527 86730 30583
rect 86798 30527 86854 30583
rect 86922 30527 86978 30583
rect 87046 30527 87102 30583
rect 86674 30403 86730 30459
rect 86798 30403 86854 30459
rect 86922 30403 86978 30459
rect 87046 30403 87102 30459
rect 86674 30279 86730 30335
rect 86798 30279 86854 30335
rect 86922 30279 86978 30335
rect 87046 30279 87102 30335
rect 86674 30155 86730 30211
rect 86798 30155 86854 30211
rect 86922 30155 86978 30211
rect 87046 30155 87102 30211
rect 86674 30031 86730 30087
rect 86798 30031 86854 30087
rect 86922 30031 86978 30087
rect 87046 30031 87102 30087
rect 86674 29907 86730 29963
rect 86798 29907 86854 29963
rect 86922 29907 86978 29963
rect 87046 29907 87102 29963
rect 86550 26200 86606 26256
rect 86550 26076 86606 26132
rect 86550 25952 86606 26008
rect 86550 25828 86606 25884
rect 86550 25704 86606 25760
rect 86550 25580 86606 25636
rect 86550 25456 86606 25512
rect 86550 25332 86606 25388
rect 86674 26200 86730 26256
rect 86798 26200 86854 26256
rect 86922 26200 86978 26256
rect 87046 26200 87102 26256
rect 86674 26076 86730 26132
rect 86798 26076 86854 26132
rect 86922 26076 86978 26132
rect 87046 26076 87102 26132
rect 86674 25952 86730 26008
rect 86798 25952 86854 26008
rect 86922 25952 86978 26008
rect 87046 25952 87102 26008
rect 86674 25828 86730 25884
rect 86798 25828 86854 25884
rect 86922 25828 86978 25884
rect 87046 25828 87102 25884
rect 86674 25704 86730 25760
rect 86798 25704 86854 25760
rect 86922 25704 86978 25760
rect 87046 25704 87102 25760
rect 86674 25580 86730 25636
rect 86798 25580 86854 25636
rect 86922 25580 86978 25636
rect 87046 25580 87102 25636
rect 86674 25456 86730 25512
rect 86798 25456 86854 25512
rect 86922 25456 86978 25512
rect 87046 25456 87102 25512
rect 86674 25332 86730 25388
rect 86798 25332 86854 25388
rect 86922 25332 86978 25388
rect 87046 25332 87102 25388
rect 1068 24544 1124 24600
rect 1068 24420 1124 24476
rect 1068 24296 1124 24352
rect 1068 24172 1124 24228
rect 1068 24048 1124 24104
rect 1068 23924 1124 23980
rect 1068 23800 1124 23856
rect 1068 23676 1124 23732
rect 1192 24544 1248 24600
rect 1316 24544 1372 24600
rect 1440 24544 1496 24600
rect 1564 24544 1620 24600
rect 1192 24420 1248 24476
rect 1316 24420 1372 24476
rect 1440 24420 1496 24476
rect 1564 24420 1620 24476
rect 1192 24296 1248 24352
rect 1316 24296 1372 24352
rect 1440 24296 1496 24352
rect 1564 24296 1620 24352
rect 1192 24172 1248 24228
rect 1316 24172 1372 24228
rect 1440 24172 1496 24228
rect 1564 24172 1620 24228
rect 1192 24048 1248 24104
rect 1316 24048 1372 24104
rect 1440 24048 1496 24104
rect 1564 24048 1620 24104
rect 1192 23924 1248 23980
rect 1316 23924 1372 23980
rect 1440 23924 1496 23980
rect 1564 23924 1620 23980
rect 1192 23800 1248 23856
rect 1316 23800 1372 23856
rect 1440 23800 1496 23856
rect 1564 23800 1620 23856
rect 1192 23676 1248 23732
rect 1316 23676 1372 23732
rect 1440 23676 1496 23732
rect 1564 23676 1620 23732
rect 85750 24544 85806 24600
rect 85750 24420 85806 24476
rect 85750 24296 85806 24352
rect 85750 24172 85806 24228
rect 85750 24048 85806 24104
rect 85750 23924 85806 23980
rect 85750 23800 85806 23856
rect 85750 23676 85806 23732
rect 85874 24544 85930 24600
rect 85998 24544 86054 24600
rect 86122 24544 86178 24600
rect 86246 24544 86302 24600
rect 85874 24420 85930 24476
rect 85998 24420 86054 24476
rect 86122 24420 86178 24476
rect 86246 24420 86302 24476
rect 85874 24296 85930 24352
rect 85998 24296 86054 24352
rect 86122 24296 86178 24352
rect 86246 24296 86302 24352
rect 85874 24172 85930 24228
rect 85998 24172 86054 24228
rect 86122 24172 86178 24228
rect 86246 24172 86302 24228
rect 85874 24048 85930 24104
rect 85998 24048 86054 24104
rect 86122 24048 86178 24104
rect 86246 24048 86302 24104
rect 85874 23924 85930 23980
rect 85998 23924 86054 23980
rect 86122 23924 86178 23980
rect 86246 23924 86302 23980
rect 85874 23800 85930 23856
rect 85998 23800 86054 23856
rect 86122 23800 86178 23856
rect 86246 23800 86302 23856
rect 85874 23676 85930 23732
rect 85998 23676 86054 23732
rect 86122 23676 86178 23732
rect 86246 23676 86302 23732
rect 1930 12958 1986 13014
rect 2054 12958 2110 13014
rect 2178 12958 2234 13014
rect 2302 12958 2358 13014
rect 1930 12834 1986 12890
rect 2054 12834 2110 12890
rect 2178 12834 2234 12890
rect 2302 12834 2358 12890
rect 1930 12710 1986 12766
rect 2054 12710 2110 12766
rect 2178 12710 2234 12766
rect 2302 12710 2358 12766
rect 1930 12586 1986 12642
rect 2054 12586 2110 12642
rect 2178 12586 2234 12642
rect 2302 12586 2358 12642
rect 86612 12803 86668 12859
rect 86736 12803 86792 12859
rect 86860 12803 86916 12859
rect 86984 12803 87040 12859
rect 86612 12679 86668 12735
rect 86736 12679 86792 12735
rect 86860 12679 86916 12735
rect 86984 12679 87040 12735
rect 86612 12555 86668 12611
rect 86736 12555 86792 12611
rect 86860 12555 86916 12611
rect 86984 12555 87040 12611
rect 86612 12431 86668 12487
rect 86736 12431 86792 12487
rect 86860 12431 86916 12487
rect 86984 12431 87040 12487
rect 1130 11608 1186 11664
rect 1254 11608 1310 11664
rect 1378 11608 1434 11664
rect 1502 11608 1558 11664
rect 1130 11484 1186 11540
rect 1254 11484 1310 11540
rect 1378 11484 1434 11540
rect 1502 11484 1558 11540
rect 1130 11360 1186 11416
rect 1254 11360 1310 11416
rect 1378 11360 1434 11416
rect 1502 11360 1558 11416
rect 1130 11236 1186 11292
rect 1254 11236 1310 11292
rect 1378 11236 1434 11292
rect 1502 11236 1558 11292
rect 85812 11608 85868 11664
rect 85936 11608 85992 11664
rect 86060 11608 86116 11664
rect 86184 11608 86240 11664
rect 85812 11484 85868 11540
rect 85936 11484 85992 11540
rect 86060 11484 86116 11540
rect 86184 11484 86240 11540
rect 85812 11360 85868 11416
rect 85936 11360 85992 11416
rect 86060 11360 86116 11416
rect 86184 11360 86240 11416
rect 85812 11236 85868 11292
rect 85936 11236 85992 11292
rect 86060 11236 86116 11292
rect 86184 11236 86240 11292
rect 86612 10708 86668 10764
rect 86736 10708 86792 10764
rect 86860 10708 86916 10764
rect 86984 10708 87040 10764
rect 1930 10584 1986 10640
rect 2054 10584 2110 10640
rect 2178 10584 2234 10640
rect 2302 10584 2358 10640
rect 1930 10460 1986 10516
rect 2054 10460 2110 10516
rect 2178 10460 2234 10516
rect 2302 10460 2358 10516
rect 86612 10584 86668 10640
rect 86736 10584 86792 10640
rect 86860 10584 86916 10640
rect 86984 10584 87040 10640
rect 86612 10460 86668 10516
rect 86736 10460 86792 10516
rect 86860 10460 86916 10516
rect 86984 10460 87040 10516
rect 86612 10336 86668 10392
rect 86736 10336 86792 10392
rect 86860 10336 86916 10392
rect 86984 10336 87040 10392
rect 1130 9808 1186 9864
rect 1254 9808 1310 9864
rect 1378 9808 1434 9864
rect 1502 9808 1558 9864
rect 1130 9684 1186 9740
rect 1254 9684 1310 9740
rect 1378 9684 1434 9740
rect 1502 9684 1558 9740
rect 1130 9560 1186 9616
rect 1254 9560 1310 9616
rect 1378 9560 1434 9616
rect 1502 9560 1558 9616
rect 1130 9436 1186 9492
rect 1254 9436 1310 9492
rect 1378 9436 1434 9492
rect 1502 9436 1558 9492
rect 85812 9808 85868 9864
rect 85936 9808 85992 9864
rect 86060 9808 86116 9864
rect 86184 9808 86240 9864
rect 85812 9684 85868 9740
rect 85936 9684 85992 9740
rect 86060 9684 86116 9740
rect 86184 9684 86240 9740
rect 85812 9560 85868 9616
rect 85936 9560 85992 9616
rect 86060 9560 86116 9616
rect 86184 9560 86240 9616
rect 85812 9436 85868 9492
rect 85936 9436 85992 9492
rect 86060 9436 86116 9492
rect 86184 9436 86240 9492
rect 86612 8908 86668 8964
rect 86736 8908 86792 8964
rect 86860 8908 86916 8964
rect 86984 8908 87040 8964
rect 1930 8784 1986 8840
rect 2054 8784 2110 8840
rect 2178 8784 2234 8840
rect 2302 8784 2358 8840
rect 1930 8660 1986 8716
rect 2054 8660 2110 8716
rect 2178 8660 2234 8716
rect 2302 8660 2358 8716
rect 86612 8784 86668 8840
rect 86736 8784 86792 8840
rect 86860 8784 86916 8840
rect 86984 8784 87040 8840
rect 86612 8660 86668 8716
rect 86736 8660 86792 8716
rect 86860 8660 86916 8716
rect 86984 8660 87040 8716
rect 86612 8536 86668 8592
rect 86736 8536 86792 8592
rect 86860 8536 86916 8592
rect 86984 8536 87040 8592
rect 1130 8008 1186 8064
rect 1254 8008 1310 8064
rect 1378 8008 1434 8064
rect 1502 8008 1558 8064
rect 1130 7884 1186 7940
rect 1254 7884 1310 7940
rect 1378 7884 1434 7940
rect 1502 7884 1558 7940
rect 1130 7760 1186 7816
rect 1254 7760 1310 7816
rect 1378 7760 1434 7816
rect 1502 7760 1558 7816
rect 1130 7636 1186 7692
rect 1254 7636 1310 7692
rect 1378 7636 1434 7692
rect 1502 7636 1558 7692
rect 85812 8008 85868 8064
rect 85936 8008 85992 8064
rect 86060 8008 86116 8064
rect 86184 8008 86240 8064
rect 85812 7884 85868 7940
rect 85936 7884 85992 7940
rect 86060 7884 86116 7940
rect 86184 7884 86240 7940
rect 85812 7760 85868 7816
rect 85936 7760 85992 7816
rect 86060 7760 86116 7816
rect 86184 7760 86240 7816
rect 85812 7636 85868 7692
rect 85936 7636 85992 7692
rect 86060 7636 86116 7692
rect 86184 7636 86240 7692
rect 86612 7108 86668 7164
rect 86736 7108 86792 7164
rect 86860 7108 86916 7164
rect 86984 7108 87040 7164
rect 1930 6984 1986 7040
rect 2054 6984 2110 7040
rect 2178 6984 2234 7040
rect 2302 6984 2358 7040
rect 1930 6860 1986 6916
rect 2054 6860 2110 6916
rect 2178 6860 2234 6916
rect 2302 6860 2358 6916
rect 86612 6984 86668 7040
rect 86736 6984 86792 7040
rect 86860 6984 86916 7040
rect 86984 6984 87040 7040
rect 86612 6860 86668 6916
rect 86736 6860 86792 6916
rect 86860 6860 86916 6916
rect 86984 6860 87040 6916
rect 86612 6736 86668 6792
rect 86736 6736 86792 6792
rect 86860 6736 86916 6792
rect 86984 6736 87040 6792
rect 1130 6208 1186 6264
rect 1254 6208 1310 6264
rect 1378 6208 1434 6264
rect 1502 6208 1558 6264
rect 1130 6084 1186 6140
rect 1254 6084 1310 6140
rect 1378 6084 1434 6140
rect 1502 6084 1558 6140
rect 1130 5960 1186 6016
rect 1254 5960 1310 6016
rect 1378 5960 1434 6016
rect 1502 5960 1558 6016
rect 1130 5836 1186 5892
rect 1254 5836 1310 5892
rect 1378 5836 1434 5892
rect 1502 5836 1558 5892
rect 85812 6208 85868 6264
rect 85936 6208 85992 6264
rect 86060 6208 86116 6264
rect 86184 6208 86240 6264
rect 85812 6084 85868 6140
rect 85936 6084 85992 6140
rect 86060 6084 86116 6140
rect 86184 6084 86240 6140
rect 85812 5960 85868 6016
rect 85936 5960 85992 6016
rect 86060 5960 86116 6016
rect 86184 5960 86240 6016
rect 85812 5836 85868 5892
rect 85936 5836 85992 5892
rect 86060 5836 86116 5892
rect 86184 5836 86240 5892
rect 86612 5308 86668 5364
rect 86736 5308 86792 5364
rect 86860 5308 86916 5364
rect 86984 5308 87040 5364
rect 1930 5184 1986 5240
rect 2054 5184 2110 5240
rect 2178 5184 2234 5240
rect 2302 5184 2358 5240
rect 1930 5060 1986 5116
rect 2054 5060 2110 5116
rect 2178 5060 2234 5116
rect 2302 5060 2358 5116
rect 86612 5184 86668 5240
rect 86736 5184 86792 5240
rect 86860 5184 86916 5240
rect 86984 5184 87040 5240
rect 86612 5060 86668 5116
rect 86736 5060 86792 5116
rect 86860 5060 86916 5116
rect 86984 5060 87040 5116
rect 86612 4936 86668 4992
rect 86736 4936 86792 4992
rect 86860 4936 86916 4992
rect 86984 4936 87040 4992
rect 1130 4408 1186 4464
rect 1254 4408 1310 4464
rect 1378 4408 1434 4464
rect 1502 4408 1558 4464
rect 1130 4284 1186 4340
rect 1254 4284 1310 4340
rect 1378 4284 1434 4340
rect 1502 4284 1558 4340
rect 1130 4160 1186 4216
rect 1254 4160 1310 4216
rect 1378 4160 1434 4216
rect 1502 4160 1558 4216
rect 1130 4036 1186 4092
rect 1254 4036 1310 4092
rect 1378 4036 1434 4092
rect 1502 4036 1558 4092
rect 85812 4408 85868 4464
rect 85936 4408 85992 4464
rect 86060 4408 86116 4464
rect 86184 4408 86240 4464
rect 85812 4284 85868 4340
rect 85936 4284 85992 4340
rect 86060 4284 86116 4340
rect 86184 4284 86240 4340
rect 85812 4160 85868 4216
rect 85936 4160 85992 4216
rect 86060 4160 86116 4216
rect 86184 4160 86240 4216
rect 85812 4036 85868 4092
rect 85936 4036 85992 4092
rect 86060 4036 86116 4092
rect 86184 4036 86240 4092
rect 86612 3576 86668 3632
rect 86736 3576 86792 3632
rect 86860 3576 86916 3632
rect 86984 3576 87040 3632
rect 1930 3384 1986 3440
rect 2054 3384 2110 3440
rect 2178 3384 2234 3440
rect 2302 3384 2358 3440
rect 1930 3260 1986 3316
rect 2054 3260 2110 3316
rect 2178 3260 2234 3316
rect 2302 3260 2358 3316
rect 86612 3452 86668 3508
rect 86736 3452 86792 3508
rect 86860 3452 86916 3508
rect 86984 3452 87040 3508
rect 86612 3328 86668 3384
rect 86736 3328 86792 3384
rect 86860 3328 86916 3384
rect 86984 3328 87040 3384
rect 86612 3204 86668 3260
rect 86736 3204 86792 3260
rect 86860 3204 86916 3260
rect 86984 3204 87040 3260
<< metal4 >>
rect 1044 45436 1644 45472
rect 1044 45380 1130 45436
rect 1186 45380 1254 45436
rect 1310 45380 1378 45436
rect 1434 45380 1502 45436
rect 1558 45380 1644 45436
rect 1044 35489 1644 45380
rect 1044 35433 1068 35489
rect 1124 35433 1192 35489
rect 1248 35433 1316 35489
rect 1372 35433 1440 35489
rect 1496 35433 1564 35489
rect 1620 35433 1644 35489
rect 1044 35365 1644 35433
rect 1044 35309 1068 35365
rect 1124 35309 1192 35365
rect 1248 35309 1316 35365
rect 1372 35309 1440 35365
rect 1496 35309 1564 35365
rect 1620 35309 1644 35365
rect 1044 35241 1644 35309
rect 1044 35185 1068 35241
rect 1124 35185 1192 35241
rect 1248 35185 1316 35241
rect 1372 35185 1440 35241
rect 1496 35185 1564 35241
rect 1620 35185 1644 35241
rect 1044 35117 1644 35185
rect 1044 35061 1068 35117
rect 1124 35061 1192 35117
rect 1248 35061 1316 35117
rect 1372 35061 1440 35117
rect 1496 35061 1564 35117
rect 1620 35061 1644 35117
rect 1044 34993 1644 35061
rect 1044 34937 1068 34993
rect 1124 34937 1192 34993
rect 1248 34937 1316 34993
rect 1372 34937 1440 34993
rect 1496 34937 1564 34993
rect 1620 34937 1644 34993
rect 1044 34869 1644 34937
rect 1044 34813 1068 34869
rect 1124 34813 1192 34869
rect 1248 34813 1316 34869
rect 1372 34813 1440 34869
rect 1496 34813 1564 34869
rect 1620 34813 1644 34869
rect 1044 34745 1644 34813
rect 1044 34689 1068 34745
rect 1124 34689 1192 34745
rect 1248 34689 1316 34745
rect 1372 34689 1440 34745
rect 1496 34689 1564 34745
rect 1620 34689 1644 34745
rect 1044 34621 1644 34689
rect 1044 34565 1068 34621
rect 1124 34565 1192 34621
rect 1248 34565 1316 34621
rect 1372 34565 1440 34621
rect 1496 34565 1564 34621
rect 1620 34565 1644 34621
rect 1044 34497 1644 34565
rect 1044 34441 1068 34497
rect 1124 34441 1192 34497
rect 1248 34441 1316 34497
rect 1372 34441 1440 34497
rect 1496 34441 1564 34497
rect 1620 34441 1644 34497
rect 1044 34373 1644 34441
rect 1044 34317 1068 34373
rect 1124 34317 1192 34373
rect 1248 34317 1316 34373
rect 1372 34317 1440 34373
rect 1496 34317 1564 34373
rect 1620 34317 1644 34373
rect 1044 34249 1644 34317
rect 1044 34193 1068 34249
rect 1124 34193 1192 34249
rect 1248 34193 1316 34249
rect 1372 34193 1440 34249
rect 1496 34193 1564 34249
rect 1620 34193 1644 34249
rect 1044 34125 1644 34193
rect 1044 34069 1068 34125
rect 1124 34069 1192 34125
rect 1248 34069 1316 34125
rect 1372 34069 1440 34125
rect 1496 34069 1564 34125
rect 1620 34069 1644 34125
rect 1044 34001 1644 34069
rect 1044 33945 1068 34001
rect 1124 33945 1192 34001
rect 1248 33945 1316 34001
rect 1372 33945 1440 34001
rect 1496 33945 1564 34001
rect 1620 33945 1644 34001
rect 1044 33877 1644 33945
rect 1044 33821 1068 33877
rect 1124 33821 1192 33877
rect 1248 33821 1316 33877
rect 1372 33821 1440 33877
rect 1496 33821 1564 33877
rect 1620 33821 1644 33877
rect 1044 33753 1644 33821
rect 1044 33697 1068 33753
rect 1124 33697 1192 33753
rect 1248 33697 1316 33753
rect 1372 33697 1440 33753
rect 1496 33697 1564 33753
rect 1620 33697 1644 33753
rect 1044 33629 1644 33697
rect 1044 33573 1068 33629
rect 1124 33573 1192 33629
rect 1248 33573 1316 33629
rect 1372 33573 1440 33629
rect 1496 33573 1564 33629
rect 1620 33573 1644 33629
rect 1044 33505 1644 33573
rect 1044 33449 1068 33505
rect 1124 33449 1192 33505
rect 1248 33449 1316 33505
rect 1372 33449 1440 33505
rect 1496 33449 1564 33505
rect 1620 33449 1644 33505
rect 1044 24600 1644 33449
rect 1044 24544 1068 24600
rect 1124 24544 1192 24600
rect 1248 24544 1316 24600
rect 1372 24544 1440 24600
rect 1496 24544 1564 24600
rect 1620 24544 1644 24600
rect 1044 24476 1644 24544
rect 1044 24420 1068 24476
rect 1124 24420 1192 24476
rect 1248 24420 1316 24476
rect 1372 24420 1440 24476
rect 1496 24420 1564 24476
rect 1620 24420 1644 24476
rect 1044 24352 1644 24420
rect 1044 24296 1068 24352
rect 1124 24296 1192 24352
rect 1248 24296 1316 24352
rect 1372 24296 1440 24352
rect 1496 24296 1564 24352
rect 1620 24296 1644 24352
rect 1044 24228 1644 24296
rect 1044 24172 1068 24228
rect 1124 24172 1192 24228
rect 1248 24172 1316 24228
rect 1372 24172 1440 24228
rect 1496 24172 1564 24228
rect 1620 24172 1644 24228
rect 1044 24104 1644 24172
rect 1044 24048 1068 24104
rect 1124 24048 1192 24104
rect 1248 24048 1316 24104
rect 1372 24048 1440 24104
rect 1496 24048 1564 24104
rect 1620 24048 1644 24104
rect 1044 23980 1644 24048
rect 1044 23924 1068 23980
rect 1124 23924 1192 23980
rect 1248 23924 1316 23980
rect 1372 23924 1440 23980
rect 1496 23924 1564 23980
rect 1620 23924 1644 23980
rect 1044 23856 1644 23924
rect 1044 23800 1068 23856
rect 1124 23800 1192 23856
rect 1248 23800 1316 23856
rect 1372 23800 1440 23856
rect 1496 23800 1564 23856
rect 1620 23800 1644 23856
rect 1044 23732 1644 23800
rect 1044 23676 1068 23732
rect 1124 23676 1192 23732
rect 1248 23676 1316 23732
rect 1372 23676 1440 23732
rect 1496 23676 1564 23732
rect 1620 23676 1644 23732
rect 1044 11664 1644 23676
rect 1044 11608 1130 11664
rect 1186 11608 1254 11664
rect 1310 11608 1378 11664
rect 1434 11608 1502 11664
rect 1558 11608 1644 11664
rect 1044 11540 1644 11608
rect 1044 11484 1130 11540
rect 1186 11484 1254 11540
rect 1310 11484 1378 11540
rect 1434 11484 1502 11540
rect 1558 11484 1644 11540
rect 1044 11416 1644 11484
rect 1044 11360 1130 11416
rect 1186 11360 1254 11416
rect 1310 11360 1378 11416
rect 1434 11360 1502 11416
rect 1558 11360 1644 11416
rect 1044 11292 1644 11360
rect 1044 11236 1130 11292
rect 1186 11236 1254 11292
rect 1310 11236 1378 11292
rect 1434 11236 1502 11292
rect 1558 11236 1644 11292
rect 1044 9864 1644 11236
rect 1044 9808 1130 9864
rect 1186 9808 1254 9864
rect 1310 9808 1378 9864
rect 1434 9808 1502 9864
rect 1558 9808 1644 9864
rect 1044 9740 1644 9808
rect 1044 9684 1130 9740
rect 1186 9684 1254 9740
rect 1310 9684 1378 9740
rect 1434 9684 1502 9740
rect 1558 9684 1644 9740
rect 1044 9616 1644 9684
rect 1044 9560 1130 9616
rect 1186 9560 1254 9616
rect 1310 9560 1378 9616
rect 1434 9560 1502 9616
rect 1558 9560 1644 9616
rect 1044 9492 1644 9560
rect 1044 9436 1130 9492
rect 1186 9436 1254 9492
rect 1310 9436 1378 9492
rect 1434 9436 1502 9492
rect 1558 9436 1644 9492
rect 1044 8064 1644 9436
rect 1044 8008 1130 8064
rect 1186 8008 1254 8064
rect 1310 8008 1378 8064
rect 1434 8008 1502 8064
rect 1558 8008 1644 8064
rect 1044 7940 1644 8008
rect 1044 7884 1130 7940
rect 1186 7884 1254 7940
rect 1310 7884 1378 7940
rect 1434 7884 1502 7940
rect 1558 7884 1644 7940
rect 1044 7816 1644 7884
rect 1044 7760 1130 7816
rect 1186 7760 1254 7816
rect 1310 7760 1378 7816
rect 1434 7760 1502 7816
rect 1558 7760 1644 7816
rect 1044 7692 1644 7760
rect 1044 7636 1130 7692
rect 1186 7636 1254 7692
rect 1310 7636 1378 7692
rect 1434 7636 1502 7692
rect 1558 7636 1644 7692
rect 1044 6264 1644 7636
rect 1044 6208 1130 6264
rect 1186 6208 1254 6264
rect 1310 6208 1378 6264
rect 1434 6208 1502 6264
rect 1558 6208 1644 6264
rect 1044 6140 1644 6208
rect 1044 6084 1130 6140
rect 1186 6084 1254 6140
rect 1310 6084 1378 6140
rect 1434 6084 1502 6140
rect 1558 6084 1644 6140
rect 1044 6016 1644 6084
rect 1044 5960 1130 6016
rect 1186 5960 1254 6016
rect 1310 5960 1378 6016
rect 1434 5960 1502 6016
rect 1558 5960 1644 6016
rect 1044 5892 1644 5960
rect 1044 5836 1130 5892
rect 1186 5836 1254 5892
rect 1310 5836 1378 5892
rect 1434 5836 1502 5892
rect 1558 5836 1644 5892
rect 1044 4464 1644 5836
rect 1044 4408 1130 4464
rect 1186 4408 1254 4464
rect 1310 4408 1378 4464
rect 1434 4408 1502 4464
rect 1558 4408 1644 4464
rect 1044 4340 1644 4408
rect 1044 4284 1130 4340
rect 1186 4284 1254 4340
rect 1310 4284 1378 4340
rect 1434 4284 1502 4340
rect 1558 4284 1644 4340
rect 1044 4216 1644 4284
rect 1044 4160 1130 4216
rect 1186 4160 1254 4216
rect 1310 4160 1378 4216
rect 1434 4160 1502 4216
rect 1558 4160 1644 4216
rect 1044 4092 1644 4160
rect 1044 4036 1130 4092
rect 1186 4036 1254 4092
rect 1310 4036 1378 4092
rect 1434 4036 1502 4092
rect 1558 4036 1644 4092
rect 1044 3136 1644 4036
rect 1844 45025 2444 45472
rect 1844 44969 1901 45025
rect 1957 44969 2444 45025
rect 1844 44901 2444 44969
rect 1844 44845 1901 44901
rect 1957 44845 2444 44901
rect 1844 44777 2444 44845
rect 1844 44721 1901 44777
rect 1957 44721 2444 44777
rect 1844 44653 2444 44721
rect 1844 44597 1901 44653
rect 1957 44597 2444 44653
rect 1844 44529 2444 44597
rect 1844 44473 1901 44529
rect 1957 44473 2444 44529
rect 1844 44405 2444 44473
rect 1844 44349 1901 44405
rect 1957 44349 2444 44405
rect 1844 44281 2444 44349
rect 1844 44225 1901 44281
rect 1957 44225 2444 44281
rect 1844 44157 2444 44225
rect 1844 44101 1901 44157
rect 1957 44101 2444 44157
rect 1844 44033 2444 44101
rect 1844 43977 1901 44033
rect 1957 43977 2444 44033
rect 1844 43909 2444 43977
rect 1844 43853 1901 43909
rect 1957 43853 2444 43909
rect 1844 40501 2444 43853
rect 1844 40445 1930 40501
rect 1986 40445 2054 40501
rect 2110 40445 2178 40501
rect 2234 40445 2302 40501
rect 2358 40445 2444 40501
rect 1844 40377 2444 40445
rect 1844 40321 1930 40377
rect 1986 40321 2054 40377
rect 2110 40321 2178 40377
rect 2234 40321 2302 40377
rect 2358 40321 2444 40377
rect 1844 40253 2444 40321
rect 1844 40197 1930 40253
rect 1986 40197 2054 40253
rect 2110 40197 2178 40253
rect 2234 40197 2302 40253
rect 2358 40197 2444 40253
rect 1844 40129 2444 40197
rect 1844 40073 1930 40129
rect 1986 40073 2054 40129
rect 2110 40073 2178 40129
rect 2234 40073 2302 40129
rect 2358 40073 2444 40129
rect 1844 33187 2444 40073
rect 1844 33131 1868 33187
rect 1924 33131 1992 33187
rect 2048 33131 2116 33187
rect 2172 33131 2240 33187
rect 2296 33131 2364 33187
rect 2420 33131 2444 33187
rect 1844 33063 2444 33131
rect 1844 33007 1868 33063
rect 1924 33007 1992 33063
rect 2048 33007 2116 33063
rect 2172 33007 2240 33063
rect 2296 33007 2364 33063
rect 2420 33007 2444 33063
rect 1844 32939 2444 33007
rect 1844 32883 1868 32939
rect 1924 32883 1992 32939
rect 2048 32883 2116 32939
rect 2172 32883 2240 32939
rect 2296 32883 2364 32939
rect 2420 32883 2444 32939
rect 1844 32815 2444 32883
rect 1844 32759 1868 32815
rect 1924 32759 1992 32815
rect 2048 32759 2116 32815
rect 2172 32759 2240 32815
rect 2296 32759 2364 32815
rect 2420 32759 2444 32815
rect 1844 32691 2444 32759
rect 1844 32635 1868 32691
rect 1924 32635 1992 32691
rect 2048 32635 2116 32691
rect 2172 32635 2240 32691
rect 2296 32635 2364 32691
rect 2420 32635 2444 32691
rect 1844 32567 2444 32635
rect 1844 32511 1868 32567
rect 1924 32511 1992 32567
rect 2048 32511 2116 32567
rect 2172 32511 2240 32567
rect 2296 32511 2364 32567
rect 2420 32511 2444 32567
rect 1844 32443 2444 32511
rect 1844 32387 1868 32443
rect 1924 32387 1992 32443
rect 2048 32387 2116 32443
rect 2172 32387 2240 32443
rect 2296 32387 2364 32443
rect 2420 32387 2444 32443
rect 1844 32319 2444 32387
rect 1844 32263 1868 32319
rect 1924 32263 1992 32319
rect 2048 32263 2116 32319
rect 2172 32263 2240 32319
rect 2296 32263 2364 32319
rect 2420 32263 2444 32319
rect 1844 32195 2444 32263
rect 1844 32139 1868 32195
rect 1924 32139 1992 32195
rect 2048 32139 2116 32195
rect 2172 32139 2240 32195
rect 2296 32139 2364 32195
rect 2420 32139 2444 32195
rect 1844 32071 2444 32139
rect 1844 32015 1868 32071
rect 1924 32015 1992 32071
rect 2048 32015 2116 32071
rect 2172 32015 2240 32071
rect 2296 32015 2364 32071
rect 2420 32015 2444 32071
rect 1844 31947 2444 32015
rect 1844 31891 1868 31947
rect 1924 31891 1992 31947
rect 2048 31891 2116 31947
rect 2172 31891 2240 31947
rect 2296 31891 2364 31947
rect 2420 31891 2444 31947
rect 1844 31823 2444 31891
rect 1844 31767 1868 31823
rect 1924 31767 1992 31823
rect 2048 31767 2116 31823
rect 2172 31767 2240 31823
rect 2296 31767 2364 31823
rect 2420 31767 2444 31823
rect 1844 31699 2444 31767
rect 1844 31643 1868 31699
rect 1924 31643 1992 31699
rect 2048 31643 2116 31699
rect 2172 31643 2240 31699
rect 2296 31643 2364 31699
rect 2420 31643 2444 31699
rect 1844 31575 2444 31643
rect 1844 31519 1868 31575
rect 1924 31519 1992 31575
rect 2048 31519 2116 31575
rect 2172 31519 2240 31575
rect 2296 31519 2364 31575
rect 2420 31519 2444 31575
rect 1844 31451 2444 31519
rect 1844 31395 1868 31451
rect 1924 31395 1992 31451
rect 2048 31395 2116 31451
rect 2172 31395 2240 31451
rect 2296 31395 2364 31451
rect 2420 31395 2444 31451
rect 1844 31327 2444 31395
rect 1844 31271 1868 31327
rect 1924 31271 1992 31327
rect 2048 31271 2116 31327
rect 2172 31271 2240 31327
rect 2296 31271 2364 31327
rect 2420 31271 2444 31327
rect 1844 31203 2444 31271
rect 1844 31147 1868 31203
rect 1924 31147 1992 31203
rect 2048 31147 2116 31203
rect 2172 31147 2240 31203
rect 2296 31147 2364 31203
rect 2420 31147 2444 31203
rect 1844 31079 2444 31147
rect 1844 31023 1868 31079
rect 1924 31023 1992 31079
rect 2048 31023 2116 31079
rect 2172 31023 2240 31079
rect 2296 31023 2364 31079
rect 2420 31023 2444 31079
rect 1844 30955 2444 31023
rect 1844 30899 1868 30955
rect 1924 30899 1992 30955
rect 2048 30899 2116 30955
rect 2172 30899 2240 30955
rect 2296 30899 2364 30955
rect 2420 30899 2444 30955
rect 1844 30831 2444 30899
rect 1844 30775 1868 30831
rect 1924 30775 1992 30831
rect 2048 30775 2116 30831
rect 2172 30775 2240 30831
rect 2296 30775 2364 30831
rect 2420 30775 2444 30831
rect 1844 30707 2444 30775
rect 1844 30651 1868 30707
rect 1924 30651 1992 30707
rect 2048 30651 2116 30707
rect 2172 30651 2240 30707
rect 2296 30651 2364 30707
rect 2420 30651 2444 30707
rect 1844 30583 2444 30651
rect 1844 30527 1868 30583
rect 1924 30527 1992 30583
rect 2048 30527 2116 30583
rect 2172 30527 2240 30583
rect 2296 30527 2364 30583
rect 2420 30527 2444 30583
rect 1844 30459 2444 30527
rect 1844 30403 1868 30459
rect 1924 30403 1992 30459
rect 2048 30403 2116 30459
rect 2172 30403 2240 30459
rect 2296 30403 2364 30459
rect 2420 30403 2444 30459
rect 1844 30335 2444 30403
rect 1844 30279 1868 30335
rect 1924 30279 1992 30335
rect 2048 30279 2116 30335
rect 2172 30279 2240 30335
rect 2296 30279 2364 30335
rect 2420 30279 2444 30335
rect 1844 30211 2444 30279
rect 1844 30155 1868 30211
rect 1924 30155 1992 30211
rect 2048 30155 2116 30211
rect 2172 30155 2240 30211
rect 2296 30155 2364 30211
rect 2420 30155 2444 30211
rect 1844 30087 2444 30155
rect 1844 30031 1868 30087
rect 1924 30031 1992 30087
rect 2048 30031 2116 30087
rect 2172 30031 2240 30087
rect 2296 30031 2364 30087
rect 2420 30031 2444 30087
rect 1844 29963 2444 30031
rect 1844 29907 1868 29963
rect 1924 29907 1992 29963
rect 2048 29907 2116 29963
rect 2172 29907 2240 29963
rect 2296 29907 2364 29963
rect 2420 29907 2444 29963
rect 1844 13014 2444 29907
rect 1844 12958 1930 13014
rect 1986 12958 2054 13014
rect 2110 12958 2178 13014
rect 2234 12958 2302 13014
rect 2358 12958 2444 13014
rect 1844 12890 2444 12958
rect 1844 12834 1930 12890
rect 1986 12834 2054 12890
rect 2110 12834 2178 12890
rect 2234 12834 2302 12890
rect 2358 12834 2444 12890
rect 1844 12766 2444 12834
rect 1844 12710 1930 12766
rect 1986 12710 2054 12766
rect 2110 12710 2178 12766
rect 2234 12710 2302 12766
rect 2358 12710 2444 12766
rect 1844 12642 2444 12710
rect 1844 12586 1930 12642
rect 1986 12586 2054 12642
rect 2110 12586 2178 12642
rect 2234 12586 2302 12642
rect 2358 12586 2444 12642
rect 1844 10640 2444 12586
rect 1844 10584 1930 10640
rect 1986 10584 2054 10640
rect 2110 10584 2178 10640
rect 2234 10584 2302 10640
rect 2358 10584 2444 10640
rect 1844 10516 2444 10584
rect 1844 10460 1930 10516
rect 1986 10460 2054 10516
rect 2110 10460 2178 10516
rect 2234 10460 2302 10516
rect 2358 10460 2444 10516
rect 1844 8840 2444 10460
rect 1844 8784 1930 8840
rect 1986 8784 2054 8840
rect 2110 8784 2178 8840
rect 2234 8784 2302 8840
rect 2358 8784 2444 8840
rect 1844 8716 2444 8784
rect 1844 8660 1930 8716
rect 1986 8660 2054 8716
rect 2110 8660 2178 8716
rect 2234 8660 2302 8716
rect 2358 8660 2444 8716
rect 1844 7040 2444 8660
rect 1844 6984 1930 7040
rect 1986 6984 2054 7040
rect 2110 6984 2178 7040
rect 2234 6984 2302 7040
rect 2358 6984 2444 7040
rect 1844 6916 2444 6984
rect 1844 6860 1930 6916
rect 1986 6860 2054 6916
rect 2110 6860 2178 6916
rect 2234 6860 2302 6916
rect 2358 6860 2444 6916
rect 1844 5240 2444 6860
rect 1844 5184 1930 5240
rect 1986 5184 2054 5240
rect 2110 5184 2178 5240
rect 2234 5184 2302 5240
rect 2358 5184 2444 5240
rect 1844 5116 2444 5184
rect 1844 5060 1930 5116
rect 1986 5060 2054 5116
rect 2110 5060 2178 5116
rect 2234 5060 2302 5116
rect 2358 5060 2444 5116
rect 1844 3440 2444 5060
rect 1844 3384 1930 3440
rect 1986 3384 2054 3440
rect 2110 3384 2178 3440
rect 2234 3384 2302 3440
rect 2358 3384 2444 3440
rect 1844 3316 2444 3384
rect 1844 3260 1930 3316
rect 1986 3260 2054 3316
rect 2110 3260 2178 3316
rect 2234 3260 2302 3316
rect 2358 3260 2444 3316
rect 1844 3136 2444 3260
rect 85726 45436 86326 45472
rect 85726 45380 85812 45436
rect 85868 45380 85936 45436
rect 85992 45380 86060 45436
rect 86116 45380 86184 45436
rect 86240 45380 86326 45436
rect 85726 39391 86326 45380
rect 85726 39335 85750 39391
rect 85806 39335 85874 39391
rect 85930 39335 85998 39391
rect 86054 39335 86122 39391
rect 86178 39335 86246 39391
rect 86302 39335 86326 39391
rect 85726 39267 86326 39335
rect 85726 39211 85750 39267
rect 85806 39211 85874 39267
rect 85930 39211 85998 39267
rect 86054 39211 86122 39267
rect 86178 39211 86246 39267
rect 86302 39211 86326 39267
rect 85726 39143 86326 39211
rect 85726 39087 85750 39143
rect 85806 39087 85874 39143
rect 85930 39087 85998 39143
rect 86054 39087 86122 39143
rect 86178 39087 86246 39143
rect 86302 39087 86326 39143
rect 85726 39019 86326 39087
rect 85726 38963 85750 39019
rect 85806 38963 85874 39019
rect 85930 38963 85998 39019
rect 86054 38963 86122 39019
rect 86178 38963 86246 39019
rect 86302 38963 86326 39019
rect 85726 38895 86326 38963
rect 85726 38839 85750 38895
rect 85806 38839 85874 38895
rect 85930 38839 85998 38895
rect 86054 38839 86122 38895
rect 86178 38839 86246 38895
rect 86302 38839 86326 38895
rect 85726 38771 86326 38839
rect 85726 38715 85750 38771
rect 85806 38715 85874 38771
rect 85930 38715 85998 38771
rect 86054 38715 86122 38771
rect 86178 38715 86246 38771
rect 86302 38715 86326 38771
rect 85726 38647 86326 38715
rect 85726 38591 85750 38647
rect 85806 38591 85874 38647
rect 85930 38591 85998 38647
rect 86054 38591 86122 38647
rect 86178 38591 86246 38647
rect 86302 38591 86326 38647
rect 85726 38523 86326 38591
rect 85726 38467 85750 38523
rect 85806 38467 85874 38523
rect 85930 38467 85998 38523
rect 86054 38467 86122 38523
rect 86178 38467 86246 38523
rect 86302 38467 86326 38523
rect 85726 38399 86326 38467
rect 85726 38343 85750 38399
rect 85806 38343 85874 38399
rect 85930 38343 85998 38399
rect 86054 38343 86122 38399
rect 86178 38343 86246 38399
rect 86302 38343 86326 38399
rect 85726 38275 86326 38343
rect 85726 38219 85750 38275
rect 85806 38219 85874 38275
rect 85930 38219 85998 38275
rect 86054 38219 86122 38275
rect 86178 38219 86246 38275
rect 86302 38219 86326 38275
rect 85726 38151 86326 38219
rect 85726 38095 85750 38151
rect 85806 38095 85874 38151
rect 85930 38095 85998 38151
rect 86054 38095 86122 38151
rect 86178 38095 86246 38151
rect 86302 38095 86326 38151
rect 85726 35489 86326 38095
rect 85726 35433 85750 35489
rect 85806 35433 85874 35489
rect 85930 35433 85998 35489
rect 86054 35433 86122 35489
rect 86178 35433 86246 35489
rect 86302 35433 86326 35489
rect 85726 35365 86326 35433
rect 85726 35309 85750 35365
rect 85806 35309 85874 35365
rect 85930 35309 85998 35365
rect 86054 35309 86122 35365
rect 86178 35309 86246 35365
rect 86302 35309 86326 35365
rect 85726 35241 86326 35309
rect 85726 35185 85750 35241
rect 85806 35185 85874 35241
rect 85930 35185 85998 35241
rect 86054 35185 86122 35241
rect 86178 35185 86246 35241
rect 86302 35185 86326 35241
rect 85726 35117 86326 35185
rect 85726 35061 85750 35117
rect 85806 35061 85874 35117
rect 85930 35061 85998 35117
rect 86054 35061 86122 35117
rect 86178 35061 86246 35117
rect 86302 35061 86326 35117
rect 85726 34993 86326 35061
rect 85726 34937 85750 34993
rect 85806 34937 85874 34993
rect 85930 34937 85998 34993
rect 86054 34937 86122 34993
rect 86178 34937 86246 34993
rect 86302 34937 86326 34993
rect 85726 34869 86326 34937
rect 85726 34813 85750 34869
rect 85806 34813 85874 34869
rect 85930 34813 85998 34869
rect 86054 34813 86122 34869
rect 86178 34813 86246 34869
rect 86302 34813 86326 34869
rect 85726 34745 86326 34813
rect 85726 34689 85750 34745
rect 85806 34689 85874 34745
rect 85930 34689 85998 34745
rect 86054 34689 86122 34745
rect 86178 34689 86246 34745
rect 86302 34689 86326 34745
rect 85726 34621 86326 34689
rect 85726 34565 85750 34621
rect 85806 34565 85874 34621
rect 85930 34565 85998 34621
rect 86054 34565 86122 34621
rect 86178 34565 86246 34621
rect 86302 34565 86326 34621
rect 85726 34497 86326 34565
rect 85726 34441 85750 34497
rect 85806 34441 85874 34497
rect 85930 34441 85998 34497
rect 86054 34441 86122 34497
rect 86178 34441 86246 34497
rect 86302 34441 86326 34497
rect 85726 34373 86326 34441
rect 85726 34317 85750 34373
rect 85806 34317 85874 34373
rect 85930 34317 85998 34373
rect 86054 34317 86122 34373
rect 86178 34317 86246 34373
rect 86302 34317 86326 34373
rect 85726 34249 86326 34317
rect 85726 34193 85750 34249
rect 85806 34193 85874 34249
rect 85930 34193 85998 34249
rect 86054 34193 86122 34249
rect 86178 34193 86246 34249
rect 86302 34193 86326 34249
rect 85726 34125 86326 34193
rect 85726 34069 85750 34125
rect 85806 34069 85874 34125
rect 85930 34069 85998 34125
rect 86054 34069 86122 34125
rect 86178 34069 86246 34125
rect 86302 34069 86326 34125
rect 85726 34001 86326 34069
rect 85726 33945 85750 34001
rect 85806 33945 85874 34001
rect 85930 33945 85998 34001
rect 86054 33945 86122 34001
rect 86178 33945 86246 34001
rect 86302 33945 86326 34001
rect 85726 33877 86326 33945
rect 85726 33821 85750 33877
rect 85806 33821 85874 33877
rect 85930 33821 85998 33877
rect 86054 33821 86122 33877
rect 86178 33821 86246 33877
rect 86302 33821 86326 33877
rect 85726 33753 86326 33821
rect 85726 33697 85750 33753
rect 85806 33697 85874 33753
rect 85930 33697 85998 33753
rect 86054 33697 86122 33753
rect 86178 33697 86246 33753
rect 86302 33697 86326 33753
rect 85726 33629 86326 33697
rect 85726 33573 85750 33629
rect 85806 33573 85874 33629
rect 85930 33573 85998 33629
rect 86054 33573 86122 33629
rect 86178 33573 86246 33629
rect 86302 33573 86326 33629
rect 85726 33505 86326 33573
rect 85726 33449 85750 33505
rect 85806 33449 85874 33505
rect 85930 33449 85998 33505
rect 86054 33449 86122 33505
rect 86178 33449 86246 33505
rect 86302 33449 86326 33505
rect 85726 24600 86326 33449
rect 85726 24544 85750 24600
rect 85806 24544 85874 24600
rect 85930 24544 85998 24600
rect 86054 24544 86122 24600
rect 86178 24544 86246 24600
rect 86302 24544 86326 24600
rect 85726 24476 86326 24544
rect 85726 24420 85750 24476
rect 85806 24420 85874 24476
rect 85930 24420 85998 24476
rect 86054 24420 86122 24476
rect 86178 24420 86246 24476
rect 86302 24420 86326 24476
rect 85726 24352 86326 24420
rect 85726 24296 85750 24352
rect 85806 24296 85874 24352
rect 85930 24296 85998 24352
rect 86054 24296 86122 24352
rect 86178 24296 86246 24352
rect 86302 24296 86326 24352
rect 85726 24228 86326 24296
rect 85726 24172 85750 24228
rect 85806 24172 85874 24228
rect 85930 24172 85998 24228
rect 86054 24172 86122 24228
rect 86178 24172 86246 24228
rect 86302 24172 86326 24228
rect 85726 24104 86326 24172
rect 85726 24048 85750 24104
rect 85806 24048 85874 24104
rect 85930 24048 85998 24104
rect 86054 24048 86122 24104
rect 86178 24048 86246 24104
rect 86302 24048 86326 24104
rect 85726 23980 86326 24048
rect 85726 23924 85750 23980
rect 85806 23924 85874 23980
rect 85930 23924 85998 23980
rect 86054 23924 86122 23980
rect 86178 23924 86246 23980
rect 86302 23924 86326 23980
rect 85726 23856 86326 23924
rect 85726 23800 85750 23856
rect 85806 23800 85874 23856
rect 85930 23800 85998 23856
rect 86054 23800 86122 23856
rect 86178 23800 86246 23856
rect 86302 23800 86326 23856
rect 85726 23732 86326 23800
rect 85726 23676 85750 23732
rect 85806 23676 85874 23732
rect 85930 23676 85998 23732
rect 86054 23676 86122 23732
rect 86178 23676 86246 23732
rect 86302 23676 86326 23732
rect 85726 11664 86326 23676
rect 85726 11608 85812 11664
rect 85868 11608 85936 11664
rect 85992 11608 86060 11664
rect 86116 11608 86184 11664
rect 86240 11608 86326 11664
rect 85726 11540 86326 11608
rect 85726 11484 85812 11540
rect 85868 11484 85936 11540
rect 85992 11484 86060 11540
rect 86116 11484 86184 11540
rect 86240 11484 86326 11540
rect 85726 11416 86326 11484
rect 85726 11360 85812 11416
rect 85868 11360 85936 11416
rect 85992 11360 86060 11416
rect 86116 11360 86184 11416
rect 86240 11360 86326 11416
rect 85726 11292 86326 11360
rect 85726 11236 85812 11292
rect 85868 11236 85936 11292
rect 85992 11236 86060 11292
rect 86116 11236 86184 11292
rect 86240 11236 86326 11292
rect 85726 9864 86326 11236
rect 85726 9808 85812 9864
rect 85868 9808 85936 9864
rect 85992 9808 86060 9864
rect 86116 9808 86184 9864
rect 86240 9808 86326 9864
rect 85726 9740 86326 9808
rect 85726 9684 85812 9740
rect 85868 9684 85936 9740
rect 85992 9684 86060 9740
rect 86116 9684 86184 9740
rect 86240 9684 86326 9740
rect 85726 9616 86326 9684
rect 85726 9560 85812 9616
rect 85868 9560 85936 9616
rect 85992 9560 86060 9616
rect 86116 9560 86184 9616
rect 86240 9560 86326 9616
rect 85726 9492 86326 9560
rect 85726 9436 85812 9492
rect 85868 9436 85936 9492
rect 85992 9436 86060 9492
rect 86116 9436 86184 9492
rect 86240 9436 86326 9492
rect 85726 8064 86326 9436
rect 85726 8008 85812 8064
rect 85868 8008 85936 8064
rect 85992 8008 86060 8064
rect 86116 8008 86184 8064
rect 86240 8008 86326 8064
rect 85726 7940 86326 8008
rect 85726 7884 85812 7940
rect 85868 7884 85936 7940
rect 85992 7884 86060 7940
rect 86116 7884 86184 7940
rect 86240 7884 86326 7940
rect 85726 7816 86326 7884
rect 85726 7760 85812 7816
rect 85868 7760 85936 7816
rect 85992 7760 86060 7816
rect 86116 7760 86184 7816
rect 86240 7760 86326 7816
rect 85726 7692 86326 7760
rect 85726 7636 85812 7692
rect 85868 7636 85936 7692
rect 85992 7636 86060 7692
rect 86116 7636 86184 7692
rect 86240 7636 86326 7692
rect 85726 6264 86326 7636
rect 85726 6208 85812 6264
rect 85868 6208 85936 6264
rect 85992 6208 86060 6264
rect 86116 6208 86184 6264
rect 86240 6208 86326 6264
rect 85726 6140 86326 6208
rect 85726 6084 85812 6140
rect 85868 6084 85936 6140
rect 85992 6084 86060 6140
rect 86116 6084 86184 6140
rect 86240 6084 86326 6140
rect 85726 6016 86326 6084
rect 85726 5960 85812 6016
rect 85868 5960 85936 6016
rect 85992 5960 86060 6016
rect 86116 5960 86184 6016
rect 86240 5960 86326 6016
rect 85726 5892 86326 5960
rect 85726 5836 85812 5892
rect 85868 5836 85936 5892
rect 85992 5836 86060 5892
rect 86116 5836 86184 5892
rect 86240 5836 86326 5892
rect 85726 4464 86326 5836
rect 85726 4408 85812 4464
rect 85868 4408 85936 4464
rect 85992 4408 86060 4464
rect 86116 4408 86184 4464
rect 86240 4408 86326 4464
rect 85726 4340 86326 4408
rect 85726 4284 85812 4340
rect 85868 4284 85936 4340
rect 85992 4284 86060 4340
rect 86116 4284 86184 4340
rect 86240 4284 86326 4340
rect 85726 4216 86326 4284
rect 85726 4160 85812 4216
rect 85868 4160 85936 4216
rect 85992 4160 86060 4216
rect 86116 4160 86184 4216
rect 86240 4160 86326 4216
rect 85726 4092 86326 4160
rect 85726 4036 85812 4092
rect 85868 4036 85936 4092
rect 85992 4036 86060 4092
rect 86116 4036 86184 4092
rect 86240 4036 86326 4092
rect 85726 3136 86326 4036
rect 86526 45025 87126 45472
rect 86526 44969 86550 45025
rect 86606 44969 86674 45025
rect 86730 44969 86798 45025
rect 86854 44969 86922 45025
rect 86978 44969 87046 45025
rect 87102 44969 87126 45025
rect 86526 44901 87126 44969
rect 86526 44845 86550 44901
rect 86606 44845 86674 44901
rect 86730 44845 86798 44901
rect 86854 44845 86922 44901
rect 86978 44845 87046 44901
rect 87102 44845 87126 44901
rect 86526 44777 87126 44845
rect 86526 44721 86550 44777
rect 86606 44721 86674 44777
rect 86730 44721 86798 44777
rect 86854 44721 86922 44777
rect 86978 44721 87046 44777
rect 87102 44721 87126 44777
rect 86526 44653 87126 44721
rect 86526 44597 86550 44653
rect 86606 44597 86674 44653
rect 86730 44597 86798 44653
rect 86854 44597 86922 44653
rect 86978 44597 87046 44653
rect 87102 44597 87126 44653
rect 86526 44529 87126 44597
rect 86526 44473 86550 44529
rect 86606 44473 86674 44529
rect 86730 44473 86798 44529
rect 86854 44473 86922 44529
rect 86978 44473 87046 44529
rect 87102 44473 87126 44529
rect 86526 44405 87126 44473
rect 86526 44349 86550 44405
rect 86606 44349 86674 44405
rect 86730 44349 86798 44405
rect 86854 44349 86922 44405
rect 86978 44349 87046 44405
rect 87102 44349 87126 44405
rect 86526 44281 87126 44349
rect 86526 44225 86550 44281
rect 86606 44225 86674 44281
rect 86730 44225 86798 44281
rect 86854 44225 86922 44281
rect 86978 44225 87046 44281
rect 87102 44225 87126 44281
rect 86526 44157 87126 44225
rect 86526 44101 86550 44157
rect 86606 44101 86674 44157
rect 86730 44101 86798 44157
rect 86854 44101 86922 44157
rect 86978 44101 87046 44157
rect 87102 44101 87126 44157
rect 86526 44033 87126 44101
rect 86526 43977 86550 44033
rect 86606 43977 86674 44033
rect 86730 43977 86798 44033
rect 86854 43977 86922 44033
rect 86978 43977 87046 44033
rect 87102 43977 87126 44033
rect 86526 43909 87126 43977
rect 86526 43853 86550 43909
rect 86606 43853 86674 43909
rect 86730 43853 86798 43909
rect 86854 43853 86922 43909
rect 86978 43853 87046 43909
rect 87102 43853 87126 43909
rect 86526 41791 87126 43853
rect 86526 41735 86550 41791
rect 86606 41735 86674 41791
rect 86730 41735 86798 41791
rect 86854 41735 86922 41791
rect 86978 41735 87046 41791
rect 87102 41735 87126 41791
rect 86526 41667 87126 41735
rect 86526 41611 86550 41667
rect 86606 41611 86674 41667
rect 86730 41611 86798 41667
rect 86854 41611 86922 41667
rect 86978 41611 87046 41667
rect 87102 41611 87126 41667
rect 86526 41543 87126 41611
rect 86526 41487 86550 41543
rect 86606 41487 86674 41543
rect 86730 41487 86798 41543
rect 86854 41487 86922 41543
rect 86978 41487 87046 41543
rect 87102 41487 87126 41543
rect 86526 41419 87126 41487
rect 86526 41363 86550 41419
rect 86606 41363 86674 41419
rect 86730 41363 86798 41419
rect 86854 41363 86922 41419
rect 86978 41363 87046 41419
rect 87102 41363 87126 41419
rect 86526 41295 87126 41363
rect 86526 41239 86550 41295
rect 86606 41239 86674 41295
rect 86730 41239 86798 41295
rect 86854 41239 86922 41295
rect 86978 41239 87046 41295
rect 87102 41239 87126 41295
rect 86526 41171 87126 41239
rect 86526 41115 86550 41171
rect 86606 41115 86674 41171
rect 86730 41115 86798 41171
rect 86854 41115 86922 41171
rect 86978 41115 87046 41171
rect 87102 41115 87126 41171
rect 86526 41047 87126 41115
rect 86526 40991 86550 41047
rect 86606 40991 86674 41047
rect 86730 40991 86798 41047
rect 86854 40991 86922 41047
rect 86978 40991 87046 41047
rect 87102 40991 87126 41047
rect 86526 40923 87126 40991
rect 86526 40867 86550 40923
rect 86606 40867 86674 40923
rect 86730 40867 86798 40923
rect 86854 40867 86922 40923
rect 86978 40867 87046 40923
rect 87102 40867 87126 40923
rect 86526 40799 87126 40867
rect 86526 40743 86550 40799
rect 86606 40743 86674 40799
rect 86730 40743 86798 40799
rect 86854 40743 86922 40799
rect 86978 40743 87046 40799
rect 87102 40743 87126 40799
rect 86526 40675 87126 40743
rect 86526 40619 86550 40675
rect 86606 40619 86674 40675
rect 86730 40619 86798 40675
rect 86854 40619 86922 40675
rect 86978 40619 87046 40675
rect 87102 40619 87126 40675
rect 86526 40551 87126 40619
rect 86526 40495 86550 40551
rect 86606 40495 86674 40551
rect 86730 40495 86798 40551
rect 86854 40495 86922 40551
rect 86978 40495 87046 40551
rect 87102 40495 87126 40551
rect 86526 40427 87126 40495
rect 86526 40371 86550 40427
rect 86606 40371 86674 40427
rect 86730 40371 86798 40427
rect 86854 40371 86922 40427
rect 86978 40371 87046 40427
rect 87102 40371 87126 40427
rect 86526 40303 87126 40371
rect 86526 40247 86550 40303
rect 86606 40247 86674 40303
rect 86730 40247 86798 40303
rect 86854 40247 86922 40303
rect 86978 40247 87046 40303
rect 87102 40247 87126 40303
rect 86526 40179 87126 40247
rect 86526 40123 86550 40179
rect 86606 40123 86674 40179
rect 86730 40123 86798 40179
rect 86854 40123 86922 40179
rect 86978 40123 87046 40179
rect 87102 40123 87126 40179
rect 86526 40055 87126 40123
rect 86526 39999 86550 40055
rect 86606 39999 86674 40055
rect 86730 39999 86798 40055
rect 86854 39999 86922 40055
rect 86978 39999 87046 40055
rect 87102 39999 87126 40055
rect 86526 33187 87126 39999
rect 86526 33131 86550 33187
rect 86606 33131 86674 33187
rect 86730 33131 86798 33187
rect 86854 33131 86922 33187
rect 86978 33131 87046 33187
rect 87102 33131 87126 33187
rect 86526 33063 87126 33131
rect 86526 33007 86550 33063
rect 86606 33007 86674 33063
rect 86730 33007 86798 33063
rect 86854 33007 86922 33063
rect 86978 33007 87046 33063
rect 87102 33007 87126 33063
rect 86526 32939 87126 33007
rect 86526 32883 86550 32939
rect 86606 32883 86674 32939
rect 86730 32883 86798 32939
rect 86854 32883 86922 32939
rect 86978 32883 87046 32939
rect 87102 32883 87126 32939
rect 86526 32815 87126 32883
rect 86526 32759 86550 32815
rect 86606 32759 86674 32815
rect 86730 32759 86798 32815
rect 86854 32759 86922 32815
rect 86978 32759 87046 32815
rect 87102 32759 87126 32815
rect 86526 32691 87126 32759
rect 86526 32635 86550 32691
rect 86606 32635 86674 32691
rect 86730 32635 86798 32691
rect 86854 32635 86922 32691
rect 86978 32635 87046 32691
rect 87102 32635 87126 32691
rect 86526 32567 87126 32635
rect 86526 32511 86550 32567
rect 86606 32511 86674 32567
rect 86730 32511 86798 32567
rect 86854 32511 86922 32567
rect 86978 32511 87046 32567
rect 87102 32511 87126 32567
rect 86526 32443 87126 32511
rect 86526 32387 86550 32443
rect 86606 32387 86674 32443
rect 86730 32387 86798 32443
rect 86854 32387 86922 32443
rect 86978 32387 87046 32443
rect 87102 32387 87126 32443
rect 86526 32319 87126 32387
rect 86526 32263 86550 32319
rect 86606 32263 86674 32319
rect 86730 32263 86798 32319
rect 86854 32263 86922 32319
rect 86978 32263 87046 32319
rect 87102 32263 87126 32319
rect 86526 32195 87126 32263
rect 86526 32139 86550 32195
rect 86606 32139 86674 32195
rect 86730 32139 86798 32195
rect 86854 32139 86922 32195
rect 86978 32139 87046 32195
rect 87102 32139 87126 32195
rect 86526 32071 87126 32139
rect 86526 32015 86550 32071
rect 86606 32015 86674 32071
rect 86730 32015 86798 32071
rect 86854 32015 86922 32071
rect 86978 32015 87046 32071
rect 87102 32015 87126 32071
rect 86526 31947 87126 32015
rect 86526 31891 86550 31947
rect 86606 31891 86674 31947
rect 86730 31891 86798 31947
rect 86854 31891 86922 31947
rect 86978 31891 87046 31947
rect 87102 31891 87126 31947
rect 86526 31823 87126 31891
rect 86526 31767 86550 31823
rect 86606 31767 86674 31823
rect 86730 31767 86798 31823
rect 86854 31767 86922 31823
rect 86978 31767 87046 31823
rect 87102 31767 87126 31823
rect 86526 31699 87126 31767
rect 86526 31643 86550 31699
rect 86606 31643 86674 31699
rect 86730 31643 86798 31699
rect 86854 31643 86922 31699
rect 86978 31643 87046 31699
rect 87102 31643 87126 31699
rect 86526 31575 87126 31643
rect 86526 31519 86550 31575
rect 86606 31519 86674 31575
rect 86730 31519 86798 31575
rect 86854 31519 86922 31575
rect 86978 31519 87046 31575
rect 87102 31519 87126 31575
rect 86526 31451 87126 31519
rect 86526 31395 86550 31451
rect 86606 31395 86674 31451
rect 86730 31395 86798 31451
rect 86854 31395 86922 31451
rect 86978 31395 87046 31451
rect 87102 31395 87126 31451
rect 86526 31327 87126 31395
rect 86526 31271 86550 31327
rect 86606 31271 86674 31327
rect 86730 31271 86798 31327
rect 86854 31271 86922 31327
rect 86978 31271 87046 31327
rect 87102 31271 87126 31327
rect 86526 31203 87126 31271
rect 86526 31147 86550 31203
rect 86606 31147 86674 31203
rect 86730 31147 86798 31203
rect 86854 31147 86922 31203
rect 86978 31147 87046 31203
rect 87102 31147 87126 31203
rect 86526 31079 87126 31147
rect 86526 31023 86550 31079
rect 86606 31023 86674 31079
rect 86730 31023 86798 31079
rect 86854 31023 86922 31079
rect 86978 31023 87046 31079
rect 87102 31023 87126 31079
rect 86526 30955 87126 31023
rect 86526 30899 86550 30955
rect 86606 30899 86674 30955
rect 86730 30899 86798 30955
rect 86854 30899 86922 30955
rect 86978 30899 87046 30955
rect 87102 30899 87126 30955
rect 86526 30831 87126 30899
rect 86526 30775 86550 30831
rect 86606 30775 86674 30831
rect 86730 30775 86798 30831
rect 86854 30775 86922 30831
rect 86978 30775 87046 30831
rect 87102 30775 87126 30831
rect 86526 30707 87126 30775
rect 86526 30651 86550 30707
rect 86606 30651 86674 30707
rect 86730 30651 86798 30707
rect 86854 30651 86922 30707
rect 86978 30651 87046 30707
rect 87102 30651 87126 30707
rect 86526 30583 87126 30651
rect 86526 30527 86550 30583
rect 86606 30527 86674 30583
rect 86730 30527 86798 30583
rect 86854 30527 86922 30583
rect 86978 30527 87046 30583
rect 87102 30527 87126 30583
rect 86526 30459 87126 30527
rect 86526 30403 86550 30459
rect 86606 30403 86674 30459
rect 86730 30403 86798 30459
rect 86854 30403 86922 30459
rect 86978 30403 87046 30459
rect 87102 30403 87126 30459
rect 86526 30335 87126 30403
rect 86526 30279 86550 30335
rect 86606 30279 86674 30335
rect 86730 30279 86798 30335
rect 86854 30279 86922 30335
rect 86978 30279 87046 30335
rect 87102 30279 87126 30335
rect 86526 30211 87126 30279
rect 86526 30155 86550 30211
rect 86606 30155 86674 30211
rect 86730 30155 86798 30211
rect 86854 30155 86922 30211
rect 86978 30155 87046 30211
rect 87102 30155 87126 30211
rect 86526 30087 87126 30155
rect 86526 30031 86550 30087
rect 86606 30031 86674 30087
rect 86730 30031 86798 30087
rect 86854 30031 86922 30087
rect 86978 30031 87046 30087
rect 87102 30031 87126 30087
rect 86526 29963 87126 30031
rect 86526 29907 86550 29963
rect 86606 29907 86674 29963
rect 86730 29907 86798 29963
rect 86854 29907 86922 29963
rect 86978 29907 87046 29963
rect 87102 29907 87126 29963
rect 86526 26256 87126 29907
rect 86526 26200 86550 26256
rect 86606 26200 86674 26256
rect 86730 26200 86798 26256
rect 86854 26200 86922 26256
rect 86978 26200 87046 26256
rect 87102 26200 87126 26256
rect 86526 26132 87126 26200
rect 86526 26076 86550 26132
rect 86606 26076 86674 26132
rect 86730 26076 86798 26132
rect 86854 26076 86922 26132
rect 86978 26076 87046 26132
rect 87102 26076 87126 26132
rect 86526 26008 87126 26076
rect 86526 25952 86550 26008
rect 86606 25952 86674 26008
rect 86730 25952 86798 26008
rect 86854 25952 86922 26008
rect 86978 25952 87046 26008
rect 87102 25952 87126 26008
rect 86526 25884 87126 25952
rect 86526 25828 86550 25884
rect 86606 25828 86674 25884
rect 86730 25828 86798 25884
rect 86854 25828 86922 25884
rect 86978 25828 87046 25884
rect 87102 25828 87126 25884
rect 86526 25760 87126 25828
rect 86526 25704 86550 25760
rect 86606 25704 86674 25760
rect 86730 25704 86798 25760
rect 86854 25704 86922 25760
rect 86978 25704 87046 25760
rect 87102 25704 87126 25760
rect 86526 25636 87126 25704
rect 86526 25580 86550 25636
rect 86606 25580 86674 25636
rect 86730 25580 86798 25636
rect 86854 25580 86922 25636
rect 86978 25580 87046 25636
rect 87102 25580 87126 25636
rect 86526 25512 87126 25580
rect 86526 25456 86550 25512
rect 86606 25456 86674 25512
rect 86730 25456 86798 25512
rect 86854 25456 86922 25512
rect 86978 25456 87046 25512
rect 87102 25456 87126 25512
rect 86526 25388 87126 25456
rect 86526 25332 86550 25388
rect 86606 25332 86674 25388
rect 86730 25332 86798 25388
rect 86854 25332 86922 25388
rect 86978 25332 87046 25388
rect 87102 25332 87126 25388
rect 86526 12859 87126 25332
rect 86526 12803 86612 12859
rect 86668 12803 86736 12859
rect 86792 12803 86860 12859
rect 86916 12803 86984 12859
rect 87040 12803 87126 12859
rect 86526 12735 87126 12803
rect 86526 12679 86612 12735
rect 86668 12679 86736 12735
rect 86792 12679 86860 12735
rect 86916 12679 86984 12735
rect 87040 12679 87126 12735
rect 86526 12611 87126 12679
rect 86526 12555 86612 12611
rect 86668 12555 86736 12611
rect 86792 12555 86860 12611
rect 86916 12555 86984 12611
rect 87040 12555 87126 12611
rect 86526 12487 87126 12555
rect 86526 12431 86612 12487
rect 86668 12431 86736 12487
rect 86792 12431 86860 12487
rect 86916 12431 86984 12487
rect 87040 12431 87126 12487
rect 86526 10764 87126 12431
rect 86526 10708 86612 10764
rect 86668 10708 86736 10764
rect 86792 10708 86860 10764
rect 86916 10708 86984 10764
rect 87040 10708 87126 10764
rect 86526 10640 87126 10708
rect 86526 10584 86612 10640
rect 86668 10584 86736 10640
rect 86792 10584 86860 10640
rect 86916 10584 86984 10640
rect 87040 10584 87126 10640
rect 86526 10516 87126 10584
rect 86526 10460 86612 10516
rect 86668 10460 86736 10516
rect 86792 10460 86860 10516
rect 86916 10460 86984 10516
rect 87040 10460 87126 10516
rect 86526 10392 87126 10460
rect 86526 10336 86612 10392
rect 86668 10336 86736 10392
rect 86792 10336 86860 10392
rect 86916 10336 86984 10392
rect 87040 10336 87126 10392
rect 86526 8964 87126 10336
rect 86526 8908 86612 8964
rect 86668 8908 86736 8964
rect 86792 8908 86860 8964
rect 86916 8908 86984 8964
rect 87040 8908 87126 8964
rect 86526 8840 87126 8908
rect 86526 8784 86612 8840
rect 86668 8784 86736 8840
rect 86792 8784 86860 8840
rect 86916 8784 86984 8840
rect 87040 8784 87126 8840
rect 86526 8716 87126 8784
rect 86526 8660 86612 8716
rect 86668 8660 86736 8716
rect 86792 8660 86860 8716
rect 86916 8660 86984 8716
rect 87040 8660 87126 8716
rect 86526 8592 87126 8660
rect 86526 8536 86612 8592
rect 86668 8536 86736 8592
rect 86792 8536 86860 8592
rect 86916 8536 86984 8592
rect 87040 8536 87126 8592
rect 86526 7164 87126 8536
rect 86526 7108 86612 7164
rect 86668 7108 86736 7164
rect 86792 7108 86860 7164
rect 86916 7108 86984 7164
rect 87040 7108 87126 7164
rect 86526 7040 87126 7108
rect 86526 6984 86612 7040
rect 86668 6984 86736 7040
rect 86792 6984 86860 7040
rect 86916 6984 86984 7040
rect 87040 6984 87126 7040
rect 86526 6916 87126 6984
rect 86526 6860 86612 6916
rect 86668 6860 86736 6916
rect 86792 6860 86860 6916
rect 86916 6860 86984 6916
rect 87040 6860 87126 6916
rect 86526 6792 87126 6860
rect 86526 6736 86612 6792
rect 86668 6736 86736 6792
rect 86792 6736 86860 6792
rect 86916 6736 86984 6792
rect 87040 6736 87126 6792
rect 86526 5364 87126 6736
rect 86526 5308 86612 5364
rect 86668 5308 86736 5364
rect 86792 5308 86860 5364
rect 86916 5308 86984 5364
rect 87040 5308 87126 5364
rect 86526 5240 87126 5308
rect 86526 5184 86612 5240
rect 86668 5184 86736 5240
rect 86792 5184 86860 5240
rect 86916 5184 86984 5240
rect 87040 5184 87126 5240
rect 86526 5116 87126 5184
rect 86526 5060 86612 5116
rect 86668 5060 86736 5116
rect 86792 5060 86860 5116
rect 86916 5060 86984 5116
rect 87040 5060 87126 5116
rect 86526 4992 87126 5060
rect 86526 4936 86612 4992
rect 86668 4936 86736 4992
rect 86792 4936 86860 4992
rect 86916 4936 86984 4992
rect 87040 4936 87126 4992
rect 86526 3632 87126 4936
rect 86526 3576 86612 3632
rect 86668 3576 86736 3632
rect 86792 3576 86860 3632
rect 86916 3576 86984 3632
rect 87040 3576 87126 3632
rect 86526 3508 87126 3576
rect 86526 3452 86612 3508
rect 86668 3452 86736 3508
rect 86792 3452 86860 3508
rect 86916 3452 86984 3508
rect 87040 3452 87126 3508
rect 86526 3384 87126 3452
rect 86526 3328 86612 3384
rect 86668 3328 86736 3384
rect 86792 3328 86860 3384
rect 86916 3328 86984 3384
rect 87040 3328 87126 3384
rect 86526 3260 87126 3328
rect 86526 3204 86612 3260
rect 86668 3204 86736 3260
rect 86792 3204 86860 3260
rect 86916 3204 86984 3260
rect 87040 3204 87126 3260
rect 86526 3136 87126 3204
use gf180mcu_fd_ip_sram__sram64x8m8wm1  RAM
timestamp 0
transform -1 0 87372 0 -1 47576
box 0 0 86372 46576
<< labels >>
flabel metal2 s 52944 47976 53056 48776 0 FreeSans 448 90 0 0 A[0]
port 0 nsew signal input
flabel metal2 s 54644 47976 54756 48776 0 FreeSans 448 90 0 0 A[1]
port 1 nsew signal input
flabel metal2 s 56344 47976 56456 48776 0 FreeSans 448 90 0 0 A[2]
port 2 nsew signal input
flabel metal2 s 30944 47976 31056 48776 0 FreeSans 448 90 0 0 A[3]
port 3 nsew signal input
flabel metal2 s 31944 47976 32056 48776 0 FreeSans 448 90 0 0 A[4]
port 4 nsew signal input
flabel metal2 s 32744 47976 32856 48776 0 FreeSans 448 90 0 0 A[5]
port 5 nsew signal input
flabel metal2 s 36844 47976 36956 48776 0 FreeSans 448 90 0 0 CEN
port 6 nsew signal input
flabel metal2 s 59244 47976 59356 48776 0 FreeSans 448 90 0 0 CLK
port 7 nsew signal input
flabel metal2 s 85344 47976 85456 48776 0 FreeSans 448 90 0 0 D[0]
port 8 nsew signal input
flabel metal2 s 74944 47976 75056 48776 0 FreeSans 448 90 0 0 D[1]
port 9 nsew signal input
flabel metal2 s 73744 47976 73856 48776 0 FreeSans 448 90 0 0 D[2]
port 10 nsew signal input
flabel metal2 s 63344 47976 63456 48776 0 FreeSans 448 90 0 0 D[3]
port 11 nsew signal input
flabel metal2 s 25744 47976 25856 48776 0 FreeSans 448 90 0 0 D[4]
port 12 nsew signal input
flabel metal2 s 15444 47976 15556 48776 0 FreeSans 448 90 0 0 D[5]
port 13 nsew signal input
flabel metal2 s 14144 47976 14256 48776 0 FreeSans 448 90 0 0 D[6]
port 14 nsew signal input
flabel metal2 s 3744 47976 3856 48776 0 FreeSans 448 90 0 0 D[7]
port 15 nsew signal input
flabel metal2 s 46568 47976 46680 48776 0 FreeSans 448 90 0 0 GWEN
port 16 nsew signal input
flabel metal2 s 83844 47976 83956 48776 0 FreeSans 448 90 0 0 Q[0]
port 17 nsew signal tristate
flabel metal2 s 75644 47976 75756 48776 0 FreeSans 448 90 0 0 Q[1]
port 18 nsew signal tristate
flabel metal2 s 73044 47976 73156 48776 0 FreeSans 448 90 0 0 Q[2]
port 19 nsew signal tristate
flabel metal2 s 64944 47976 65056 48776 0 FreeSans 448 90 0 0 Q[3]
port 20 nsew signal tristate
flabel metal2 s 24244 47976 24356 48776 0 FreeSans 448 90 0 0 Q[4]
port 21 nsew signal tristate
flabel metal2 s 16044 47976 16156 48776 0 FreeSans 448 90 0 0 Q[5]
port 22 nsew signal tristate
flabel metal2 s 13444 47976 13556 48776 0 FreeSans 448 90 0 0 Q[6]
port 23 nsew signal tristate
flabel metal2 s 5344 47976 5456 48776 0 FreeSans 448 90 0 0 Q[7]
port 24 nsew signal tristate
flabel metal4 s 1044 3136 1644 45472 0 FreeSans 2560 90 0 0 VDD
port 25 nsew power bidirectional
flabel metal4 s 85726 3136 86326 45472 0 FreeSans 2560 90 0 0 VDD
port 25 nsew power bidirectional
flabel metal4 s 1844 3136 2444 45472 0 FreeSans 2560 90 0 0 VSS
port 26 nsew ground bidirectional
flabel metal4 s 86526 3136 87126 45472 0 FreeSans 2560 90 0 0 VSS
port 26 nsew ground bidirectional
flabel metal2 s 84644 47976 84756 48776 0 FreeSans 448 90 0 0 WEN[0]
port 27 nsew signal input
flabel metal2 s 74544 47976 74656 48776 0 FreeSans 448 90 0 0 WEN[1]
port 28 nsew signal input
flabel metal2 s 74144 47976 74256 48776 0 FreeSans 448 90 0 0 WEN[2]
port 29 nsew signal input
flabel metal2 s 63744 47976 63856 48776 0 FreeSans 448 90 0 0 WEN[3]
port 30 nsew signal input
flabel metal2 s 25044 47976 25156 48776 0 FreeSans 448 90 0 0 WEN[4]
port 31 nsew signal input
flabel metal2 s 14994 47976 15106 48776 0 FreeSans 448 90 0 0 WEN[5]
port 32 nsew signal input
flabel metal2 s 14544 47976 14656 48776 0 FreeSans 448 90 0 0 WEN[6]
port 33 nsew signal input
flabel metal2 s 4444 47976 4556 48776 0 FreeSans 448 90 0 0 WEN[7]
port 34 nsew signal input
rlabel via3 86212 45408 86212 45408 0 VDD
rlabel via3 87074 44997 87074 44997 0 VSS
rlabel metal2 53032 47824 53032 47824 0 A[0]
rlabel metal2 54712 47824 54712 47824 0 A[1]
rlabel metal2 56392 47824 56392 47824 0 A[2]
rlabel metal2 30968 47824 30968 47824 0 A[3]
rlabel metal2 32032 47670 32032 47670 0 A[4]
rlabel metal2 32760 47824 32760 47824 0 A[5]
rlabel metal2 36904 47824 36904 47824 0 CEN
rlabel metal2 59304 47824 59304 47824 0 CLK
rlabel metal2 85400 47824 85400 47824 0 D[0]
rlabel metal2 74984 47824 74984 47824 0 D[1]
rlabel metal2 73752 47824 73752 47824 0 D[2]
rlabel metal2 63448 47824 63448 47824 0 D[3]
rlabel metal2 25816 47824 25816 47824 0 D[4]
rlabel metal2 15512 47824 15512 47824 0 D[5]
rlabel metal2 14168 47824 14168 47824 0 D[6]
rlabel metal2 3808 47670 3808 47670 0 D[7]
rlabel metal2 46648 47824 46648 47824 0 GWEN
rlabel metal2 83944 47824 83944 47824 0 Q[0]
rlabel metal2 75656 47824 75656 47824 0 Q[1]
rlabel metal2 73080 47824 73080 47824 0 Q[2]
rlabel metal2 65016 47824 65016 47824 0 Q[3]
rlabel metal2 24248 47824 24248 47824 0 Q[4]
rlabel metal2 16072 47824 16072 47824 0 Q[5]
rlabel metal2 13496 47824 13496 47824 0 Q[6]
rlabel metal2 5432 47824 5432 47824 0 Q[7]
rlabel metal2 84728 47824 84728 47824 0 WEN[0]
rlabel metal2 74648 47824 74648 47824 0 WEN[1]
rlabel metal2 74200 47824 74200 47824 0 WEN[2]
rlabel metal2 63784 47824 63784 47824 0 WEN[3]
rlabel metal2 25144 47824 25144 47824 0 WEN[4]
rlabel metal2 15064 47824 15064 47824 0 WEN[5]
rlabel metal2 14616 47824 14616 47824 0 WEN[6]
rlabel metal2 4536 47824 4536 47824 0 WEN[7]
<< properties >>
string FIXED_BBOX 0 0 88972 48776
<< end >>
