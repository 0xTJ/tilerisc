magic
tech gf180mcuD
magscale 1 5
timestamp 1700157470
<< obsm1 >>
rect 500 500 43686 34588
<< metal2 >>
rect 1872 34788 1928 35188
rect 2222 34788 2278 35188
rect 2672 34788 2728 35188
rect 6722 34788 6778 35188
rect 7072 34788 7128 35188
rect 7272 34788 7328 35188
rect 7497 34788 7553 35188
rect 7722 34788 7778 35188
rect 8022 34788 8078 35188
rect 12122 34788 12178 35188
rect 12522 34788 12578 35188
rect 12872 34788 12928 35188
rect 15472 34788 15528 35188
rect 15972 34788 16028 35188
rect 16372 34788 16428 35188
rect 16672 34788 16728 35188
rect 18422 34788 18478 35188
rect 23284 34788 23340 35188
rect 26472 34788 26528 35188
rect 27322 34788 27378 35188
rect 28172 34788 28228 35188
rect 28722 34788 28778 35188
rect 29622 34788 29678 35188
rect 31672 34788 31728 35188
rect 31872 34788 31928 35188
rect 32472 34788 32528 35188
rect 36522 34788 36578 35188
rect 36872 34788 36928 35188
rect 37072 34788 37128 35188
rect 37272 34788 37328 35188
rect 37472 34788 37528 35188
rect 37822 34788 37878 35188
rect 41922 34788 41978 35188
rect 42322 34788 42378 35188
rect 42672 34788 42728 35188
<< obsm2 >>
rect 500 34758 1842 34804
rect 1958 34758 2192 34804
rect 2308 34758 2642 34804
rect 2758 34758 6692 34804
rect 6808 34758 7042 34804
rect 7158 34758 7242 34804
rect 7358 34758 7467 34804
rect 7583 34758 7692 34804
rect 7808 34758 7992 34804
rect 8108 34758 12092 34804
rect 12208 34758 12492 34804
rect 12608 34758 12842 34804
rect 12958 34758 15442 34804
rect 15558 34758 15942 34804
rect 16058 34758 16342 34804
rect 16458 34758 16642 34804
rect 16758 34758 18392 34804
rect 18508 34758 23254 34804
rect 23370 34758 26442 34804
rect 26558 34758 27292 34804
rect 27408 34758 28142 34804
rect 28258 34758 28692 34804
rect 28808 34758 29592 34804
rect 29708 34758 31642 34804
rect 31758 34758 31842 34804
rect 31958 34758 32442 34804
rect 32558 34758 36492 34804
rect 36608 34758 36842 34804
rect 36958 34758 37042 34804
rect 37158 34758 37242 34804
rect 37358 34758 37442 34804
rect 37558 34758 37792 34804
rect 37908 34758 41892 34804
rect 42008 34758 42292 34804
rect 42408 34758 42642 34804
rect 42758 34758 43686 34804
rect 500 500 43686 34758
<< obsm3 >>
rect 500 500 43686 34588
<< metal4 >>
rect 522 1568 822 33320
rect 922 1568 1222 33320
rect 42863 1568 43163 33320
rect 43263 1568 43563 33320
<< labels >>
rlabel metal2 s 26472 34788 26528 35188 6 A[0]
port 1 nsew signal input
rlabel metal2 s 27322 34788 27378 35188 6 A[1]
port 2 nsew signal input
rlabel metal2 s 28172 34788 28228 35188 6 A[2]
port 3 nsew signal input
rlabel metal2 s 15472 34788 15528 35188 6 A[3]
port 4 nsew signal input
rlabel metal2 s 15972 34788 16028 35188 6 A[4]
port 5 nsew signal input
rlabel metal2 s 16372 34788 16428 35188 6 A[5]
port 6 nsew signal input
rlabel metal2 s 16672 34788 16728 35188 6 A[6]
port 7 nsew signal input
rlabel metal2 s 28722 34788 28778 35188 6 A[7]
port 8 nsew signal input
rlabel metal2 s 18422 34788 18478 35188 6 CEN
port 9 nsew signal input
rlabel metal2 s 29622 34788 29678 35188 6 CLK
port 10 nsew signal input
rlabel metal2 s 42672 34788 42728 35188 6 D[0]
port 11 nsew signal input
rlabel metal2 s 37472 34788 37528 35188 6 D[1]
port 12 nsew signal input
rlabel metal2 s 36872 34788 36928 35188 6 D[2]
port 13 nsew signal input
rlabel metal2 s 31672 34788 31728 35188 6 D[3]
port 14 nsew signal input
rlabel metal2 s 12872 34788 12928 35188 6 D[4]
port 15 nsew signal input
rlabel metal2 s 7722 34788 7778 35188 6 D[5]
port 16 nsew signal input
rlabel metal2 s 7072 34788 7128 35188 6 D[6]
port 17 nsew signal input
rlabel metal2 s 1872 34788 1928 35188 6 D[7]
port 18 nsew signal input
rlabel metal2 s 23284 34788 23340 35188 6 GWEN
port 19 nsew signal input
rlabel metal2 s 41922 34788 41978 35188 6 Q[0]
port 20 nsew signal output
rlabel metal2 s 37822 34788 37878 35188 6 Q[1]
port 21 nsew signal output
rlabel metal2 s 36522 34788 36578 35188 6 Q[2]
port 22 nsew signal output
rlabel metal2 s 32472 34788 32528 35188 6 Q[3]
port 23 nsew signal output
rlabel metal2 s 12122 34788 12178 35188 6 Q[4]
port 24 nsew signal output
rlabel metal2 s 8022 34788 8078 35188 6 Q[5]
port 25 nsew signal output
rlabel metal2 s 6722 34788 6778 35188 6 Q[6]
port 26 nsew signal output
rlabel metal2 s 2672 34788 2728 35188 6 Q[7]
port 27 nsew signal output
rlabel metal4 s 522 1568 822 33320 6 VDD
port 28 nsew power bidirectional
rlabel metal4 s 42863 1568 43163 33320 6 VDD
port 28 nsew power bidirectional
rlabel metal4 s 922 1568 1222 33320 6 VSS
port 29 nsew ground bidirectional
rlabel metal4 s 43263 1568 43563 33320 6 VSS
port 29 nsew ground bidirectional
rlabel metal2 s 42322 34788 42378 35188 6 WEN[0]
port 30 nsew signal input
rlabel metal2 s 37272 34788 37328 35188 6 WEN[1]
port 31 nsew signal input
rlabel metal2 s 37072 34788 37128 35188 6 WEN[2]
port 32 nsew signal input
rlabel metal2 s 31872 34788 31928 35188 6 WEN[3]
port 33 nsew signal input
rlabel metal2 s 12522 34788 12578 35188 6 WEN[4]
port 34 nsew signal input
rlabel metal2 s 7497 34788 7553 35188 6 WEN[5]
port 35 nsew signal input
rlabel metal2 s 7272 34788 7328 35188 6 WEN[6]
port 36 nsew signal input
rlabel metal2 s 2222 34788 2278 35188 6 WEN[7]
port 37 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 44486 35188
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2585266
string GDS_FILE /home/thomas/Documents/Projects/tilerisc/openlane/gf180_ram_256x8_wrapper/runs/23_11_16_12_57/results/signoff/gf180_ram_256x8_wrapper.magic.gds
string GDS_START 2452566
<< end >>

