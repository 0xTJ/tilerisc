magic
tech gf180mcuD
magscale 1 10
timestamp 1700487504
<< metal1 >>
rect 1344 36874 58576 36908
rect 1344 36822 8367 36874
rect 8419 36822 8471 36874
rect 8523 36822 8575 36874
rect 8627 36822 22674 36874
rect 22726 36822 22778 36874
rect 22830 36822 22882 36874
rect 22934 36822 36981 36874
rect 37033 36822 37085 36874
rect 37137 36822 37189 36874
rect 37241 36822 51288 36874
rect 51340 36822 51392 36874
rect 51444 36822 51496 36874
rect 51548 36822 58576 36874
rect 1344 36788 58576 36822
rect 41918 36594 41970 36606
rect 4610 36542 4622 36594
rect 4674 36542 4686 36594
rect 8754 36542 8766 36594
rect 8818 36542 8830 36594
rect 12562 36542 12574 36594
rect 12626 36542 12638 36594
rect 14802 36542 14814 36594
rect 14866 36542 14878 36594
rect 17378 36542 17390 36594
rect 17442 36542 17454 36594
rect 19282 36542 19294 36594
rect 19346 36542 19358 36594
rect 21522 36542 21534 36594
rect 21586 36542 21598 36594
rect 23202 36542 23214 36594
rect 23266 36542 23278 36594
rect 25666 36542 25678 36594
rect 25730 36542 25742 36594
rect 27346 36542 27358 36594
rect 27410 36542 27422 36594
rect 31266 36542 31278 36594
rect 31330 36542 31342 36594
rect 35410 36542 35422 36594
rect 35474 36542 35486 36594
rect 36530 36542 36542 36594
rect 36594 36542 36606 36594
rect 41918 36530 41970 36542
rect 43038 36594 43090 36606
rect 55022 36594 55074 36606
rect 43922 36542 43934 36594
rect 43986 36542 43998 36594
rect 43038 36530 43090 36542
rect 55022 36530 55074 36542
rect 56926 36594 56978 36606
rect 56926 36530 56978 36542
rect 14366 36482 14418 36494
rect 42254 36482 42306 36494
rect 48862 36482 48914 36494
rect 1810 36430 1822 36482
rect 1874 36430 1886 36482
rect 5842 36430 5854 36482
rect 5906 36430 5918 36482
rect 9762 36430 9774 36482
rect 9826 36430 9838 36482
rect 24994 36430 25006 36482
rect 25058 36430 25070 36482
rect 28466 36430 28478 36482
rect 28530 36430 28542 36482
rect 32610 36430 32622 36482
rect 32674 36430 32686 36482
rect 37202 36430 37214 36482
rect 37266 36430 37278 36482
rect 37986 36430 37998 36482
rect 38050 36430 38062 36482
rect 38546 36430 38558 36482
rect 38610 36430 38622 36482
rect 40786 36430 40798 36482
rect 40850 36430 40862 36482
rect 41346 36430 41358 36482
rect 41410 36430 41422 36482
rect 46722 36430 46734 36482
rect 46786 36430 46798 36482
rect 49410 36430 49422 36482
rect 49474 36430 49486 36482
rect 52770 36430 52782 36482
rect 52834 36430 52846 36482
rect 53106 36430 53118 36482
rect 53170 36430 53182 36482
rect 53778 36430 53790 36482
rect 53842 36430 53854 36482
rect 55458 36430 55470 36482
rect 55522 36430 55534 36482
rect 14366 36418 14418 36430
rect 42254 36418 42306 36430
rect 48862 36418 48914 36430
rect 15822 36370 15874 36382
rect 47406 36370 47458 36382
rect 2482 36318 2494 36370
rect 2546 36318 2558 36370
rect 6626 36318 6638 36370
rect 6690 36318 6702 36370
rect 10434 36318 10446 36370
rect 10498 36318 10510 36370
rect 29138 36318 29150 36370
rect 29202 36318 29214 36370
rect 33282 36318 33294 36370
rect 33346 36318 33358 36370
rect 39218 36318 39230 36370
rect 39282 36318 39294 36370
rect 39890 36318 39902 36370
rect 39954 36318 39966 36370
rect 46050 36318 46062 36370
rect 46114 36318 46126 36370
rect 15822 36306 15874 36318
rect 47406 36306 47458 36318
rect 48302 36370 48354 36382
rect 48302 36306 48354 36318
rect 49198 36370 49250 36382
rect 49198 36306 49250 36318
rect 50542 36370 50594 36382
rect 56478 36370 56530 36382
rect 51650 36318 51662 36370
rect 51714 36318 51726 36370
rect 50542 36306 50594 36318
rect 56478 36306 56530 36318
rect 13246 36258 13298 36270
rect 13246 36194 13298 36206
rect 13694 36258 13746 36270
rect 13694 36194 13746 36206
rect 16158 36258 16210 36270
rect 16158 36194 16210 36206
rect 16942 36258 16994 36270
rect 16942 36194 16994 36206
rect 18510 36258 18562 36270
rect 18510 36194 18562 36206
rect 18846 36258 18898 36270
rect 18846 36194 18898 36206
rect 20302 36258 20354 36270
rect 20302 36194 20354 36206
rect 21086 36258 21138 36270
rect 21086 36194 21138 36206
rect 22542 36258 22594 36270
rect 22542 36194 22594 36206
rect 22766 36258 22818 36270
rect 22766 36194 22818 36206
rect 24110 36258 24162 36270
rect 24110 36194 24162 36206
rect 24670 36258 24722 36270
rect 24670 36194 24722 36206
rect 26686 36258 26738 36270
rect 26686 36194 26738 36206
rect 27806 36258 27858 36270
rect 27806 36194 27858 36206
rect 42590 36258 42642 36270
rect 42590 36194 42642 36206
rect 47742 36258 47794 36270
rect 47742 36194 47794 36206
rect 50206 36258 50258 36270
rect 50206 36194 50258 36206
rect 53566 36258 53618 36270
rect 53566 36194 53618 36206
rect 54462 36258 54514 36270
rect 54462 36194 54514 36206
rect 56030 36258 56082 36270
rect 56030 36194 56082 36206
rect 1344 36090 58731 36124
rect 1344 36038 15520 36090
rect 15572 36038 15624 36090
rect 15676 36038 15728 36090
rect 15780 36038 29827 36090
rect 29879 36038 29931 36090
rect 29983 36038 30035 36090
rect 30087 36038 44134 36090
rect 44186 36038 44238 36090
rect 44290 36038 44342 36090
rect 44394 36038 58441 36090
rect 58493 36038 58545 36090
rect 58597 36038 58649 36090
rect 58701 36038 58731 36090
rect 1344 36004 58731 36038
rect 9886 35922 9938 35934
rect 9886 35858 9938 35870
rect 10670 35922 10722 35934
rect 10670 35858 10722 35870
rect 21646 35922 21698 35934
rect 21646 35858 21698 35870
rect 35534 35922 35586 35934
rect 35534 35858 35586 35870
rect 51438 35922 51490 35934
rect 51438 35858 51490 35870
rect 54686 35922 54738 35934
rect 54686 35858 54738 35870
rect 54798 35922 54850 35934
rect 54798 35858 54850 35870
rect 56030 35922 56082 35934
rect 56030 35858 56082 35870
rect 16270 35810 16322 35822
rect 2930 35758 2942 35810
rect 2994 35758 3006 35810
rect 4946 35758 4958 35810
rect 5010 35758 5022 35810
rect 16270 35746 16322 35758
rect 22766 35810 22818 35822
rect 40910 35810 40962 35822
rect 47630 35810 47682 35822
rect 37762 35758 37774 35810
rect 37826 35758 37838 35810
rect 39778 35758 39790 35810
rect 39842 35758 39854 35810
rect 42690 35758 42702 35810
rect 42754 35758 42766 35810
rect 44706 35758 44718 35810
rect 44770 35758 44782 35810
rect 22766 35746 22818 35758
rect 40910 35746 40962 35758
rect 47630 35746 47682 35758
rect 48750 35810 48802 35822
rect 55582 35810 55634 35822
rect 49074 35758 49086 35810
rect 49138 35758 49150 35810
rect 50642 35758 50654 35810
rect 50706 35758 50718 35810
rect 51762 35758 51774 35810
rect 51826 35758 51838 35810
rect 48750 35746 48802 35758
rect 55582 35746 55634 35758
rect 56702 35810 56754 35822
rect 56702 35746 56754 35758
rect 1710 35698 1762 35710
rect 7646 35698 7698 35710
rect 22542 35698 22594 35710
rect 3826 35646 3838 35698
rect 3890 35646 3902 35698
rect 4162 35646 4174 35698
rect 4226 35646 4238 35698
rect 11666 35646 11678 35698
rect 11730 35646 11742 35698
rect 13122 35646 13134 35698
rect 13186 35646 13198 35698
rect 16482 35646 16494 35698
rect 16546 35646 16558 35698
rect 18274 35646 18286 35698
rect 18338 35646 18350 35698
rect 21410 35646 21422 35698
rect 21474 35646 21486 35698
rect 1710 35634 1762 35646
rect 7646 35634 7698 35646
rect 22542 35634 22594 35646
rect 22654 35698 22706 35710
rect 33070 35698 33122 35710
rect 41694 35698 41746 35710
rect 24210 35646 24222 35698
rect 24274 35646 24286 35698
rect 26002 35646 26014 35698
rect 26066 35646 26078 35698
rect 29586 35646 29598 35698
rect 29650 35646 29662 35698
rect 35858 35646 35870 35698
rect 35922 35646 35934 35698
rect 36418 35646 36430 35698
rect 36482 35646 36494 35698
rect 39890 35646 39902 35698
rect 39954 35646 39966 35698
rect 41122 35646 41134 35698
rect 41186 35646 41198 35698
rect 22654 35634 22706 35646
rect 33070 35634 33122 35646
rect 41694 35634 41746 35646
rect 43934 35698 43986 35710
rect 47966 35698 48018 35710
rect 54574 35698 54626 35710
rect 44818 35646 44830 35698
rect 44882 35646 44894 35698
rect 46386 35646 46398 35698
rect 46450 35646 46462 35698
rect 46834 35646 46846 35698
rect 46898 35646 46910 35698
rect 52770 35646 52782 35698
rect 52834 35646 52846 35698
rect 53554 35646 53566 35698
rect 53618 35646 53630 35698
rect 43934 35634 43986 35646
rect 47966 35634 48018 35646
rect 54574 35634 54626 35646
rect 55246 35698 55298 35710
rect 55246 35634 55298 35646
rect 56478 35698 56530 35710
rect 56478 35634 56530 35646
rect 56814 35698 56866 35710
rect 56814 35634 56866 35646
rect 8878 35586 8930 35598
rect 2146 35534 2158 35586
rect 2210 35534 2222 35586
rect 7074 35534 7086 35586
rect 7138 35534 7150 35586
rect 8082 35534 8094 35586
rect 8146 35534 8158 35586
rect 8878 35522 8930 35534
rect 11118 35586 11170 35598
rect 17838 35586 17890 35598
rect 25678 35586 25730 35598
rect 34526 35586 34578 35598
rect 42254 35586 42306 35598
rect 12114 35534 12126 35586
rect 12178 35534 12190 35586
rect 13794 35534 13806 35586
rect 13858 35534 13870 35586
rect 15922 35534 15934 35586
rect 15986 35534 15998 35586
rect 18946 35534 18958 35586
rect 19010 35534 19022 35586
rect 21074 35534 21086 35586
rect 21138 35534 21150 35586
rect 24434 35534 24446 35586
rect 24498 35534 24510 35586
rect 26786 35534 26798 35586
rect 26850 35534 26862 35586
rect 28914 35534 28926 35586
rect 28978 35534 28990 35586
rect 30370 35534 30382 35586
rect 30434 35534 30446 35586
rect 32498 35534 32510 35586
rect 32562 35534 32574 35586
rect 33730 35534 33742 35586
rect 33794 35534 33806 35586
rect 37426 35534 37438 35586
rect 37490 35534 37502 35586
rect 40114 35534 40126 35586
rect 40178 35534 40190 35586
rect 11118 35522 11170 35534
rect 17838 35522 17890 35534
rect 25678 35522 25730 35534
rect 34526 35522 34578 35534
rect 42254 35522 42306 35534
rect 43822 35586 43874 35598
rect 45602 35534 45614 35586
rect 45666 35534 45678 35586
rect 50866 35534 50878 35586
rect 50930 35534 50942 35586
rect 52098 35534 52110 35586
rect 52162 35534 52174 35586
rect 43822 35522 43874 35534
rect 21758 35474 21810 35486
rect 22082 35422 22094 35474
rect 22146 35422 22158 35474
rect 24546 35422 24558 35474
rect 24610 35422 24622 35474
rect 40226 35422 40238 35474
rect 40290 35422 40302 35474
rect 21758 35410 21810 35422
rect 1344 35306 58576 35340
rect 1344 35254 8367 35306
rect 8419 35254 8471 35306
rect 8523 35254 8575 35306
rect 8627 35254 22674 35306
rect 22726 35254 22778 35306
rect 22830 35254 22882 35306
rect 22934 35254 36981 35306
rect 37033 35254 37085 35306
rect 37137 35254 37189 35306
rect 37241 35254 51288 35306
rect 51340 35254 51392 35306
rect 51444 35254 51496 35306
rect 51548 35254 58576 35306
rect 1344 35220 58576 35254
rect 30494 35138 30546 35150
rect 30494 35074 30546 35086
rect 35086 35138 35138 35150
rect 35086 35074 35138 35086
rect 52894 35138 52946 35150
rect 53218 35086 53230 35138
rect 53282 35086 53294 35138
rect 52894 35074 52946 35086
rect 5070 35026 5122 35038
rect 14926 35026 14978 35038
rect 30158 35026 30210 35038
rect 5618 34974 5630 35026
rect 5682 34974 5694 35026
rect 11778 34974 11790 35026
rect 11842 34974 11854 35026
rect 16034 34974 16046 35026
rect 16098 34974 16110 35026
rect 18162 34974 18174 35026
rect 18226 34974 18238 35026
rect 25554 34974 25566 35026
rect 25618 34974 25630 35026
rect 5070 34962 5122 34974
rect 14926 34962 14978 34974
rect 30158 34962 30210 34974
rect 32174 35026 32226 35038
rect 51214 35026 51266 35038
rect 36978 34974 36990 35026
rect 37042 34974 37054 35026
rect 44034 34974 44046 35026
rect 44098 34974 44110 35026
rect 45826 34974 45838 35026
rect 45890 34974 45902 35026
rect 49074 34974 49086 35026
rect 49138 34974 49150 35026
rect 32174 34962 32226 34974
rect 51214 34962 51266 34974
rect 52670 35026 52722 35038
rect 58158 35026 58210 35038
rect 56690 34974 56702 35026
rect 56754 34974 56766 35026
rect 52670 34962 52722 34974
rect 58158 34962 58210 34974
rect 2270 34914 2322 34926
rect 1810 34862 1822 34914
rect 1874 34862 1886 34914
rect 2270 34850 2322 34862
rect 2606 34914 2658 34926
rect 2606 34850 2658 34862
rect 3166 34914 3218 34926
rect 3166 34850 3218 34862
rect 3502 34914 3554 34926
rect 3502 34850 3554 34862
rect 4062 34914 4114 34926
rect 20526 34914 20578 34926
rect 8530 34862 8542 34914
rect 8594 34862 8606 34914
rect 8978 34862 8990 34914
rect 9042 34862 9054 34914
rect 12338 34862 12350 34914
rect 12402 34862 12414 34914
rect 15250 34862 15262 34914
rect 15314 34862 15326 34914
rect 20290 34862 20302 34914
rect 20354 34862 20366 34914
rect 4062 34850 4114 34862
rect 20526 34850 20578 34862
rect 21646 34914 21698 34926
rect 22766 34914 22818 34926
rect 25902 34914 25954 34926
rect 22418 34862 22430 34914
rect 22482 34862 22494 34914
rect 23986 34862 23998 34914
rect 24050 34862 24062 34914
rect 21646 34850 21698 34862
rect 22766 34850 22818 34862
rect 25902 34850 25954 34862
rect 26462 34914 26514 34926
rect 31278 34914 31330 34926
rect 28130 34862 28142 34914
rect 28194 34862 28206 34914
rect 26462 34850 26514 34862
rect 31278 34850 31330 34862
rect 32958 34914 33010 34926
rect 32958 34850 33010 34862
rect 33742 34914 33794 34926
rect 33742 34850 33794 34862
rect 33966 34914 34018 34926
rect 40014 34914 40066 34926
rect 35746 34862 35758 34914
rect 35810 34862 35822 34914
rect 33966 34850 34018 34862
rect 40014 34850 40066 34862
rect 40462 34914 40514 34926
rect 50318 34914 50370 34926
rect 42578 34862 42590 34914
rect 42642 34862 42654 34914
rect 42914 34862 42926 34914
rect 42978 34862 42990 34914
rect 46050 34862 46062 34914
rect 46114 34862 46126 34914
rect 47618 34862 47630 34914
rect 47682 34862 47694 34914
rect 47842 34862 47854 34914
rect 47906 34862 47918 34914
rect 49410 34862 49422 34914
rect 49474 34862 49486 34914
rect 50530 34862 50542 34914
rect 50594 34862 50606 34914
rect 54562 34862 54574 34914
rect 54626 34862 54638 34914
rect 55458 34862 55470 34914
rect 55522 34862 55534 34914
rect 57138 34862 57150 34914
rect 57202 34862 57214 34914
rect 40462 34850 40514 34862
rect 50318 34850 50370 34862
rect 12126 34802 12178 34814
rect 7746 34750 7758 34802
rect 7810 34750 7822 34802
rect 9650 34750 9662 34802
rect 9714 34750 9726 34802
rect 12126 34738 12178 34750
rect 13022 34802 13074 34814
rect 13022 34738 13074 34750
rect 13806 34802 13858 34814
rect 13806 34738 13858 34750
rect 14142 34802 14194 34814
rect 14142 34738 14194 34750
rect 18734 34802 18786 34814
rect 18734 34738 18786 34750
rect 19070 34802 19122 34814
rect 19070 34738 19122 34750
rect 19630 34802 19682 34814
rect 19630 34738 19682 34750
rect 21310 34802 21362 34814
rect 21310 34738 21362 34750
rect 21422 34802 21474 34814
rect 21422 34738 21474 34750
rect 21870 34802 21922 34814
rect 21870 34738 21922 34750
rect 23438 34802 23490 34814
rect 26350 34802 26402 34814
rect 25218 34750 25230 34802
rect 25282 34750 25294 34802
rect 23438 34738 23490 34750
rect 26350 34738 26402 34750
rect 27246 34802 27298 34814
rect 27246 34738 27298 34750
rect 27582 34802 27634 34814
rect 27582 34738 27634 34750
rect 28366 34802 28418 34814
rect 28366 34738 28418 34750
rect 29374 34802 29426 34814
rect 29374 34738 29426 34750
rect 29710 34802 29762 34814
rect 29710 34738 29762 34750
rect 32734 34802 32786 34814
rect 32734 34738 32786 34750
rect 33294 34802 33346 34814
rect 33294 34738 33346 34750
rect 37102 34802 37154 34814
rect 37102 34738 37154 34750
rect 37326 34802 37378 34814
rect 37326 34738 37378 34750
rect 37886 34802 37938 34814
rect 37886 34738 37938 34750
rect 39566 34802 39618 34814
rect 39566 34738 39618 34750
rect 41022 34802 41074 34814
rect 49870 34802 49922 34814
rect 44930 34750 44942 34802
rect 44994 34750 45006 34802
rect 46834 34750 46846 34802
rect 46898 34750 46910 34802
rect 41022 34738 41074 34750
rect 49870 34738 49922 34750
rect 51550 34802 51602 34814
rect 56142 34802 56194 34814
rect 54226 34750 54238 34802
rect 54290 34750 54302 34802
rect 51550 34738 51602 34750
rect 56142 34738 56194 34750
rect 57598 34802 57650 34814
rect 57598 34738 57650 34750
rect 4622 34690 4674 34702
rect 4622 34626 4674 34638
rect 26126 34690 26178 34702
rect 26126 34626 26178 34638
rect 32846 34690 32898 34702
rect 32846 34626 32898 34638
rect 33854 34690 33906 34702
rect 33854 34626 33906 34638
rect 34190 34690 34242 34702
rect 34190 34626 34242 34638
rect 34862 34690 34914 34702
rect 34862 34626 34914 34638
rect 36430 34690 36482 34702
rect 36430 34626 36482 34638
rect 37550 34690 37602 34702
rect 37550 34626 37602 34638
rect 37774 34690 37826 34702
rect 51662 34690 51714 34702
rect 38434 34638 38446 34690
rect 38498 34638 38510 34690
rect 37774 34626 37826 34638
rect 51662 34626 51714 34638
rect 51886 34690 51938 34702
rect 51886 34626 51938 34638
rect 1344 34522 58731 34556
rect 1344 34470 15520 34522
rect 15572 34470 15624 34522
rect 15676 34470 15728 34522
rect 15780 34470 29827 34522
rect 29879 34470 29931 34522
rect 29983 34470 30035 34522
rect 30087 34470 44134 34522
rect 44186 34470 44238 34522
rect 44290 34470 44342 34522
rect 44394 34470 58441 34522
rect 58493 34470 58545 34522
rect 58597 34470 58649 34522
rect 58701 34470 58731 34522
rect 1344 34436 58731 34470
rect 2718 34354 2770 34366
rect 2718 34290 2770 34302
rect 4062 34354 4114 34366
rect 4062 34290 4114 34302
rect 5406 34354 5458 34366
rect 5406 34290 5458 34302
rect 6638 34354 6690 34366
rect 6638 34290 6690 34302
rect 6974 34354 7026 34366
rect 6974 34290 7026 34302
rect 7870 34354 7922 34366
rect 7870 34290 7922 34302
rect 8766 34354 8818 34366
rect 8766 34290 8818 34302
rect 9886 34354 9938 34366
rect 9886 34290 9938 34302
rect 11902 34354 11954 34366
rect 11902 34290 11954 34302
rect 17838 34354 17890 34366
rect 17838 34290 17890 34302
rect 20414 34354 20466 34366
rect 20414 34290 20466 34302
rect 21758 34354 21810 34366
rect 21758 34290 21810 34302
rect 24222 34354 24274 34366
rect 24222 34290 24274 34302
rect 28814 34354 28866 34366
rect 30942 34354 30994 34366
rect 29362 34302 29374 34354
rect 29426 34302 29438 34354
rect 28814 34290 28866 34302
rect 30942 34290 30994 34302
rect 33182 34354 33234 34366
rect 33182 34290 33234 34302
rect 36542 34354 36594 34366
rect 36542 34290 36594 34302
rect 36766 34354 36818 34366
rect 48190 34354 48242 34366
rect 42690 34302 42702 34354
rect 42754 34302 42766 34354
rect 36766 34290 36818 34302
rect 48190 34290 48242 34302
rect 50542 34354 50594 34366
rect 50542 34290 50594 34302
rect 55134 34354 55186 34366
rect 55134 34290 55186 34302
rect 3054 34242 3106 34254
rect 3054 34178 3106 34190
rect 3502 34242 3554 34254
rect 3502 34178 3554 34190
rect 4622 34242 4674 34254
rect 4622 34178 4674 34190
rect 16606 34242 16658 34254
rect 16606 34178 16658 34190
rect 21534 34242 21586 34254
rect 21534 34178 21586 34190
rect 22094 34242 22146 34254
rect 22094 34178 22146 34190
rect 28254 34242 28306 34254
rect 28254 34178 28306 34190
rect 33518 34242 33570 34254
rect 33518 34178 33570 34190
rect 35310 34242 35362 34254
rect 40014 34242 40066 34254
rect 37986 34190 37998 34242
rect 38050 34190 38062 34242
rect 35310 34178 35362 34190
rect 40014 34178 40066 34190
rect 43710 34242 43762 34254
rect 43710 34178 43762 34190
rect 45166 34242 45218 34254
rect 45166 34178 45218 34190
rect 48862 34242 48914 34254
rect 48862 34178 48914 34190
rect 49086 34242 49138 34254
rect 49086 34178 49138 34190
rect 49422 34242 49474 34254
rect 49422 34178 49474 34190
rect 50430 34242 50482 34254
rect 50430 34178 50482 34190
rect 54686 34242 54738 34254
rect 54686 34178 54738 34190
rect 56590 34242 56642 34254
rect 56590 34178 56642 34190
rect 1710 34130 1762 34142
rect 1710 34066 1762 34078
rect 3390 34130 3442 34142
rect 3390 34066 3442 34078
rect 3726 34130 3778 34142
rect 3726 34066 3778 34078
rect 4174 34130 4226 34142
rect 4174 34066 4226 34078
rect 4398 34130 4450 34142
rect 4398 34066 4450 34078
rect 4734 34130 4786 34142
rect 4734 34066 4786 34078
rect 7310 34130 7362 34142
rect 7310 34066 7362 34078
rect 8206 34130 8258 34142
rect 8206 34066 8258 34078
rect 10222 34130 10274 34142
rect 16270 34130 16322 34142
rect 12786 34078 12798 34130
rect 12850 34078 12862 34130
rect 10222 34066 10274 34078
rect 16270 34066 16322 34078
rect 18958 34130 19010 34142
rect 19854 34130 19906 34142
rect 19506 34078 19518 34130
rect 19570 34078 19582 34130
rect 18958 34066 19010 34078
rect 19854 34066 19906 34078
rect 20302 34130 20354 34142
rect 20302 34066 20354 34078
rect 20526 34130 20578 34142
rect 20526 34066 20578 34078
rect 20974 34130 21026 34142
rect 20974 34066 21026 34078
rect 21758 34130 21810 34142
rect 23998 34130 24050 34142
rect 31502 34130 31554 34142
rect 36878 34130 36930 34142
rect 39566 34130 39618 34142
rect 23090 34078 23102 34130
rect 23154 34078 23166 34130
rect 24546 34078 24558 34130
rect 24610 34078 24622 34130
rect 25666 34078 25678 34130
rect 25730 34078 25742 34130
rect 27570 34078 27582 34130
rect 27634 34078 27646 34130
rect 32162 34078 32174 34130
rect 32226 34078 32238 34130
rect 34738 34078 34750 34130
rect 34802 34078 34814 34130
rect 35970 34078 35982 34130
rect 36034 34078 36046 34130
rect 38210 34078 38222 34130
rect 38274 34078 38286 34130
rect 39106 34078 39118 34130
rect 39170 34078 39182 34130
rect 21758 34066 21810 34078
rect 23998 34066 24050 34078
rect 31502 34066 31554 34078
rect 36878 34066 36930 34078
rect 39566 34066 39618 34078
rect 40126 34130 40178 34142
rect 40126 34066 40178 34078
rect 41022 34130 41074 34142
rect 46286 34130 46338 34142
rect 47742 34130 47794 34142
rect 41570 34078 41582 34130
rect 41634 34078 41646 34130
rect 44146 34078 44158 34130
rect 44210 34078 44222 34130
rect 47058 34078 47070 34130
rect 47122 34078 47134 34130
rect 47506 34078 47518 34130
rect 47570 34078 47582 34130
rect 41022 34066 41074 34078
rect 46286 34066 46338 34078
rect 47742 34066 47794 34078
rect 48750 34130 48802 34142
rect 48750 34066 48802 34078
rect 49534 34130 49586 34142
rect 50654 34130 50706 34142
rect 53342 34130 53394 34142
rect 54574 34130 54626 34142
rect 50082 34078 50094 34130
rect 50146 34078 50158 34130
rect 51538 34078 51550 34130
rect 51602 34078 51614 34130
rect 52882 34078 52894 34130
rect 52946 34078 52958 34130
rect 54226 34078 54238 34130
rect 54290 34078 54302 34130
rect 49534 34066 49586 34078
rect 50654 34066 50706 34078
rect 53342 34066 53394 34078
rect 54574 34066 54626 34078
rect 56702 34130 56754 34142
rect 57250 34078 57262 34130
rect 57314 34078 57326 34130
rect 56702 34066 56754 34078
rect 10670 34018 10722 34030
rect 2146 33966 2158 34018
rect 2210 33966 2222 34018
rect 5842 33966 5854 34018
rect 5906 33966 5918 34018
rect 10670 33954 10722 33966
rect 11118 34018 11170 34030
rect 11118 33954 11170 33966
rect 12350 34018 12402 34030
rect 18286 34018 18338 34030
rect 13458 33966 13470 34018
rect 13522 33966 13534 34018
rect 15586 33966 15598 34018
rect 15650 33966 15662 34018
rect 12350 33954 12402 33966
rect 18286 33954 18338 33966
rect 18734 34018 18786 34030
rect 18734 33954 18786 33966
rect 22430 34018 22482 34030
rect 24110 34018 24162 34030
rect 26910 34018 26962 34030
rect 29934 34018 29986 34030
rect 23314 33966 23326 34018
rect 23378 33966 23390 34018
rect 24546 33966 24558 34018
rect 24610 34015 24622 34018
rect 24770 34015 24782 34018
rect 24610 33969 24782 34015
rect 24610 33966 24622 33969
rect 24770 33966 24782 33969
rect 24834 33966 24846 34018
rect 26002 33966 26014 34018
rect 26066 33966 26078 34018
rect 27906 33966 27918 34018
rect 27970 33966 27982 34018
rect 22430 33954 22482 33966
rect 24110 33954 24162 33966
rect 26910 33954 26962 33966
rect 29934 33954 29986 33966
rect 30494 34018 30546 34030
rect 33966 34018 34018 34030
rect 40910 34018 40962 34030
rect 58158 34018 58210 34030
rect 32386 33966 32398 34018
rect 32450 33966 32462 34018
rect 34066 33966 34078 34018
rect 34130 33966 34142 34018
rect 36194 33966 36206 34018
rect 36258 33966 36270 34018
rect 51090 33966 51102 34018
rect 51154 33966 51166 34018
rect 30494 33954 30546 33966
rect 33966 33954 34018 33966
rect 40910 33954 40962 33966
rect 58158 33954 58210 33966
rect 4062 33906 4114 33918
rect 29710 33906 29762 33918
rect 25330 33854 25342 33906
rect 25394 33854 25406 33906
rect 4062 33842 4114 33854
rect 29710 33842 29762 33854
rect 40014 33906 40066 33918
rect 40014 33842 40066 33854
rect 49422 33906 49474 33918
rect 49422 33842 49474 33854
rect 1344 33738 58576 33772
rect 1344 33686 8367 33738
rect 8419 33686 8471 33738
rect 8523 33686 8575 33738
rect 8627 33686 22674 33738
rect 22726 33686 22778 33738
rect 22830 33686 22882 33738
rect 22934 33686 36981 33738
rect 37033 33686 37085 33738
rect 37137 33686 37189 33738
rect 37241 33686 51288 33738
rect 51340 33686 51392 33738
rect 51444 33686 51496 33738
rect 51548 33686 58576 33738
rect 1344 33652 58576 33686
rect 35422 33570 35474 33582
rect 35422 33506 35474 33518
rect 50766 33570 50818 33582
rect 50766 33506 50818 33518
rect 51214 33570 51266 33582
rect 51214 33506 51266 33518
rect 54462 33570 54514 33582
rect 54462 33506 54514 33518
rect 6190 33458 6242 33470
rect 11566 33458 11618 33470
rect 4610 33406 4622 33458
rect 4674 33406 4686 33458
rect 8194 33406 8206 33458
rect 8258 33406 8270 33458
rect 6190 33394 6242 33406
rect 11566 33394 11618 33406
rect 12014 33458 12066 33470
rect 12014 33394 12066 33406
rect 12574 33458 12626 33470
rect 12574 33394 12626 33406
rect 12910 33458 12962 33470
rect 12910 33394 12962 33406
rect 14366 33458 14418 33470
rect 15710 33458 15762 33470
rect 20302 33458 20354 33470
rect 14914 33406 14926 33458
rect 14978 33406 14990 33458
rect 16818 33406 16830 33458
rect 16882 33406 16894 33458
rect 18946 33406 18958 33458
rect 19010 33406 19022 33458
rect 14366 33394 14418 33406
rect 15710 33394 15762 33406
rect 20302 33394 20354 33406
rect 21982 33458 22034 33470
rect 21982 33394 22034 33406
rect 26126 33458 26178 33470
rect 26126 33394 26178 33406
rect 27918 33458 27970 33470
rect 27918 33394 27970 33406
rect 28254 33458 28306 33470
rect 33966 33458 34018 33470
rect 39006 33458 39058 33470
rect 43822 33458 43874 33470
rect 48862 33458 48914 33470
rect 28578 33406 28590 33458
rect 28642 33406 28654 33458
rect 29586 33406 29598 33458
rect 29650 33406 29662 33458
rect 30146 33406 30158 33458
rect 30210 33406 30222 33458
rect 38546 33406 38558 33458
rect 38610 33406 38622 33458
rect 41234 33406 41246 33458
rect 41298 33406 41310 33458
rect 45378 33406 45390 33458
rect 45442 33406 45454 33458
rect 46722 33406 46734 33458
rect 46786 33406 46798 33458
rect 28254 33394 28306 33406
rect 33966 33394 34018 33406
rect 39006 33394 39058 33406
rect 43822 33394 43874 33406
rect 48862 33394 48914 33406
rect 53118 33458 53170 33470
rect 55794 33406 55806 33458
rect 55858 33406 55870 33458
rect 57586 33406 57598 33458
rect 57650 33406 57662 33458
rect 53118 33394 53170 33406
rect 20190 33346 20242 33358
rect 1810 33294 1822 33346
rect 1874 33294 1886 33346
rect 11106 33294 11118 33346
rect 11170 33294 11182 33346
rect 15250 33294 15262 33346
rect 15314 33294 15326 33346
rect 16146 33294 16158 33346
rect 16210 33294 16222 33346
rect 19842 33294 19854 33346
rect 19906 33294 19918 33346
rect 20190 33282 20242 33294
rect 21198 33346 21250 33358
rect 21198 33282 21250 33294
rect 21534 33346 21586 33358
rect 24894 33346 24946 33358
rect 23202 33294 23214 33346
rect 23266 33294 23278 33346
rect 24098 33294 24110 33346
rect 24162 33294 24174 33346
rect 21534 33282 21586 33294
rect 24894 33282 24946 33294
rect 25230 33346 25282 33358
rect 34302 33346 34354 33358
rect 27234 33294 27246 33346
rect 27298 33294 27310 33346
rect 27682 33294 27694 33346
rect 27746 33294 27758 33346
rect 29474 33294 29486 33346
rect 29538 33294 29550 33346
rect 30482 33294 30494 33346
rect 30546 33294 30558 33346
rect 32610 33294 32622 33346
rect 32674 33294 32686 33346
rect 33394 33294 33406 33346
rect 33458 33294 33470 33346
rect 25230 33282 25282 33294
rect 34302 33282 34354 33294
rect 34974 33346 35026 33358
rect 34974 33282 35026 33294
rect 35534 33346 35586 33358
rect 39118 33346 39170 33358
rect 43934 33346 43986 33358
rect 37090 33294 37102 33346
rect 37154 33294 37166 33346
rect 37650 33294 37662 33346
rect 37714 33294 37726 33346
rect 39442 33294 39454 33346
rect 39506 33294 39518 33346
rect 40562 33294 40574 33346
rect 40626 33294 40638 33346
rect 42690 33294 42702 33346
rect 42754 33294 42766 33346
rect 35534 33282 35586 33294
rect 39118 33282 39170 33294
rect 43934 33282 43986 33294
rect 44382 33346 44434 33358
rect 46286 33346 46338 33358
rect 49198 33346 49250 33358
rect 49758 33346 49810 33358
rect 45154 33294 45166 33346
rect 45218 33294 45230 33346
rect 48178 33294 48190 33346
rect 48242 33294 48254 33346
rect 49522 33294 49534 33346
rect 49586 33294 49598 33346
rect 44382 33282 44434 33294
rect 46286 33282 46338 33294
rect 49198 33282 49250 33294
rect 49758 33282 49810 33294
rect 50094 33346 50146 33358
rect 53230 33346 53282 33358
rect 53790 33346 53842 33358
rect 50754 33294 50766 33346
rect 50818 33294 50830 33346
rect 53554 33294 53566 33346
rect 53618 33294 53630 33346
rect 56018 33294 56030 33346
rect 56082 33294 56094 33346
rect 57922 33294 57934 33346
rect 57986 33294 57998 33346
rect 50094 33282 50146 33294
rect 53230 33282 53282 33294
rect 53790 33282 53842 33294
rect 13582 33234 13634 33246
rect 2482 33182 2494 33234
rect 2546 33182 2558 33234
rect 10322 33182 10334 33234
rect 10386 33182 10398 33234
rect 13582 33170 13634 33182
rect 13918 33234 13970 33246
rect 34526 33234 34578 33246
rect 22754 33182 22766 33234
rect 22818 33182 22830 33234
rect 32162 33182 32174 33234
rect 32226 33182 32238 33234
rect 13918 33170 13970 33182
rect 34526 33170 34578 33182
rect 35422 33234 35474 33246
rect 35422 33170 35474 33182
rect 40350 33234 40402 33246
rect 43374 33234 43426 33246
rect 41682 33182 41694 33234
rect 41746 33182 41758 33234
rect 40350 33170 40402 33182
rect 43374 33170 43426 33182
rect 43710 33234 43762 33246
rect 43710 33170 43762 33182
rect 45838 33234 45890 33246
rect 45838 33170 45890 33182
rect 46174 33234 46226 33246
rect 49982 33234 50034 33246
rect 47282 33182 47294 33234
rect 47346 33182 47358 33234
rect 46174 33170 46226 33182
rect 49982 33170 50034 33182
rect 50430 33234 50482 33246
rect 50430 33170 50482 33182
rect 51214 33234 51266 33246
rect 51214 33170 51266 33182
rect 51326 33234 51378 33246
rect 51326 33170 51378 33182
rect 54126 33234 54178 33246
rect 54126 33170 54178 33182
rect 54574 33234 54626 33246
rect 54574 33170 54626 33182
rect 5182 33122 5234 33134
rect 5182 33058 5234 33070
rect 5854 33122 5906 33134
rect 5854 33058 5906 33070
rect 6638 33122 6690 33134
rect 6638 33058 6690 33070
rect 7086 33122 7138 33134
rect 7086 33058 7138 33070
rect 7534 33122 7586 33134
rect 7534 33058 7586 33070
rect 20862 33122 20914 33134
rect 20862 33058 20914 33070
rect 21422 33122 21474 33134
rect 25118 33122 25170 33134
rect 24322 33070 24334 33122
rect 24386 33070 24398 33122
rect 21422 33058 21474 33070
rect 25118 33058 25170 33070
rect 25678 33122 25730 33134
rect 25678 33058 25730 33070
rect 26574 33122 26626 33134
rect 26574 33058 26626 33070
rect 28478 33122 28530 33134
rect 28478 33058 28530 33070
rect 30942 33122 30994 33134
rect 30942 33058 30994 33070
rect 34638 33122 34690 33134
rect 34638 33058 34690 33070
rect 36430 33122 36482 33134
rect 36430 33058 36482 33070
rect 40798 33122 40850 33134
rect 40798 33058 40850 33070
rect 40910 33122 40962 33134
rect 40910 33058 40962 33070
rect 49310 33122 49362 33134
rect 49310 33058 49362 33070
rect 51774 33122 51826 33134
rect 51774 33058 51826 33070
rect 53006 33122 53058 33134
rect 53006 33058 53058 33070
rect 54014 33122 54066 33134
rect 54014 33058 54066 33070
rect 1344 32954 58731 32988
rect 1344 32902 15520 32954
rect 15572 32902 15624 32954
rect 15676 32902 15728 32954
rect 15780 32902 29827 32954
rect 29879 32902 29931 32954
rect 29983 32902 30035 32954
rect 30087 32902 44134 32954
rect 44186 32902 44238 32954
rect 44290 32902 44342 32954
rect 44394 32902 58441 32954
rect 58493 32902 58545 32954
rect 58597 32902 58649 32954
rect 58701 32902 58731 32954
rect 1344 32868 58731 32902
rect 2494 32786 2546 32798
rect 2494 32722 2546 32734
rect 7198 32786 7250 32798
rect 7198 32722 7250 32734
rect 8878 32786 8930 32798
rect 8878 32722 8930 32734
rect 9662 32786 9714 32798
rect 9662 32722 9714 32734
rect 11790 32786 11842 32798
rect 11790 32722 11842 32734
rect 15262 32786 15314 32798
rect 20190 32786 20242 32798
rect 23886 32786 23938 32798
rect 17714 32734 17726 32786
rect 17778 32734 17790 32786
rect 23202 32734 23214 32786
rect 23266 32734 23278 32786
rect 15262 32722 15314 32734
rect 20190 32722 20242 32734
rect 23886 32722 23938 32734
rect 24446 32786 24498 32798
rect 24446 32722 24498 32734
rect 27694 32786 27746 32798
rect 27694 32722 27746 32734
rect 29822 32786 29874 32798
rect 29822 32722 29874 32734
rect 33294 32786 33346 32798
rect 33294 32722 33346 32734
rect 38782 32786 38834 32798
rect 38782 32722 38834 32734
rect 42814 32786 42866 32798
rect 42814 32722 42866 32734
rect 43934 32786 43986 32798
rect 56142 32786 56194 32798
rect 53218 32734 53230 32786
rect 53282 32734 53294 32786
rect 43934 32722 43986 32734
rect 56142 32722 56194 32734
rect 58158 32786 58210 32798
rect 58158 32722 58210 32734
rect 1822 32674 1874 32686
rect 1822 32610 1874 32622
rect 1934 32674 1986 32686
rect 1934 32610 1986 32622
rect 2382 32674 2434 32686
rect 2382 32610 2434 32622
rect 2718 32674 2770 32686
rect 2718 32610 2770 32622
rect 6638 32674 6690 32686
rect 6638 32610 6690 32622
rect 6750 32674 6802 32686
rect 16158 32674 16210 32686
rect 26238 32674 26290 32686
rect 7970 32622 7982 32674
rect 8034 32622 8046 32674
rect 8306 32622 8318 32674
rect 8370 32622 8382 32674
rect 10770 32622 10782 32674
rect 10834 32622 10846 32674
rect 18946 32622 18958 32674
rect 19010 32622 19022 32674
rect 21746 32622 21758 32674
rect 21810 32622 21822 32674
rect 23090 32622 23102 32674
rect 23154 32622 23166 32674
rect 6750 32610 6802 32622
rect 16158 32610 16210 32622
rect 26238 32610 26290 32622
rect 30382 32674 30434 32686
rect 30382 32610 30434 32622
rect 30606 32674 30658 32686
rect 30606 32610 30658 32622
rect 34414 32674 34466 32686
rect 34414 32610 34466 32622
rect 36318 32674 36370 32686
rect 36318 32610 36370 32622
rect 36542 32674 36594 32686
rect 38670 32674 38722 32686
rect 36978 32622 36990 32674
rect 37042 32622 37054 32674
rect 36542 32610 36594 32622
rect 38670 32610 38722 32622
rect 39342 32674 39394 32686
rect 39342 32610 39394 32622
rect 41918 32674 41970 32686
rect 41918 32610 41970 32622
rect 43822 32674 43874 32686
rect 43822 32610 43874 32622
rect 47854 32674 47906 32686
rect 47854 32610 47906 32622
rect 48750 32674 48802 32686
rect 54910 32674 54962 32686
rect 50530 32622 50542 32674
rect 50594 32622 50606 32674
rect 51986 32622 51998 32674
rect 52050 32622 52062 32674
rect 48750 32610 48802 32622
rect 54910 32610 54962 32622
rect 55806 32674 55858 32686
rect 55806 32610 55858 32622
rect 55918 32674 55970 32686
rect 55918 32610 55970 32622
rect 56590 32674 56642 32686
rect 56590 32610 56642 32622
rect 2158 32562 2210 32574
rect 2158 32498 2210 32510
rect 2942 32562 2994 32574
rect 6414 32562 6466 32574
rect 3266 32510 3278 32562
rect 3330 32510 3342 32562
rect 2942 32498 2994 32510
rect 6414 32498 6466 32510
rect 8542 32562 8594 32574
rect 8542 32498 8594 32510
rect 9438 32562 9490 32574
rect 9438 32498 9490 32510
rect 9774 32562 9826 32574
rect 9774 32498 9826 32510
rect 10110 32562 10162 32574
rect 15150 32562 15202 32574
rect 10658 32510 10670 32562
rect 10722 32510 10734 32562
rect 13234 32510 13246 32562
rect 13298 32510 13310 32562
rect 14578 32510 14590 32562
rect 14642 32510 14654 32562
rect 10110 32498 10162 32510
rect 15150 32498 15202 32510
rect 15374 32562 15426 32574
rect 15374 32498 15426 32510
rect 15822 32562 15874 32574
rect 26126 32562 26178 32574
rect 28926 32562 28978 32574
rect 18050 32510 18062 32562
rect 18114 32510 18126 32562
rect 28578 32510 28590 32562
rect 28642 32510 28654 32562
rect 15822 32498 15874 32510
rect 26126 32498 26178 32510
rect 28926 32498 28978 32510
rect 29374 32562 29426 32574
rect 29374 32498 29426 32510
rect 30270 32562 30322 32574
rect 30270 32498 30322 32510
rect 30830 32562 30882 32574
rect 32286 32562 32338 32574
rect 31826 32510 31838 32562
rect 31890 32510 31902 32562
rect 30830 32498 30882 32510
rect 32286 32498 32338 32510
rect 33070 32562 33122 32574
rect 33070 32498 33122 32510
rect 33182 32562 33234 32574
rect 33182 32498 33234 32510
rect 34302 32562 34354 32574
rect 34302 32498 34354 32510
rect 36654 32562 36706 32574
rect 39118 32562 39170 32574
rect 37426 32510 37438 32562
rect 37490 32510 37502 32562
rect 38434 32510 38446 32562
rect 38498 32510 38510 32562
rect 36654 32498 36706 32510
rect 39118 32498 39170 32510
rect 39454 32562 39506 32574
rect 39454 32498 39506 32510
rect 40350 32562 40402 32574
rect 40350 32498 40402 32510
rect 41470 32562 41522 32574
rect 41470 32498 41522 32510
rect 42030 32562 42082 32574
rect 42030 32498 42082 32510
rect 43374 32562 43426 32574
rect 43374 32498 43426 32510
rect 44046 32562 44098 32574
rect 46622 32562 46674 32574
rect 44818 32510 44830 32562
rect 44882 32510 44894 32562
rect 46274 32510 46286 32562
rect 46338 32510 46350 32562
rect 48066 32510 48078 32562
rect 48130 32510 48142 32562
rect 49410 32510 49422 32562
rect 49474 32510 49486 32562
rect 52882 32510 52894 32562
rect 52946 32510 52958 32562
rect 54226 32510 54238 32562
rect 54290 32510 54302 32562
rect 57474 32510 57486 32562
rect 57538 32510 57550 32562
rect 44046 32498 44098 32510
rect 46622 32498 46674 32510
rect 11454 32450 11506 32462
rect 16830 32450 16882 32462
rect 20750 32450 20802 32462
rect 4050 32398 4062 32450
rect 4114 32398 4126 32450
rect 6178 32398 6190 32450
rect 6242 32398 6254 32450
rect 14690 32398 14702 32450
rect 14754 32398 14766 32450
rect 16034 32398 16046 32450
rect 16098 32398 16110 32450
rect 19506 32398 19518 32450
rect 19570 32398 19582 32450
rect 11454 32386 11506 32398
rect 16830 32386 16882 32398
rect 20750 32386 20802 32398
rect 21422 32450 21474 32462
rect 21422 32386 21474 32398
rect 28030 32450 28082 32462
rect 28030 32386 28082 32398
rect 28254 32450 28306 32462
rect 40238 32450 40290 32462
rect 31378 32398 31390 32450
rect 31442 32398 31454 32450
rect 37762 32398 37774 32450
rect 37826 32398 37838 32450
rect 28254 32386 28306 32398
rect 40238 32386 40290 32398
rect 40910 32450 40962 32462
rect 40910 32386 40962 32398
rect 43262 32450 43314 32462
rect 45390 32450 45442 32462
rect 44482 32398 44494 32450
rect 44546 32398 44558 32450
rect 43262 32386 43314 32398
rect 45390 32386 45442 32398
rect 46734 32450 46786 32462
rect 46734 32386 46786 32398
rect 47182 32450 47234 32462
rect 55470 32450 55522 32462
rect 50866 32398 50878 32450
rect 50930 32398 50942 32450
rect 51426 32398 51438 32450
rect 51490 32398 51502 32450
rect 54002 32398 54014 32450
rect 54066 32398 54078 32450
rect 57138 32398 57150 32450
rect 57202 32398 57214 32450
rect 47182 32386 47234 32398
rect 55470 32386 55522 32398
rect 16382 32338 16434 32350
rect 13010 32286 13022 32338
rect 13074 32286 13086 32338
rect 16382 32274 16434 32286
rect 26238 32338 26290 32350
rect 26238 32274 26290 32286
rect 29150 32338 29202 32350
rect 29150 32274 29202 32286
rect 34414 32338 34466 32350
rect 34414 32274 34466 32286
rect 38782 32338 38834 32350
rect 38782 32274 38834 32286
rect 41246 32338 41298 32350
rect 41246 32274 41298 32286
rect 41918 32338 41970 32350
rect 41918 32274 41970 32286
rect 1344 32170 58576 32204
rect 1344 32118 8367 32170
rect 8419 32118 8471 32170
rect 8523 32118 8575 32170
rect 8627 32118 22674 32170
rect 22726 32118 22778 32170
rect 22830 32118 22882 32170
rect 22934 32118 36981 32170
rect 37033 32118 37085 32170
rect 37137 32118 37189 32170
rect 37241 32118 51288 32170
rect 51340 32118 51392 32170
rect 51444 32118 51496 32170
rect 51548 32118 58576 32170
rect 1344 32084 58576 32118
rect 32398 32002 32450 32014
rect 32398 31938 32450 31950
rect 33406 32002 33458 32014
rect 37426 31950 37438 32002
rect 37490 31950 37502 32002
rect 46946 31950 46958 32002
rect 47010 31950 47022 32002
rect 53330 31950 53342 32002
rect 53394 31950 53406 32002
rect 55794 31950 55806 32002
rect 55858 31950 55870 32002
rect 33406 31938 33458 31950
rect 7198 31890 7250 31902
rect 7198 31826 7250 31838
rect 7534 31890 7586 31902
rect 21534 31890 21586 31902
rect 18498 31838 18510 31890
rect 18562 31838 18574 31890
rect 20178 31838 20190 31890
rect 20242 31838 20254 31890
rect 7534 31826 7586 31838
rect 21534 31826 21586 31838
rect 27134 31890 27186 31902
rect 33854 31890 33906 31902
rect 31826 31838 31838 31890
rect 31890 31838 31902 31890
rect 27134 31826 27186 31838
rect 33854 31826 33906 31838
rect 36430 31890 36482 31902
rect 43710 31890 43762 31902
rect 37762 31838 37774 31890
rect 37826 31838 37838 31890
rect 36430 31826 36482 31838
rect 43710 31826 43762 31838
rect 45726 31890 45778 31902
rect 45726 31826 45778 31838
rect 51326 31890 51378 31902
rect 53666 31838 53678 31890
rect 53730 31838 53742 31890
rect 51326 31826 51378 31838
rect 2270 31778 2322 31790
rect 1810 31726 1822 31778
rect 1874 31726 1886 31778
rect 2270 31714 2322 31726
rect 3838 31778 3890 31790
rect 3838 31714 3890 31726
rect 3950 31778 4002 31790
rect 3950 31714 4002 31726
rect 5966 31778 6018 31790
rect 5966 31714 6018 31726
rect 8430 31778 8482 31790
rect 8430 31714 8482 31726
rect 9550 31778 9602 31790
rect 9550 31714 9602 31726
rect 10670 31778 10722 31790
rect 10670 31714 10722 31726
rect 14254 31778 14306 31790
rect 15150 31778 15202 31790
rect 16158 31778 16210 31790
rect 14802 31726 14814 31778
rect 14866 31726 14878 31778
rect 15810 31726 15822 31778
rect 15874 31726 15886 31778
rect 14254 31714 14306 31726
rect 15150 31714 15202 31726
rect 16158 31714 16210 31726
rect 16494 31778 16546 31790
rect 16494 31714 16546 31726
rect 17054 31778 17106 31790
rect 19742 31778 19794 31790
rect 25902 31778 25954 31790
rect 18274 31726 18286 31778
rect 18338 31726 18350 31778
rect 19394 31726 19406 31778
rect 19458 31726 19470 31778
rect 20290 31726 20302 31778
rect 20354 31726 20366 31778
rect 17054 31714 17106 31726
rect 19742 31714 19794 31726
rect 25902 31714 25954 31726
rect 26238 31778 26290 31790
rect 27358 31778 27410 31790
rect 26562 31726 26574 31778
rect 26626 31726 26638 31778
rect 26238 31714 26290 31726
rect 27358 31714 27410 31726
rect 27694 31778 27746 31790
rect 33294 31778 33346 31790
rect 34750 31778 34802 31790
rect 30146 31726 30158 31778
rect 30210 31726 30222 31778
rect 34514 31726 34526 31778
rect 34578 31726 34590 31778
rect 27694 31714 27746 31726
rect 33294 31714 33346 31726
rect 34750 31714 34802 31726
rect 35534 31778 35586 31790
rect 39678 31778 39730 31790
rect 40574 31778 40626 31790
rect 35970 31726 35982 31778
rect 36034 31726 36046 31778
rect 37874 31726 37886 31778
rect 37938 31726 37950 31778
rect 40114 31726 40126 31778
rect 40178 31726 40190 31778
rect 35534 31714 35586 31726
rect 39678 31714 39730 31726
rect 40574 31714 40626 31726
rect 41022 31778 41074 31790
rect 41022 31714 41074 31726
rect 41358 31778 41410 31790
rect 42702 31778 42754 31790
rect 42466 31726 42478 31778
rect 42530 31726 42542 31778
rect 41358 31714 41410 31726
rect 42702 31714 42754 31726
rect 44718 31778 44770 31790
rect 44718 31714 44770 31726
rect 45054 31778 45106 31790
rect 45054 31714 45106 31726
rect 45614 31778 45666 31790
rect 55134 31778 55186 31790
rect 56926 31778 56978 31790
rect 46162 31726 46174 31778
rect 46226 31726 46238 31778
rect 48178 31726 48190 31778
rect 48242 31726 48254 31778
rect 49074 31726 49086 31778
rect 49138 31726 49150 31778
rect 51986 31726 51998 31778
rect 52050 31726 52062 31778
rect 53554 31726 53566 31778
rect 53618 31726 53630 31778
rect 54674 31726 54686 31778
rect 54738 31726 54750 31778
rect 54898 31726 54910 31778
rect 54962 31726 54974 31778
rect 56018 31726 56030 31778
rect 56082 31726 56094 31778
rect 57250 31726 57262 31778
rect 57314 31726 57326 31778
rect 45614 31714 45666 31726
rect 55134 31714 55186 31726
rect 56926 31714 56978 31726
rect 3278 31666 3330 31678
rect 3278 31602 3330 31614
rect 4286 31666 4338 31678
rect 4286 31602 4338 31614
rect 4622 31666 4674 31678
rect 4622 31602 4674 31614
rect 4958 31666 5010 31678
rect 4958 31602 5010 31614
rect 5630 31666 5682 31678
rect 5630 31602 5682 31614
rect 5742 31666 5794 31678
rect 8318 31666 8370 31678
rect 6626 31614 6638 31666
rect 6690 31614 6702 31666
rect 6962 31614 6974 31666
rect 7026 31614 7038 31666
rect 5742 31602 5794 31614
rect 8318 31602 8370 31614
rect 9214 31666 9266 31678
rect 9214 31602 9266 31614
rect 9326 31666 9378 31678
rect 16382 31666 16434 31678
rect 15586 31614 15598 31666
rect 15650 31614 15662 31666
rect 9326 31602 9378 31614
rect 16382 31602 16434 31614
rect 17390 31666 17442 31678
rect 25566 31666 25618 31678
rect 32734 31666 32786 31678
rect 18722 31614 18734 31666
rect 18786 31614 18798 31666
rect 21634 31614 21646 31666
rect 21698 31614 21710 31666
rect 23314 31614 23326 31666
rect 23378 31614 23390 31666
rect 29138 31614 29150 31666
rect 29202 31614 29214 31666
rect 31490 31614 31502 31666
rect 31554 31614 31566 31666
rect 17390 31602 17442 31614
rect 25566 31602 25618 31614
rect 32734 31602 32786 31614
rect 33406 31666 33458 31678
rect 41134 31666 41186 31678
rect 38882 31614 38894 31666
rect 38946 31614 38958 31666
rect 33406 31602 33458 31614
rect 41134 31602 41186 31614
rect 42926 31666 42978 31678
rect 42926 31602 42978 31614
rect 44942 31666 44994 31678
rect 47058 31614 47070 31666
rect 47122 31614 47134 31666
rect 48066 31614 48078 31666
rect 48130 31614 48142 31666
rect 50082 31614 50094 31666
rect 50146 31614 50158 31666
rect 44942 31602 44994 31614
rect 2718 31554 2770 31566
rect 2718 31490 2770 31502
rect 2942 31554 2994 31566
rect 2942 31490 2994 31502
rect 3166 31554 3218 31566
rect 3166 31490 3218 31502
rect 4062 31554 4114 31566
rect 4062 31490 4114 31502
rect 8094 31554 8146 31566
rect 8094 31490 8146 31502
rect 8878 31554 8930 31566
rect 8878 31490 8930 31502
rect 9886 31554 9938 31566
rect 9886 31490 9938 31502
rect 10334 31554 10386 31566
rect 10334 31490 10386 31502
rect 10782 31554 10834 31566
rect 10782 31490 10834 31502
rect 11006 31554 11058 31566
rect 11006 31490 11058 31502
rect 17278 31554 17330 31566
rect 17278 31490 17330 31502
rect 17950 31554 18002 31566
rect 24110 31554 24162 31566
rect 23202 31502 23214 31554
rect 23266 31502 23278 31554
rect 17950 31490 18002 31502
rect 24110 31490 24162 31502
rect 24334 31554 24386 31566
rect 24334 31490 24386 31502
rect 24446 31554 24498 31566
rect 24446 31490 24498 31502
rect 24558 31554 24610 31566
rect 24558 31490 24610 31502
rect 25678 31554 25730 31566
rect 25678 31490 25730 31502
rect 27582 31554 27634 31566
rect 27582 31490 27634 31502
rect 28590 31554 28642 31566
rect 28590 31490 28642 31502
rect 32510 31554 32562 31566
rect 32510 31490 32562 31502
rect 39230 31554 39282 31566
rect 39230 31490 39282 31502
rect 43598 31554 43650 31566
rect 43598 31490 43650 31502
rect 43822 31554 43874 31566
rect 43822 31490 43874 31502
rect 44046 31554 44098 31566
rect 44046 31490 44098 31502
rect 50878 31554 50930 31566
rect 50878 31490 50930 31502
rect 51774 31554 51826 31566
rect 51774 31490 51826 31502
rect 1344 31386 58731 31420
rect 1344 31334 15520 31386
rect 15572 31334 15624 31386
rect 15676 31334 15728 31386
rect 15780 31334 29827 31386
rect 29879 31334 29931 31386
rect 29983 31334 30035 31386
rect 30087 31334 44134 31386
rect 44186 31334 44238 31386
rect 44290 31334 44342 31386
rect 44394 31334 58441 31386
rect 58493 31334 58545 31386
rect 58597 31334 58649 31386
rect 58701 31334 58731 31386
rect 1344 31300 58731 31334
rect 15822 31218 15874 31230
rect 15822 31154 15874 31166
rect 16382 31218 16434 31230
rect 19294 31218 19346 31230
rect 18946 31166 18958 31218
rect 19010 31166 19022 31218
rect 16382 31154 16434 31166
rect 19294 31154 19346 31166
rect 19406 31218 19458 31230
rect 19406 31154 19458 31166
rect 20302 31218 20354 31230
rect 20302 31154 20354 31166
rect 21422 31218 21474 31230
rect 33182 31218 33234 31230
rect 45390 31218 45442 31230
rect 23874 31166 23886 31218
rect 23938 31166 23950 31218
rect 40002 31166 40014 31218
rect 40066 31166 40078 31218
rect 40898 31166 40910 31218
rect 40962 31166 40974 31218
rect 21422 31154 21474 31166
rect 33182 31154 33234 31166
rect 45390 31154 45442 31166
rect 15710 31106 15762 31118
rect 15710 31042 15762 31054
rect 19742 31106 19794 31118
rect 26014 31106 26066 31118
rect 22306 31054 22318 31106
rect 22370 31054 22382 31106
rect 23986 31054 23998 31106
rect 24050 31054 24062 31106
rect 19742 31042 19794 31054
rect 26014 31042 26066 31054
rect 28254 31106 28306 31118
rect 28254 31042 28306 31054
rect 33294 31106 33346 31118
rect 45502 31106 45554 31118
rect 55246 31106 55298 31118
rect 34738 31054 34750 31106
rect 34802 31054 34814 31106
rect 35186 31054 35198 31106
rect 35250 31054 35262 31106
rect 36306 31054 36318 31106
rect 36370 31054 36382 31106
rect 38658 31054 38670 31106
rect 38722 31054 38734 31106
rect 45938 31054 45950 31106
rect 46002 31054 46014 31106
rect 33294 31042 33346 31054
rect 45502 31042 45554 31054
rect 55246 31042 55298 31054
rect 56590 31106 56642 31118
rect 56590 31042 56642 31054
rect 58046 31106 58098 31118
rect 58046 31042 58098 31054
rect 1710 30994 1762 31006
rect 14814 30994 14866 31006
rect 2818 30942 2830 30994
rect 2882 30942 2894 30994
rect 6178 30942 6190 30994
rect 6242 30942 6254 30994
rect 10098 30942 10110 30994
rect 10162 30942 10174 30994
rect 1710 30930 1762 30942
rect 14814 30930 14866 30942
rect 15038 30994 15090 31006
rect 15038 30930 15090 30942
rect 15486 30994 15538 31006
rect 15486 30930 15538 30942
rect 19518 30994 19570 31006
rect 19518 30930 19570 30942
rect 20414 30994 20466 31006
rect 26910 30994 26962 31006
rect 34078 30994 34130 31006
rect 40350 30994 40402 31006
rect 45166 30994 45218 31006
rect 22866 30942 22878 30994
rect 22930 30942 22942 30994
rect 26674 30942 26686 30994
rect 26738 30942 26750 30994
rect 29138 30942 29150 30994
rect 29202 30942 29214 30994
rect 29810 30942 29822 30994
rect 29874 30942 29886 30994
rect 31602 30942 31614 30994
rect 31666 30942 31678 30994
rect 37538 30942 37550 30994
rect 37602 30942 37614 30994
rect 42578 30942 42590 30994
rect 42642 30942 42654 30994
rect 43922 30942 43934 30994
rect 43986 30942 43998 30994
rect 46386 30942 46398 30994
rect 46450 30942 46462 30994
rect 46722 30942 46734 30994
rect 46786 30942 46798 30994
rect 47954 30942 47966 30994
rect 48018 30942 48030 30994
rect 49074 30942 49086 30994
rect 49138 30942 49150 30994
rect 49410 30942 49422 30994
rect 49474 30942 49486 30994
rect 51650 30942 51662 30994
rect 51714 30942 51726 30994
rect 52994 30942 53006 30994
rect 53058 30942 53070 30994
rect 53778 30942 53790 30994
rect 53842 30942 53854 30994
rect 55458 30942 55470 30994
rect 55522 30942 55534 30994
rect 57026 30942 57038 30994
rect 57090 30942 57102 30994
rect 20414 30930 20466 30942
rect 26910 30930 26962 30942
rect 34078 30930 34130 30942
rect 40350 30930 40402 30942
rect 45166 30930 45218 30942
rect 2270 30882 2322 30894
rect 9662 30882 9714 30894
rect 14926 30882 14978 30894
rect 3602 30830 3614 30882
rect 3666 30830 3678 30882
rect 5730 30830 5742 30882
rect 5794 30830 5806 30882
rect 6850 30830 6862 30882
rect 6914 30830 6926 30882
rect 8978 30830 8990 30882
rect 9042 30830 9054 30882
rect 10770 30830 10782 30882
rect 10834 30830 10846 30882
rect 12898 30830 12910 30882
rect 12962 30830 12974 30882
rect 2270 30818 2322 30830
rect 9662 30818 9714 30830
rect 14926 30818 14978 30830
rect 17614 30882 17666 30894
rect 17614 30818 17666 30830
rect 18398 30882 18450 30894
rect 18398 30818 18450 30830
rect 20862 30882 20914 30894
rect 20862 30818 20914 30830
rect 28366 30882 28418 30894
rect 30606 30882 30658 30894
rect 32286 30882 32338 30894
rect 28914 30830 28926 30882
rect 28978 30830 28990 30882
rect 29362 30830 29374 30882
rect 29426 30830 29438 30882
rect 31826 30830 31838 30882
rect 31890 30830 31902 30882
rect 28366 30818 28418 30830
rect 30606 30818 30658 30830
rect 32286 30818 32338 30830
rect 33070 30882 33122 30894
rect 33070 30818 33122 30830
rect 34414 30882 34466 30894
rect 41470 30882 41522 30894
rect 56142 30882 56194 30894
rect 36082 30830 36094 30882
rect 36146 30830 36158 30882
rect 42466 30830 42478 30882
rect 42530 30830 42542 30882
rect 48850 30830 48862 30882
rect 48914 30830 48926 30882
rect 49298 30830 49310 30882
rect 49362 30830 49374 30882
rect 51762 30830 51774 30882
rect 51826 30830 51838 30882
rect 54226 30830 54238 30882
rect 54290 30830 54302 30882
rect 57362 30830 57374 30882
rect 57426 30830 57438 30882
rect 34414 30818 34466 30830
rect 41470 30818 41522 30830
rect 56142 30818 56194 30830
rect 15822 30770 15874 30782
rect 15822 30706 15874 30718
rect 18622 30770 18674 30782
rect 18622 30706 18674 30718
rect 28478 30770 28530 30782
rect 28478 30706 28530 30718
rect 41246 30770 41298 30782
rect 44482 30718 44494 30770
rect 44546 30718 44558 30770
rect 50754 30718 50766 30770
rect 50818 30718 50830 30770
rect 41246 30706 41298 30718
rect 1344 30602 58576 30636
rect 1344 30550 8367 30602
rect 8419 30550 8471 30602
rect 8523 30550 8575 30602
rect 8627 30550 22674 30602
rect 22726 30550 22778 30602
rect 22830 30550 22882 30602
rect 22934 30550 36981 30602
rect 37033 30550 37085 30602
rect 37137 30550 37189 30602
rect 37241 30550 51288 30602
rect 51340 30550 51392 30602
rect 51444 30550 51496 30602
rect 51548 30550 58576 30602
rect 1344 30516 58576 30550
rect 19630 30434 19682 30446
rect 6962 30382 6974 30434
rect 7026 30431 7038 30434
rect 7298 30431 7310 30434
rect 7026 30385 7310 30431
rect 7026 30382 7038 30385
rect 7298 30382 7310 30385
rect 7362 30382 7374 30434
rect 19630 30370 19682 30382
rect 19966 30434 20018 30446
rect 19966 30370 20018 30382
rect 23998 30434 24050 30446
rect 23998 30370 24050 30382
rect 31726 30434 31778 30446
rect 55346 30382 55358 30434
rect 55410 30382 55422 30434
rect 31726 30370 31778 30382
rect 10670 30322 10722 30334
rect 10670 30258 10722 30270
rect 16606 30322 16658 30334
rect 21534 30322 21586 30334
rect 34078 30322 34130 30334
rect 40686 30322 40738 30334
rect 18498 30270 18510 30322
rect 18562 30270 18574 30322
rect 24546 30270 24558 30322
rect 24610 30270 24622 30322
rect 27682 30270 27694 30322
rect 27746 30270 27758 30322
rect 38546 30270 38558 30322
rect 38610 30270 38622 30322
rect 16606 30258 16658 30270
rect 21534 30258 21586 30270
rect 34078 30258 34130 30270
rect 40686 30258 40738 30270
rect 43038 30322 43090 30334
rect 45826 30270 45838 30322
rect 45890 30270 45902 30322
rect 48962 30270 48974 30322
rect 49026 30270 49038 30322
rect 54450 30270 54462 30322
rect 54514 30270 54526 30322
rect 57138 30270 57150 30322
rect 57202 30270 57214 30322
rect 43038 30258 43090 30270
rect 2942 30210 2994 30222
rect 2942 30146 2994 30158
rect 3614 30210 3666 30222
rect 3614 30146 3666 30158
rect 4398 30210 4450 30222
rect 4398 30146 4450 30158
rect 5630 30210 5682 30222
rect 5630 30146 5682 30158
rect 5966 30210 6018 30222
rect 5966 30146 6018 30158
rect 7534 30210 7586 30222
rect 7534 30146 7586 30158
rect 7870 30210 7922 30222
rect 7870 30146 7922 30158
rect 9998 30210 10050 30222
rect 9998 30146 10050 30158
rect 10558 30210 10610 30222
rect 28590 30210 28642 30222
rect 11330 30158 11342 30210
rect 11394 30158 11406 30210
rect 15026 30158 15038 30210
rect 15090 30158 15102 30210
rect 18834 30158 18846 30210
rect 18898 30158 18910 30210
rect 26002 30158 26014 30210
rect 26066 30158 26078 30210
rect 27906 30158 27918 30210
rect 27970 30158 27982 30210
rect 10558 30146 10610 30158
rect 28590 30146 28642 30158
rect 29150 30210 29202 30222
rect 29150 30146 29202 30158
rect 29486 30210 29538 30222
rect 29486 30146 29538 30158
rect 30046 30210 30098 30222
rect 30046 30146 30098 30158
rect 31390 30210 31442 30222
rect 31390 30146 31442 30158
rect 32398 30210 32450 30222
rect 32398 30146 32450 30158
rect 33182 30210 33234 30222
rect 37662 30210 37714 30222
rect 33618 30158 33630 30210
rect 33682 30158 33694 30210
rect 40002 30158 40014 30210
rect 40066 30158 40078 30210
rect 43474 30158 43486 30210
rect 43538 30158 43550 30210
rect 44258 30158 44270 30210
rect 44322 30158 44334 30210
rect 47170 30158 47182 30210
rect 47234 30158 47246 30210
rect 50418 30158 50430 30210
rect 50482 30158 50494 30210
rect 52658 30158 52670 30210
rect 52722 30158 52734 30210
rect 53218 30158 53230 30210
rect 53282 30158 53294 30210
rect 55682 30158 55694 30210
rect 55746 30158 55758 30210
rect 56690 30158 56702 30210
rect 56754 30158 56766 30210
rect 57922 30158 57934 30210
rect 57986 30158 57998 30210
rect 33182 30146 33234 30158
rect 37662 30146 37714 30158
rect 1710 30098 1762 30110
rect 1710 30034 1762 30046
rect 2046 30098 2098 30110
rect 2046 30034 2098 30046
rect 4734 30098 4786 30110
rect 4734 30034 4786 30046
rect 4958 30098 5010 30110
rect 4958 30034 5010 30046
rect 6414 30098 6466 30110
rect 6414 30034 6466 30046
rect 6638 30098 6690 30110
rect 6638 30034 6690 30046
rect 6750 30098 6802 30110
rect 6750 30034 6802 30046
rect 8094 30098 8146 30110
rect 8094 30034 8146 30046
rect 10222 30098 10274 30110
rect 10222 30034 10274 30046
rect 10782 30098 10834 30110
rect 10782 30034 10834 30046
rect 11118 30098 11170 30110
rect 19294 30098 19346 30110
rect 14914 30046 14926 30098
rect 14978 30046 14990 30098
rect 16370 30046 16382 30098
rect 16434 30046 16446 30098
rect 11118 30034 11170 30046
rect 19294 30034 19346 30046
rect 20190 30098 20242 30110
rect 23886 30098 23938 30110
rect 29374 30098 29426 30110
rect 21634 30046 21646 30098
rect 21698 30046 21710 30098
rect 23314 30046 23326 30098
rect 23378 30046 23390 30098
rect 24770 30046 24782 30098
rect 24834 30046 24846 30098
rect 20190 30034 20242 30046
rect 23886 30034 23938 30046
rect 29374 30034 29426 30046
rect 31614 30098 31666 30110
rect 31614 30034 31666 30046
rect 36990 30098 37042 30110
rect 36990 30034 37042 30046
rect 37214 30098 37266 30110
rect 54126 30098 54178 30110
rect 38770 30046 38782 30098
rect 38834 30046 38846 30098
rect 42802 30046 42814 30098
rect 42866 30046 42878 30098
rect 46274 30046 46286 30098
rect 46338 30046 46350 30098
rect 48514 30046 48526 30098
rect 48578 30046 48590 30098
rect 49410 30046 49422 30098
rect 49474 30046 49486 30098
rect 53330 30046 53342 30098
rect 53394 30046 53406 30098
rect 37214 30034 37266 30046
rect 54126 30034 54178 30046
rect 57598 30098 57650 30110
rect 57598 30034 57650 30046
rect 2382 29986 2434 29998
rect 2382 29922 2434 29934
rect 3726 29986 3778 29998
rect 3726 29922 3778 29934
rect 3950 29986 4002 29998
rect 3950 29922 4002 29934
rect 4510 29986 4562 29998
rect 4510 29922 4562 29934
rect 5742 29986 5794 29998
rect 5742 29922 5794 29934
rect 7198 29986 7250 29998
rect 7198 29922 7250 29934
rect 7646 29986 7698 29998
rect 7646 29922 7698 29934
rect 8542 29986 8594 29998
rect 8542 29922 8594 29934
rect 13694 29986 13746 29998
rect 13694 29922 13746 29934
rect 17054 29986 17106 29998
rect 23998 29986 24050 29998
rect 37326 29986 37378 29998
rect 23202 29934 23214 29986
rect 23266 29934 23278 29986
rect 26562 29934 26574 29986
rect 26626 29934 26638 29986
rect 17054 29922 17106 29934
rect 23998 29922 24050 29934
rect 37326 29922 37378 29934
rect 45166 29986 45218 29998
rect 45166 29922 45218 29934
rect 51774 29986 51826 29998
rect 54350 29986 54402 29998
rect 52770 29934 52782 29986
rect 52834 29934 52846 29986
rect 51774 29922 51826 29934
rect 54350 29922 54402 29934
rect 57710 29986 57762 29998
rect 57710 29922 57762 29934
rect 1344 29818 58731 29852
rect 1344 29766 15520 29818
rect 15572 29766 15624 29818
rect 15676 29766 15728 29818
rect 15780 29766 29827 29818
rect 29879 29766 29931 29818
rect 29983 29766 30035 29818
rect 30087 29766 44134 29818
rect 44186 29766 44238 29818
rect 44290 29766 44342 29818
rect 44394 29766 58441 29818
rect 58493 29766 58545 29818
rect 58597 29766 58649 29818
rect 58701 29766 58731 29818
rect 1344 29732 58731 29766
rect 19966 29650 20018 29662
rect 13794 29598 13806 29650
rect 13858 29598 13870 29650
rect 19966 29586 20018 29598
rect 20526 29650 20578 29662
rect 20526 29586 20578 29598
rect 20750 29650 20802 29662
rect 20750 29586 20802 29598
rect 21534 29650 21586 29662
rect 21534 29586 21586 29598
rect 25678 29650 25730 29662
rect 31950 29650 32002 29662
rect 29250 29598 29262 29650
rect 29314 29598 29326 29650
rect 25678 29586 25730 29598
rect 31950 29586 32002 29598
rect 32062 29650 32114 29662
rect 32062 29586 32114 29598
rect 32398 29650 32450 29662
rect 32398 29586 32450 29598
rect 35534 29650 35586 29662
rect 35534 29586 35586 29598
rect 42926 29650 42978 29662
rect 42926 29586 42978 29598
rect 47966 29650 48018 29662
rect 47966 29586 48018 29598
rect 48078 29650 48130 29662
rect 48962 29598 48974 29650
rect 49026 29598 49038 29650
rect 48078 29586 48130 29598
rect 15374 29538 15426 29550
rect 20190 29538 20242 29550
rect 18162 29486 18174 29538
rect 18226 29486 18238 29538
rect 15374 29474 15426 29486
rect 20190 29474 20242 29486
rect 20862 29538 20914 29550
rect 20862 29474 20914 29486
rect 21310 29538 21362 29550
rect 21310 29474 21362 29486
rect 23662 29538 23714 29550
rect 29934 29538 29986 29550
rect 28018 29486 28030 29538
rect 28082 29486 28094 29538
rect 23662 29474 23714 29486
rect 29934 29474 29986 29486
rect 34526 29538 34578 29550
rect 34526 29474 34578 29486
rect 34638 29538 34690 29550
rect 34638 29474 34690 29486
rect 35422 29538 35474 29550
rect 35422 29474 35474 29486
rect 36990 29538 37042 29550
rect 36990 29474 37042 29486
rect 42814 29538 42866 29550
rect 42814 29474 42866 29486
rect 45726 29538 45778 29550
rect 54350 29538 54402 29550
rect 50194 29486 50206 29538
rect 50258 29486 50270 29538
rect 51538 29486 51550 29538
rect 51602 29486 51614 29538
rect 53778 29486 53790 29538
rect 53842 29486 53854 29538
rect 45726 29474 45778 29486
rect 54350 29474 54402 29486
rect 55806 29538 55858 29550
rect 55806 29474 55858 29486
rect 55918 29538 55970 29550
rect 56914 29486 56926 29538
rect 56978 29486 56990 29538
rect 55918 29474 55970 29486
rect 19742 29426 19794 29438
rect 1810 29374 1822 29426
rect 1874 29374 1886 29426
rect 5282 29374 5294 29426
rect 5346 29374 5358 29426
rect 10210 29374 10222 29426
rect 10274 29374 10286 29426
rect 13570 29374 13582 29426
rect 13634 29374 13646 29426
rect 14690 29374 14702 29426
rect 14754 29374 14766 29426
rect 19282 29374 19294 29426
rect 19346 29374 19358 29426
rect 19742 29362 19794 29374
rect 20302 29426 20354 29438
rect 20302 29362 20354 29374
rect 21198 29426 21250 29438
rect 21198 29362 21250 29374
rect 23774 29426 23826 29438
rect 32174 29426 32226 29438
rect 38222 29426 38274 29438
rect 54574 29426 54626 29438
rect 56142 29426 56194 29438
rect 24322 29374 24334 29426
rect 24386 29374 24398 29426
rect 29026 29374 29038 29426
rect 29090 29374 29102 29426
rect 30594 29374 30606 29426
rect 30658 29374 30670 29426
rect 31602 29374 31614 29426
rect 31666 29374 31678 29426
rect 33618 29374 33630 29426
rect 33682 29374 33694 29426
rect 36530 29374 36542 29426
rect 36594 29374 36606 29426
rect 37762 29374 37774 29426
rect 37826 29374 37838 29426
rect 39890 29374 39902 29426
rect 39954 29374 39966 29426
rect 44146 29374 44158 29426
rect 44210 29374 44222 29426
rect 45266 29374 45278 29426
rect 45330 29374 45342 29426
rect 50082 29374 50094 29426
rect 50146 29374 50158 29426
rect 52994 29374 53006 29426
rect 53058 29374 53070 29426
rect 54786 29374 54798 29426
rect 54850 29374 54862 29426
rect 56578 29374 56590 29426
rect 56642 29374 56654 29426
rect 57698 29374 57710 29426
rect 57762 29374 57774 29426
rect 23774 29362 23826 29374
rect 32174 29362 32226 29374
rect 38222 29362 38274 29374
rect 54574 29362 54626 29374
rect 56142 29362 56194 29374
rect 17726 29314 17778 29326
rect 2594 29262 2606 29314
rect 2658 29262 2670 29314
rect 4722 29262 4734 29314
rect 4786 29262 4798 29314
rect 6066 29262 6078 29314
rect 6130 29262 6142 29314
rect 8194 29262 8206 29314
rect 8258 29262 8270 29314
rect 10882 29262 10894 29314
rect 10946 29262 10958 29314
rect 13010 29262 13022 29314
rect 13074 29262 13086 29314
rect 14914 29262 14926 29314
rect 14978 29262 14990 29314
rect 17726 29250 17778 29262
rect 21870 29314 21922 29326
rect 21870 29250 21922 29262
rect 25790 29314 25842 29326
rect 31390 29314 31442 29326
rect 34078 29314 34130 29326
rect 37326 29314 37378 29326
rect 40350 29314 40402 29326
rect 46174 29314 46226 29326
rect 58158 29314 58210 29326
rect 27458 29262 27470 29314
rect 27522 29262 27534 29314
rect 30258 29262 30270 29314
rect 30322 29262 30334 29314
rect 33282 29262 33294 29314
rect 33346 29262 33358 29314
rect 36082 29262 36094 29314
rect 36146 29262 36158 29314
rect 39554 29262 39566 29314
rect 39618 29262 39630 29314
rect 43922 29262 43934 29314
rect 43986 29262 43998 29314
rect 44930 29262 44942 29314
rect 44994 29262 45006 29314
rect 51202 29262 51214 29314
rect 51266 29262 51278 29314
rect 57138 29262 57150 29314
rect 57202 29262 57214 29314
rect 25790 29250 25842 29262
rect 31390 29250 31442 29262
rect 34078 29250 34130 29262
rect 37326 29250 37378 29262
rect 40350 29250 40402 29262
rect 46174 29250 46226 29262
rect 58158 29250 58210 29262
rect 31278 29202 31330 29214
rect 31278 29138 31330 29150
rect 34526 29202 34578 29214
rect 34526 29138 34578 29150
rect 35646 29202 35698 29214
rect 48190 29202 48242 29214
rect 43586 29150 43598 29202
rect 43650 29150 43662 29202
rect 35646 29138 35698 29150
rect 48190 29138 48242 29150
rect 1344 29034 58576 29068
rect 1344 28982 8367 29034
rect 8419 28982 8471 29034
rect 8523 28982 8575 29034
rect 8627 28982 22674 29034
rect 22726 28982 22778 29034
rect 22830 28982 22882 29034
rect 22934 28982 36981 29034
rect 37033 28982 37085 29034
rect 37137 28982 37189 29034
rect 37241 28982 51288 29034
rect 51340 28982 51392 29034
rect 51444 28982 51496 29034
rect 51548 28982 58576 29034
rect 1344 28948 58576 28982
rect 8318 28866 8370 28878
rect 8318 28802 8370 28814
rect 8654 28866 8706 28878
rect 8654 28802 8706 28814
rect 9886 28866 9938 28878
rect 9886 28802 9938 28814
rect 12798 28866 12850 28878
rect 21982 28866 22034 28878
rect 14914 28814 14926 28866
rect 14978 28814 14990 28866
rect 12798 28802 12850 28814
rect 21982 28802 22034 28814
rect 25118 28866 25170 28878
rect 25118 28802 25170 28814
rect 27918 28866 27970 28878
rect 27918 28802 27970 28814
rect 33854 28866 33906 28878
rect 43710 28866 43762 28878
rect 37426 28814 37438 28866
rect 37490 28863 37502 28866
rect 38210 28863 38222 28866
rect 37490 28817 38222 28863
rect 37490 28814 37502 28817
rect 38210 28814 38222 28817
rect 38274 28814 38286 28866
rect 33854 28802 33906 28814
rect 43710 28802 43762 28814
rect 44046 28866 44098 28878
rect 44046 28802 44098 28814
rect 44942 28866 44994 28878
rect 44942 28802 44994 28814
rect 49198 28866 49250 28878
rect 49198 28802 49250 28814
rect 55694 28866 55746 28878
rect 55694 28802 55746 28814
rect 3054 28754 3106 28766
rect 3054 28690 3106 28702
rect 5070 28754 5122 28766
rect 5070 28690 5122 28702
rect 5742 28754 5794 28766
rect 5742 28690 5794 28702
rect 10446 28754 10498 28766
rect 19742 28754 19794 28766
rect 15138 28702 15150 28754
rect 15202 28702 15214 28754
rect 10446 28690 10498 28702
rect 19742 28690 19794 28702
rect 20638 28754 20690 28766
rect 20638 28690 20690 28702
rect 23438 28754 23490 28766
rect 23438 28690 23490 28702
rect 24446 28754 24498 28766
rect 24446 28690 24498 28702
rect 24894 28754 24946 28766
rect 24894 28690 24946 28702
rect 25902 28754 25954 28766
rect 28478 28754 28530 28766
rect 27122 28702 27134 28754
rect 27186 28702 27198 28754
rect 25902 28690 25954 28702
rect 28478 28690 28530 28702
rect 30046 28754 30098 28766
rect 33294 28754 33346 28766
rect 30482 28702 30494 28754
rect 30546 28702 30558 28754
rect 31154 28702 31166 28754
rect 31218 28702 31230 28754
rect 30046 28690 30098 28702
rect 33294 28690 33346 28702
rect 37662 28754 37714 28766
rect 43374 28754 43426 28766
rect 50318 28754 50370 28766
rect 42690 28702 42702 28754
rect 42754 28702 42766 28754
rect 46386 28702 46398 28754
rect 46450 28702 46462 28754
rect 49746 28702 49758 28754
rect 49810 28702 49822 28754
rect 52770 28702 52782 28754
rect 52834 28702 52846 28754
rect 57922 28702 57934 28754
rect 57986 28702 57998 28754
rect 37662 28690 37714 28702
rect 43374 28690 43426 28702
rect 50318 28690 50370 28702
rect 1934 28642 1986 28654
rect 1934 28578 1986 28590
rect 2158 28642 2210 28654
rect 2158 28578 2210 28590
rect 2830 28642 2882 28654
rect 2830 28578 2882 28590
rect 3278 28642 3330 28654
rect 3278 28578 3330 28590
rect 3726 28642 3778 28654
rect 3726 28578 3778 28590
rect 4734 28642 4786 28654
rect 4734 28578 4786 28590
rect 5518 28642 5570 28654
rect 5518 28578 5570 28590
rect 5966 28642 6018 28654
rect 5966 28578 6018 28590
rect 6078 28642 6130 28654
rect 6078 28578 6130 28590
rect 6750 28642 6802 28654
rect 6750 28578 6802 28590
rect 9438 28642 9490 28654
rect 9438 28578 9490 28590
rect 10222 28642 10274 28654
rect 10222 28578 10274 28590
rect 10670 28642 10722 28654
rect 10670 28578 10722 28590
rect 11118 28642 11170 28654
rect 11118 28578 11170 28590
rect 11454 28642 11506 28654
rect 11454 28578 11506 28590
rect 11678 28642 11730 28654
rect 11678 28578 11730 28590
rect 12014 28642 12066 28654
rect 18846 28642 18898 28654
rect 21198 28642 21250 28654
rect 23326 28642 23378 28654
rect 33182 28642 33234 28654
rect 14242 28590 14254 28642
rect 14306 28590 14318 28642
rect 15362 28590 15374 28642
rect 15426 28590 15438 28642
rect 19058 28590 19070 28642
rect 19122 28590 19134 28642
rect 22978 28590 22990 28642
rect 23042 28590 23054 28642
rect 23986 28590 23998 28642
rect 24050 28590 24062 28642
rect 30594 28590 30606 28642
rect 30658 28590 30670 28642
rect 32834 28590 32846 28642
rect 32898 28590 32910 28642
rect 12014 28578 12066 28590
rect 18846 28578 18898 28590
rect 21198 28578 21250 28590
rect 23326 28578 23378 28590
rect 33182 28578 33234 28590
rect 33406 28642 33458 28654
rect 33406 28578 33458 28590
rect 33742 28642 33794 28654
rect 33742 28578 33794 28590
rect 35982 28642 36034 28654
rect 35982 28578 36034 28590
rect 36878 28642 36930 28654
rect 44270 28642 44322 28654
rect 38770 28590 38782 28642
rect 38834 28590 38846 28642
rect 39554 28590 39566 28642
rect 39618 28590 39630 28642
rect 40786 28590 40798 28642
rect 40850 28590 40862 28642
rect 41570 28590 41582 28642
rect 41634 28590 41646 28642
rect 36878 28578 36930 28590
rect 44270 28578 44322 28590
rect 45278 28642 45330 28654
rect 49982 28642 50034 28654
rect 55022 28642 55074 28654
rect 48178 28590 48190 28642
rect 48242 28590 48254 28642
rect 51426 28590 51438 28642
rect 51490 28590 51502 28642
rect 51874 28590 51886 28642
rect 51938 28590 51950 28642
rect 53218 28590 53230 28642
rect 53282 28590 53294 28642
rect 54562 28590 54574 28642
rect 54626 28590 54638 28642
rect 56354 28590 56366 28642
rect 56418 28590 56430 28642
rect 45278 28578 45330 28590
rect 49982 28578 50034 28590
rect 55022 28578 55074 28590
rect 2494 28530 2546 28542
rect 2494 28466 2546 28478
rect 3502 28530 3554 28542
rect 3502 28466 3554 28478
rect 3950 28530 4002 28542
rect 3950 28466 4002 28478
rect 4062 28530 4114 28542
rect 4062 28466 4114 28478
rect 4398 28530 4450 28542
rect 4398 28466 4450 28478
rect 6974 28530 7026 28542
rect 6974 28466 7026 28478
rect 7086 28530 7138 28542
rect 9998 28530 10050 28542
rect 7634 28478 7646 28530
rect 7698 28478 7710 28530
rect 7970 28478 7982 28530
rect 8034 28478 8046 28530
rect 7086 28466 7138 28478
rect 9998 28466 10050 28478
rect 10894 28530 10946 28542
rect 10894 28466 10946 28478
rect 12238 28530 12290 28542
rect 12238 28466 12290 28478
rect 12350 28530 12402 28542
rect 12350 28466 12402 28478
rect 12686 28530 12738 28542
rect 12686 28466 12738 28478
rect 12798 28530 12850 28542
rect 20190 28530 20242 28542
rect 14466 28478 14478 28530
rect 14530 28478 14542 28530
rect 12798 28466 12850 28478
rect 20190 28466 20242 28478
rect 21534 28530 21586 28542
rect 21534 28466 21586 28478
rect 21982 28530 22034 28542
rect 21982 28466 22034 28478
rect 22094 28530 22146 28542
rect 22094 28466 22146 28478
rect 24334 28530 24386 28542
rect 31502 28530 31554 28542
rect 27122 28478 27134 28530
rect 27186 28478 27198 28530
rect 24334 28466 24386 28478
rect 31502 28466 31554 28478
rect 36318 28530 36370 28542
rect 36318 28466 36370 28478
rect 37102 28530 37154 28542
rect 37102 28466 37154 28478
rect 37214 28530 37266 28542
rect 45054 28530 45106 28542
rect 39666 28478 39678 28530
rect 39730 28478 39742 28530
rect 40674 28478 40686 28530
rect 40738 28478 40750 28530
rect 37214 28466 37266 28478
rect 45054 28466 45106 28478
rect 45502 28530 45554 28542
rect 45502 28466 45554 28478
rect 45614 28530 45666 28542
rect 52110 28530 52162 28542
rect 46610 28478 46622 28530
rect 46674 28478 46686 28530
rect 57362 28478 57374 28530
rect 57426 28478 57438 28530
rect 45614 28466 45666 28478
rect 52110 28466 52162 28478
rect 4510 28418 4562 28430
rect 4510 28354 4562 28366
rect 9886 28418 9938 28430
rect 9886 28354 9938 28366
rect 11454 28418 11506 28430
rect 11454 28354 11506 28366
rect 13918 28418 13970 28430
rect 13918 28354 13970 28366
rect 21422 28418 21474 28430
rect 21422 28354 21474 28366
rect 24558 28418 24610 28430
rect 25790 28418 25842 28430
rect 25442 28366 25454 28418
rect 25506 28366 25518 28418
rect 24558 28354 24610 28366
rect 25790 28354 25842 28366
rect 31278 28418 31330 28430
rect 31278 28354 31330 28366
rect 34526 28418 34578 28430
rect 34526 28354 34578 28366
rect 35758 28418 35810 28430
rect 35758 28354 35810 28366
rect 36206 28418 36258 28430
rect 36206 28354 36258 28366
rect 38222 28418 38274 28430
rect 44942 28418 44994 28430
rect 38658 28366 38670 28418
rect 38722 28366 38734 28418
rect 38222 28354 38274 28366
rect 44942 28354 44994 28366
rect 1344 28250 58731 28284
rect 1344 28198 15520 28250
rect 15572 28198 15624 28250
rect 15676 28198 15728 28250
rect 15780 28198 29827 28250
rect 29879 28198 29931 28250
rect 29983 28198 30035 28250
rect 30087 28198 44134 28250
rect 44186 28198 44238 28250
rect 44290 28198 44342 28250
rect 44394 28198 58441 28250
rect 58493 28198 58545 28250
rect 58597 28198 58649 28250
rect 58701 28198 58731 28250
rect 1344 28164 58731 28198
rect 1710 28082 1762 28094
rect 4734 28082 4786 28094
rect 9550 28082 9602 28094
rect 2706 28030 2718 28082
rect 2770 28030 2782 28082
rect 3042 28030 3054 28082
rect 3106 28030 3118 28082
rect 7410 28030 7422 28082
rect 7474 28030 7486 28082
rect 1710 28018 1762 28030
rect 4734 28018 4786 28030
rect 9550 28018 9602 28030
rect 10334 28082 10386 28094
rect 10334 28018 10386 28030
rect 10782 28082 10834 28094
rect 10782 28018 10834 28030
rect 11006 28082 11058 28094
rect 18062 28082 18114 28094
rect 16482 28030 16494 28082
rect 16546 28030 16558 28082
rect 11006 28018 11058 28030
rect 18062 28018 18114 28030
rect 18510 28082 18562 28094
rect 18510 28018 18562 28030
rect 20526 28082 20578 28094
rect 20526 28018 20578 28030
rect 22318 28082 22370 28094
rect 22318 28018 22370 28030
rect 22542 28082 22594 28094
rect 22542 28018 22594 28030
rect 35422 28082 35474 28094
rect 35422 28018 35474 28030
rect 39902 28082 39954 28094
rect 39902 28018 39954 28030
rect 41022 28082 41074 28094
rect 41022 28018 41074 28030
rect 49310 28082 49362 28094
rect 49310 28018 49362 28030
rect 49534 28082 49586 28094
rect 52222 28082 52274 28094
rect 49746 28030 49758 28082
rect 49810 28030 49822 28082
rect 49534 28018 49586 28030
rect 52222 28018 52274 28030
rect 54238 28082 54290 28094
rect 54238 28018 54290 28030
rect 57262 28082 57314 28094
rect 57262 28018 57314 28030
rect 2046 27970 2098 27982
rect 2046 27906 2098 27918
rect 4286 27970 4338 27982
rect 4286 27906 4338 27918
rect 7982 27970 8034 27982
rect 18622 27970 18674 27982
rect 12114 27918 12126 27970
rect 12178 27918 12190 27970
rect 15250 27918 15262 27970
rect 15314 27918 15326 27970
rect 16594 27918 16606 27970
rect 16658 27918 16670 27970
rect 7982 27906 8034 27918
rect 18622 27906 18674 27918
rect 25454 27970 25506 27982
rect 25454 27906 25506 27918
rect 30270 27970 30322 27982
rect 40910 27970 40962 27982
rect 47294 27970 47346 27982
rect 32162 27918 32174 27970
rect 32226 27918 32238 27970
rect 37314 27918 37326 27970
rect 37378 27918 37390 27970
rect 39554 27918 39566 27970
rect 39618 27918 39630 27970
rect 42466 27918 42478 27970
rect 42530 27918 42542 27970
rect 30270 27906 30322 27918
rect 40910 27906 40962 27918
rect 47294 27906 47346 27918
rect 48190 27970 48242 27982
rect 52446 27970 52498 27982
rect 48190 27906 48242 27918
rect 49198 27914 49250 27926
rect 51874 27918 51886 27970
rect 51938 27918 51950 27970
rect 2382 27858 2434 27870
rect 7086 27858 7138 27870
rect 9886 27858 9938 27870
rect 3266 27806 3278 27858
rect 3330 27806 3342 27858
rect 4050 27806 4062 27858
rect 4114 27806 4126 27858
rect 8418 27806 8430 27858
rect 8482 27806 8494 27858
rect 2382 27794 2434 27806
rect 7086 27794 7138 27806
rect 9886 27794 9938 27806
rect 10670 27858 10722 27870
rect 18286 27858 18338 27870
rect 20302 27858 20354 27870
rect 22206 27858 22258 27870
rect 28030 27858 28082 27870
rect 34638 27858 34690 27870
rect 11442 27806 11454 27858
rect 11506 27806 11518 27858
rect 19394 27806 19406 27858
rect 19458 27806 19470 27858
rect 20850 27806 20862 27858
rect 20914 27806 20926 27858
rect 24210 27806 24222 27858
rect 24274 27806 24286 27858
rect 25890 27806 25902 27858
rect 25954 27806 25966 27858
rect 27682 27806 27694 27858
rect 27746 27806 27758 27858
rect 28802 27806 28814 27858
rect 28866 27806 28878 27858
rect 30930 27806 30942 27858
rect 30994 27806 31006 27858
rect 34178 27806 34190 27858
rect 34242 27806 34254 27858
rect 10670 27794 10722 27806
rect 18286 27794 18338 27806
rect 20302 27794 20354 27806
rect 22206 27794 22258 27806
rect 28030 27794 28082 27806
rect 34638 27794 34690 27806
rect 34974 27858 35026 27870
rect 34974 27794 35026 27806
rect 35310 27858 35362 27870
rect 35310 27794 35362 27806
rect 35646 27858 35698 27870
rect 43710 27858 43762 27870
rect 37426 27806 37438 27858
rect 37490 27806 37502 27858
rect 38210 27806 38222 27858
rect 38274 27806 38286 27858
rect 41234 27806 41246 27858
rect 41298 27806 41310 27858
rect 42690 27806 42702 27858
rect 42754 27806 42766 27858
rect 43362 27806 43374 27858
rect 43426 27806 43438 27858
rect 35646 27794 35698 27806
rect 43710 27794 43762 27806
rect 44270 27858 44322 27870
rect 45950 27858 46002 27870
rect 47630 27858 47682 27870
rect 45490 27806 45502 27858
rect 45554 27806 45566 27858
rect 46834 27806 46846 27858
rect 46898 27806 46910 27858
rect 44270 27794 44322 27806
rect 45950 27794 46002 27806
rect 47630 27794 47682 27806
rect 47854 27858 47906 27870
rect 47854 27794 47906 27806
rect 48078 27858 48130 27870
rect 52446 27906 52498 27918
rect 52558 27970 52610 27982
rect 52558 27906 52610 27918
rect 54126 27970 54178 27982
rect 54126 27906 54178 27918
rect 55022 27970 55074 27982
rect 55022 27906 55074 27918
rect 57822 27970 57874 27982
rect 57822 27906 57874 27918
rect 49198 27850 49250 27862
rect 50206 27858 50258 27870
rect 48078 27794 48130 27806
rect 50206 27794 50258 27806
rect 50318 27858 50370 27870
rect 53006 27858 53058 27870
rect 50530 27806 50542 27858
rect 50594 27806 50606 27858
rect 50866 27806 50878 27858
rect 50930 27806 50942 27858
rect 51426 27806 51438 27858
rect 51490 27806 51502 27858
rect 50318 27794 50370 27806
rect 53006 27794 53058 27806
rect 54350 27858 54402 27870
rect 54350 27794 54402 27806
rect 54686 27858 54738 27870
rect 54686 27794 54738 27806
rect 55134 27858 55186 27870
rect 55458 27806 55470 27858
rect 55522 27806 55534 27858
rect 57026 27806 57038 27858
rect 57090 27806 57102 27858
rect 55134 27794 55186 27806
rect 5182 27746 5234 27758
rect 5182 27682 5234 27694
rect 8990 27746 9042 27758
rect 14814 27746 14866 27758
rect 14242 27694 14254 27746
rect 14306 27694 14318 27746
rect 8990 27682 9042 27694
rect 14814 27682 14866 27694
rect 18958 27746 19010 27758
rect 20414 27746 20466 27758
rect 19842 27694 19854 27746
rect 19906 27694 19918 27746
rect 18958 27682 19010 27694
rect 20414 27682 20466 27694
rect 21758 27746 21810 27758
rect 21758 27682 21810 27694
rect 22878 27746 22930 27758
rect 24670 27746 24722 27758
rect 24322 27694 24334 27746
rect 24386 27694 24398 27746
rect 22878 27682 22930 27694
rect 24670 27682 24722 27694
rect 25230 27746 25282 27758
rect 28142 27746 28194 27758
rect 25554 27694 25566 27746
rect 25618 27694 25630 27746
rect 25230 27682 25282 27694
rect 28142 27682 28194 27694
rect 28478 27746 28530 27758
rect 28478 27682 28530 27694
rect 28590 27746 28642 27758
rect 28590 27682 28642 27694
rect 32286 27746 32338 27758
rect 40014 27746 40066 27758
rect 48862 27746 48914 27758
rect 52894 27746 52946 27758
rect 33730 27694 33742 27746
rect 33794 27694 33806 27746
rect 42354 27694 42366 27746
rect 42418 27694 42430 27746
rect 45042 27694 45054 27746
rect 45106 27694 45118 27746
rect 46946 27694 46958 27746
rect 47010 27694 47022 27746
rect 51538 27694 51550 27746
rect 51602 27694 51614 27746
rect 32286 27682 32338 27694
rect 40014 27682 40066 27694
rect 48862 27682 48914 27694
rect 52894 27682 52946 27694
rect 53902 27746 53954 27758
rect 57138 27694 57150 27746
rect 57202 27694 57214 27746
rect 57698 27694 57710 27746
rect 57762 27694 57774 27746
rect 53902 27682 53954 27694
rect 25902 27634 25954 27646
rect 4722 27582 4734 27634
rect 4786 27631 4798 27634
rect 5170 27631 5182 27634
rect 4786 27585 5182 27631
rect 4786 27582 4798 27585
rect 5170 27582 5182 27585
rect 5234 27582 5246 27634
rect 25902 27570 25954 27582
rect 26238 27634 26290 27646
rect 26238 27570 26290 27582
rect 58046 27634 58098 27646
rect 58046 27570 58098 27582
rect 1344 27466 58576 27500
rect 1344 27414 8367 27466
rect 8419 27414 8471 27466
rect 8523 27414 8575 27466
rect 8627 27414 22674 27466
rect 22726 27414 22778 27466
rect 22830 27414 22882 27466
rect 22934 27414 36981 27466
rect 37033 27414 37085 27466
rect 37137 27414 37189 27466
rect 37241 27414 51288 27466
rect 51340 27414 51392 27466
rect 51444 27414 51496 27466
rect 51548 27414 58576 27466
rect 1344 27380 58576 27414
rect 16494 27298 16546 27310
rect 16494 27234 16546 27246
rect 20078 27298 20130 27310
rect 20078 27234 20130 27246
rect 34414 27298 34466 27310
rect 46958 27298 47010 27310
rect 43810 27246 43822 27298
rect 43874 27246 43886 27298
rect 46610 27246 46622 27298
rect 46674 27246 46686 27298
rect 34414 27234 34466 27246
rect 46958 27234 47010 27246
rect 47294 27298 47346 27310
rect 47294 27234 47346 27246
rect 47742 27298 47794 27310
rect 47742 27234 47794 27246
rect 49086 27298 49138 27310
rect 49086 27234 49138 27246
rect 50654 27298 50706 27310
rect 50654 27234 50706 27246
rect 52782 27298 52834 27310
rect 57138 27246 57150 27298
rect 57202 27246 57214 27298
rect 52782 27234 52834 27246
rect 15598 27186 15650 27198
rect 4610 27134 4622 27186
rect 4674 27134 4686 27186
rect 8530 27134 8542 27186
rect 8594 27134 8606 27186
rect 15598 27122 15650 27134
rect 17278 27186 17330 27198
rect 17278 27122 17330 27134
rect 26014 27186 26066 27198
rect 31726 27186 31778 27198
rect 30930 27134 30942 27186
rect 30994 27134 31006 27186
rect 26014 27122 26066 27134
rect 31726 27122 31778 27134
rect 33854 27186 33906 27198
rect 33854 27122 33906 27134
rect 35646 27186 35698 27198
rect 37998 27186 38050 27198
rect 36306 27134 36318 27186
rect 36370 27134 36382 27186
rect 35646 27122 35698 27134
rect 37998 27122 38050 27134
rect 40014 27186 40066 27198
rect 40014 27122 40066 27134
rect 42926 27186 42978 27198
rect 52110 27186 52162 27198
rect 44930 27134 44942 27186
rect 44994 27134 45006 27186
rect 42926 27122 42978 27134
rect 52110 27122 52162 27134
rect 10894 27074 10946 27086
rect 1698 27022 1710 27074
rect 1762 27022 1774 27074
rect 5618 27022 5630 27074
rect 5682 27022 5694 27074
rect 10894 27010 10946 27022
rect 11230 27074 11282 27086
rect 11230 27010 11282 27022
rect 11790 27074 11842 27086
rect 11790 27010 11842 27022
rect 15486 27074 15538 27086
rect 15486 27010 15538 27022
rect 15710 27074 15762 27086
rect 15710 27010 15762 27022
rect 16158 27074 16210 27086
rect 16158 27010 16210 27022
rect 17838 27074 17890 27086
rect 17838 27010 17890 27022
rect 18062 27074 18114 27086
rect 18062 27010 18114 27022
rect 18398 27074 18450 27086
rect 18398 27010 18450 27022
rect 18622 27074 18674 27086
rect 18622 27010 18674 27022
rect 18846 27074 18898 27086
rect 18846 27010 18898 27022
rect 19742 27074 19794 27086
rect 19742 27010 19794 27022
rect 21982 27074 22034 27086
rect 21982 27010 22034 27022
rect 22206 27074 22258 27086
rect 22206 27010 22258 27022
rect 22542 27074 22594 27086
rect 22542 27010 22594 27022
rect 22990 27074 23042 27086
rect 24222 27074 24274 27086
rect 34078 27074 34130 27086
rect 23650 27022 23662 27074
rect 23714 27022 23726 27074
rect 27458 27022 27470 27074
rect 27522 27022 27534 27074
rect 31266 27022 31278 27074
rect 31330 27022 31342 27074
rect 22990 27010 23042 27022
rect 24222 27010 24274 27022
rect 34078 27010 34130 27022
rect 34638 27074 34690 27086
rect 37102 27074 37154 27086
rect 39678 27074 39730 27086
rect 36082 27022 36094 27074
rect 36146 27022 36158 27074
rect 37314 27022 37326 27074
rect 37378 27022 37390 27074
rect 34638 27010 34690 27022
rect 37102 27010 37154 27022
rect 39678 27010 39730 27022
rect 42030 27074 42082 27086
rect 43262 27074 43314 27086
rect 42242 27022 42254 27074
rect 42306 27022 42318 27074
rect 42030 27010 42082 27022
rect 43262 27010 43314 27022
rect 43486 27074 43538 27086
rect 43486 27010 43538 27022
rect 45390 27074 45442 27086
rect 45390 27010 45442 27022
rect 46062 27074 46114 27086
rect 46062 27010 46114 27022
rect 46286 27074 46338 27086
rect 46286 27010 46338 27022
rect 47854 27074 47906 27086
rect 47854 27010 47906 27022
rect 48526 27074 48578 27086
rect 57262 27074 57314 27086
rect 51538 27022 51550 27074
rect 51602 27022 51614 27074
rect 51874 27022 51886 27074
rect 51938 27022 51950 27074
rect 55122 27022 55134 27074
rect 55186 27022 55198 27074
rect 56018 27022 56030 27074
rect 56082 27022 56094 27074
rect 57474 27022 57486 27074
rect 57538 27022 57550 27074
rect 48526 27010 48578 27022
rect 57262 27010 57314 27022
rect 9998 26962 10050 26974
rect 2482 26910 2494 26962
rect 2546 26910 2558 26962
rect 6402 26910 6414 26962
rect 6466 26910 6478 26962
rect 9998 26898 10050 26910
rect 10334 26962 10386 26974
rect 10334 26898 10386 26910
rect 11566 26962 11618 26974
rect 11566 26898 11618 26910
rect 12014 26962 12066 26974
rect 12014 26898 12066 26910
rect 12126 26962 12178 26974
rect 12126 26898 12178 26910
rect 12686 26962 12738 26974
rect 12686 26898 12738 26910
rect 16382 26962 16434 26974
rect 16382 26898 16434 26910
rect 18174 26962 18226 26974
rect 18174 26898 18226 26910
rect 19518 26962 19570 26974
rect 19518 26898 19570 26910
rect 22654 26962 22706 26974
rect 22654 26898 22706 26910
rect 22878 26962 22930 26974
rect 22878 26898 22930 26910
rect 24334 26962 24386 26974
rect 29262 26962 29314 26974
rect 26226 26910 26238 26962
rect 26290 26910 26302 26962
rect 27906 26910 27918 26962
rect 27970 26910 27982 26962
rect 24334 26898 24386 26910
rect 29262 26898 29314 26910
rect 30494 26962 30546 26974
rect 30494 26898 30546 26910
rect 32062 26962 32114 26974
rect 32062 26898 32114 26910
rect 33294 26962 33346 26974
rect 33294 26898 33346 26910
rect 34302 26962 34354 26974
rect 34302 26898 34354 26910
rect 34862 26962 34914 26974
rect 34862 26898 34914 26910
rect 34974 26962 35026 26974
rect 34974 26898 35026 26910
rect 39790 26962 39842 26974
rect 39790 26898 39842 26910
rect 40126 26962 40178 26974
rect 40126 26898 40178 26910
rect 47182 26962 47234 26974
rect 47182 26898 47234 26910
rect 47742 26962 47794 26974
rect 47742 26898 47794 26910
rect 48190 26962 48242 26974
rect 48190 26898 48242 26910
rect 49198 26962 49250 26974
rect 49198 26898 49250 26910
rect 50542 26962 50594 26974
rect 52894 26962 52946 26974
rect 50542 26898 50594 26910
rect 50654 26906 50706 26918
rect 10670 26850 10722 26862
rect 10670 26786 10722 26798
rect 11230 26850 11282 26862
rect 11230 26786 11282 26798
rect 16494 26850 16546 26862
rect 21534 26850 21586 26862
rect 19170 26798 19182 26850
rect 19234 26798 19246 26850
rect 16494 26786 16546 26798
rect 21534 26786 21586 26798
rect 22318 26850 22370 26862
rect 22318 26786 22370 26798
rect 24782 26850 24834 26862
rect 24782 26786 24834 26798
rect 30046 26850 30098 26862
rect 30046 26786 30098 26798
rect 32174 26850 32226 26862
rect 32174 26786 32226 26798
rect 32398 26850 32450 26862
rect 32398 26786 32450 26798
rect 32846 26850 32898 26862
rect 32846 26786 32898 26798
rect 38894 26850 38946 26862
rect 38894 26786 38946 26798
rect 48302 26850 48354 26862
rect 48302 26786 48354 26798
rect 49086 26850 49138 26862
rect 49086 26786 49138 26798
rect 49870 26850 49922 26862
rect 52894 26898 52946 26910
rect 53342 26962 53394 26974
rect 53342 26898 53394 26910
rect 53454 26962 53506 26974
rect 53454 26898 53506 26910
rect 54126 26962 54178 26974
rect 56702 26962 56754 26974
rect 54786 26910 54798 26962
rect 54850 26910 54862 26962
rect 54126 26898 54178 26910
rect 56702 26898 56754 26910
rect 50654 26842 50706 26854
rect 52782 26850 52834 26862
rect 49870 26786 49922 26798
rect 52782 26786 52834 26798
rect 53678 26850 53730 26862
rect 53678 26786 53730 26798
rect 1344 26682 58731 26716
rect 1344 26630 15520 26682
rect 15572 26630 15624 26682
rect 15676 26630 15728 26682
rect 15780 26630 29827 26682
rect 29879 26630 29931 26682
rect 29983 26630 30035 26682
rect 30087 26630 44134 26682
rect 44186 26630 44238 26682
rect 44290 26630 44342 26682
rect 44394 26630 58441 26682
rect 58493 26630 58545 26682
rect 58597 26630 58649 26682
rect 58701 26630 58731 26682
rect 1344 26596 58731 26630
rect 2494 26514 2546 26526
rect 2494 26450 2546 26462
rect 3054 26514 3106 26526
rect 3054 26450 3106 26462
rect 6414 26514 6466 26526
rect 6414 26450 6466 26462
rect 7198 26514 7250 26526
rect 7198 26450 7250 26462
rect 8878 26514 8930 26526
rect 8878 26450 8930 26462
rect 10446 26514 10498 26526
rect 10446 26450 10498 26462
rect 24334 26514 24386 26526
rect 30718 26514 30770 26526
rect 25218 26462 25230 26514
rect 25282 26462 25294 26514
rect 24334 26450 24386 26462
rect 30718 26450 30770 26462
rect 33406 26514 33458 26526
rect 33406 26450 33458 26462
rect 33518 26514 33570 26526
rect 33518 26450 33570 26462
rect 34526 26514 34578 26526
rect 34526 26450 34578 26462
rect 35758 26514 35810 26526
rect 35758 26450 35810 26462
rect 36206 26514 36258 26526
rect 36206 26450 36258 26462
rect 36318 26514 36370 26526
rect 40798 26514 40850 26526
rect 36754 26462 36766 26514
rect 36818 26462 36830 26514
rect 39666 26462 39678 26514
rect 39730 26462 39742 26514
rect 36318 26450 36370 26462
rect 40798 26450 40850 26462
rect 45390 26514 45442 26526
rect 47506 26462 47518 26514
rect 47570 26462 47582 26514
rect 45390 26450 45442 26462
rect 2046 26402 2098 26414
rect 2046 26338 2098 26350
rect 3502 26402 3554 26414
rect 3502 26338 3554 26350
rect 4062 26402 4114 26414
rect 4062 26338 4114 26350
rect 4622 26402 4674 26414
rect 8990 26402 9042 26414
rect 8306 26350 8318 26402
rect 8370 26350 8382 26402
rect 4622 26338 4674 26350
rect 8990 26338 9042 26350
rect 10222 26402 10274 26414
rect 20526 26402 20578 26414
rect 11442 26350 11454 26402
rect 11506 26350 11518 26402
rect 10222 26338 10274 26350
rect 20526 26338 20578 26350
rect 20638 26402 20690 26414
rect 20638 26338 20690 26350
rect 23550 26402 23602 26414
rect 23550 26338 23602 26350
rect 24558 26402 24610 26414
rect 33182 26402 33234 26414
rect 28466 26350 28478 26402
rect 28530 26350 28542 26402
rect 30930 26350 30942 26402
rect 30994 26350 31006 26402
rect 24558 26338 24610 26350
rect 33182 26338 33234 26350
rect 33742 26402 33794 26414
rect 33742 26338 33794 26350
rect 34302 26402 34354 26414
rect 34302 26338 34354 26350
rect 34862 26402 34914 26414
rect 34862 26338 34914 26350
rect 35310 26402 35362 26414
rect 35310 26338 35362 26350
rect 38334 26402 38386 26414
rect 38334 26338 38386 26350
rect 40126 26402 40178 26414
rect 40126 26338 40178 26350
rect 41022 26402 41074 26414
rect 41022 26338 41074 26350
rect 44494 26402 44546 26414
rect 44494 26338 44546 26350
rect 46622 26402 46674 26414
rect 54798 26402 54850 26414
rect 49074 26350 49086 26402
rect 49138 26350 49150 26402
rect 51650 26350 51662 26402
rect 51714 26350 51726 26402
rect 52546 26350 52558 26402
rect 52610 26350 52622 26402
rect 46622 26338 46674 26350
rect 54798 26338 54850 26350
rect 55918 26402 55970 26414
rect 55918 26338 55970 26350
rect 2830 26290 2882 26302
rect 1810 26238 1822 26290
rect 1874 26238 1886 26290
rect 2830 26226 2882 26238
rect 3278 26290 3330 26302
rect 3278 26226 3330 26238
rect 3838 26290 3890 26302
rect 3838 26226 3890 26238
rect 4174 26290 4226 26302
rect 4174 26226 4226 26238
rect 4510 26290 4562 26302
rect 4510 26226 4562 26238
rect 6078 26290 6130 26302
rect 6078 26226 6130 26238
rect 6526 26290 6578 26302
rect 6526 26226 6578 26238
rect 6750 26290 6802 26302
rect 6750 26226 6802 26238
rect 7534 26290 7586 26302
rect 8654 26290 8706 26302
rect 7970 26238 7982 26290
rect 8034 26238 8046 26290
rect 7534 26226 7586 26238
rect 8654 26226 8706 26238
rect 10110 26290 10162 26302
rect 20302 26290 20354 26302
rect 10770 26238 10782 26290
rect 10834 26238 10846 26290
rect 15026 26238 15038 26290
rect 15090 26238 15102 26290
rect 16370 26238 16382 26290
rect 16434 26238 16446 26290
rect 17938 26238 17950 26290
rect 18002 26238 18014 26290
rect 18946 26238 18958 26290
rect 19010 26238 19022 26290
rect 10110 26226 10162 26238
rect 20302 26226 20354 26238
rect 21310 26290 21362 26302
rect 21310 26226 21362 26238
rect 21534 26290 21586 26302
rect 21534 26226 21586 26238
rect 21982 26290 22034 26302
rect 21982 26226 22034 26238
rect 22654 26290 22706 26302
rect 22654 26226 22706 26238
rect 22878 26290 22930 26302
rect 22878 26226 22930 26238
rect 23774 26290 23826 26302
rect 23774 26226 23826 26238
rect 24670 26290 24722 26302
rect 24670 26226 24722 26238
rect 25566 26290 25618 26302
rect 33070 26290 33122 26302
rect 29362 26238 29374 26290
rect 29426 26238 29438 26290
rect 31042 26238 31054 26290
rect 31106 26238 31118 26290
rect 31602 26238 31614 26290
rect 31666 26238 31678 26290
rect 32386 26238 32398 26290
rect 32450 26238 32462 26290
rect 25566 26226 25618 26238
rect 33070 26226 33122 26238
rect 33854 26290 33906 26302
rect 33854 26226 33906 26238
rect 34190 26290 34242 26302
rect 34190 26226 34242 26238
rect 37102 26290 37154 26302
rect 37102 26226 37154 26238
rect 38222 26290 38274 26302
rect 38222 26226 38274 26238
rect 38558 26290 38610 26302
rect 38558 26226 38610 26238
rect 40350 26290 40402 26302
rect 40350 26226 40402 26238
rect 41134 26290 41186 26302
rect 41134 26226 41186 26238
rect 44606 26290 44658 26302
rect 46510 26290 46562 26302
rect 46050 26238 46062 26290
rect 46114 26238 46126 26290
rect 50418 26238 50430 26290
rect 50482 26238 50494 26290
rect 53218 26238 53230 26290
rect 53282 26238 53294 26290
rect 53442 26238 53454 26290
rect 53506 26238 53518 26290
rect 55122 26238 55134 26290
rect 55186 26238 55198 26290
rect 57138 26238 57150 26290
rect 57202 26238 57214 26290
rect 44606 26226 44658 26238
rect 46510 26226 46562 26238
rect 9774 26178 9826 26190
rect 21422 26178 21474 26190
rect 13570 26126 13582 26178
rect 13634 26126 13646 26178
rect 16482 26126 16494 26178
rect 16546 26126 16558 26178
rect 17714 26126 17726 26178
rect 17778 26126 17790 26178
rect 9774 26114 9826 26126
rect 21422 26114 21474 26126
rect 22318 26178 22370 26190
rect 22318 26114 22370 26126
rect 27582 26178 27634 26190
rect 37998 26178 38050 26190
rect 28466 26126 28478 26178
rect 28530 26126 28542 26178
rect 27582 26114 27634 26126
rect 37998 26114 38050 26126
rect 39118 26178 39170 26190
rect 46958 26178 47010 26190
rect 40002 26126 40014 26178
rect 40066 26126 40078 26178
rect 39118 26114 39170 26126
rect 46958 26114 47010 26126
rect 47966 26178 48018 26190
rect 52110 26178 52162 26190
rect 48962 26126 48974 26178
rect 49026 26126 49038 26178
rect 47966 26114 48018 26126
rect 52110 26114 52162 26126
rect 54910 26178 54962 26190
rect 54910 26114 54962 26126
rect 55694 26178 55746 26190
rect 55694 26114 55746 26126
rect 55806 26178 55858 26190
rect 57598 26178 57650 26190
rect 56690 26126 56702 26178
rect 56754 26126 56766 26178
rect 55806 26114 55858 26126
rect 57598 26114 57650 26126
rect 58046 26178 58098 26190
rect 58046 26114 58098 26126
rect 4622 26066 4674 26078
rect 24110 26066 24162 26078
rect 14802 26014 14814 26066
rect 14866 26014 14878 26066
rect 19170 26014 19182 26066
rect 19234 26014 19246 26066
rect 23202 26014 23214 26066
rect 23266 26014 23278 26066
rect 4622 26002 4674 26014
rect 24110 26002 24162 26014
rect 36430 26066 36482 26078
rect 36430 26002 36482 26014
rect 39342 26066 39394 26078
rect 39342 26002 39394 26014
rect 44494 26066 44546 26078
rect 44494 26002 44546 26014
rect 47182 26066 47234 26078
rect 47182 26002 47234 26014
rect 1344 25898 58576 25932
rect 1344 25846 8367 25898
rect 8419 25846 8471 25898
rect 8523 25846 8575 25898
rect 8627 25846 22674 25898
rect 22726 25846 22778 25898
rect 22830 25846 22882 25898
rect 22934 25846 36981 25898
rect 37033 25846 37085 25898
rect 37137 25846 37189 25898
rect 37241 25846 51288 25898
rect 51340 25846 51392 25898
rect 51444 25846 51496 25898
rect 51548 25846 58576 25898
rect 1344 25812 58576 25846
rect 8542 25730 8594 25742
rect 8542 25666 8594 25678
rect 32062 25730 32114 25742
rect 32062 25666 32114 25678
rect 33966 25730 34018 25742
rect 33966 25666 34018 25678
rect 36990 25730 37042 25742
rect 36990 25666 37042 25678
rect 46958 25730 47010 25742
rect 46958 25666 47010 25678
rect 54014 25730 54066 25742
rect 54014 25666 54066 25678
rect 8206 25618 8258 25630
rect 4834 25566 4846 25618
rect 4898 25566 4910 25618
rect 8206 25554 8258 25566
rect 12462 25618 12514 25630
rect 12462 25554 12514 25566
rect 13694 25618 13746 25630
rect 13694 25554 13746 25566
rect 16046 25618 16098 25630
rect 16046 25554 16098 25566
rect 17166 25618 17218 25630
rect 17166 25554 17218 25566
rect 18734 25618 18786 25630
rect 31614 25618 31666 25630
rect 19618 25566 19630 25618
rect 19682 25566 19694 25618
rect 23874 25566 23886 25618
rect 23938 25566 23950 25618
rect 29586 25566 29598 25618
rect 29650 25566 29662 25618
rect 18734 25554 18786 25566
rect 31614 25554 31666 25566
rect 31950 25618 32002 25630
rect 31950 25554 32002 25566
rect 34974 25618 35026 25630
rect 45166 25618 45218 25630
rect 47070 25618 47122 25630
rect 39442 25566 39454 25618
rect 39506 25566 39518 25618
rect 41682 25566 41694 25618
rect 41746 25566 41758 25618
rect 42466 25566 42478 25618
rect 42530 25566 42542 25618
rect 46162 25566 46174 25618
rect 46226 25566 46238 25618
rect 34974 25554 35026 25566
rect 45166 25554 45218 25566
rect 47070 25554 47122 25566
rect 47742 25618 47794 25630
rect 47742 25554 47794 25566
rect 49534 25618 49586 25630
rect 49534 25554 49586 25566
rect 51662 25618 51714 25630
rect 51662 25554 51714 25566
rect 53230 25618 53282 25630
rect 56018 25566 56030 25618
rect 56082 25566 56094 25618
rect 56466 25566 56478 25618
rect 56530 25566 56542 25618
rect 53230 25554 53282 25566
rect 11454 25506 11506 25518
rect 2034 25454 2046 25506
rect 2098 25454 2110 25506
rect 11454 25442 11506 25454
rect 12014 25506 12066 25518
rect 12014 25442 12066 25454
rect 14366 25506 14418 25518
rect 16382 25506 16434 25518
rect 21758 25506 21810 25518
rect 27918 25506 27970 25518
rect 30718 25506 30770 25518
rect 38222 25506 38274 25518
rect 15586 25454 15598 25506
rect 15650 25454 15662 25506
rect 15810 25454 15822 25506
rect 15874 25454 15886 25506
rect 19394 25454 19406 25506
rect 19458 25454 19470 25506
rect 26450 25454 26462 25506
rect 26514 25454 26526 25506
rect 29138 25454 29150 25506
rect 29202 25454 29214 25506
rect 30034 25454 30046 25506
rect 30098 25454 30110 25506
rect 31154 25454 31166 25506
rect 31218 25454 31230 25506
rect 33506 25454 33518 25506
rect 33570 25454 33582 25506
rect 34178 25454 34190 25506
rect 34242 25454 34254 25506
rect 34850 25454 34862 25506
rect 34914 25454 34926 25506
rect 35634 25454 35646 25506
rect 35698 25454 35710 25506
rect 14366 25442 14418 25454
rect 16382 25442 16434 25454
rect 21758 25442 21810 25454
rect 27918 25442 27970 25454
rect 30718 25442 30770 25454
rect 38222 25442 38274 25454
rect 38558 25506 38610 25518
rect 43150 25506 43202 25518
rect 39666 25454 39678 25506
rect 39730 25454 39742 25506
rect 41122 25454 41134 25506
rect 41186 25454 41198 25506
rect 42578 25454 42590 25506
rect 42642 25454 42654 25506
rect 38558 25442 38610 25454
rect 43150 25442 43202 25454
rect 43934 25506 43986 25518
rect 43934 25442 43986 25454
rect 44718 25506 44770 25518
rect 44718 25442 44770 25454
rect 45390 25506 45442 25518
rect 45390 25442 45442 25454
rect 48638 25506 48690 25518
rect 51550 25506 51602 25518
rect 49074 25454 49086 25506
rect 49138 25454 49150 25506
rect 51202 25454 51214 25506
rect 51266 25454 51278 25506
rect 53666 25454 53678 25506
rect 53730 25454 53742 25506
rect 55122 25454 55134 25506
rect 55186 25454 55198 25506
rect 55906 25454 55918 25506
rect 55970 25454 55982 25506
rect 57250 25454 57262 25506
rect 57314 25454 57326 25506
rect 57698 25454 57710 25506
rect 57762 25454 57774 25506
rect 48638 25442 48690 25454
rect 51550 25442 51602 25454
rect 10334 25394 10386 25406
rect 2706 25342 2718 25394
rect 2770 25342 2782 25394
rect 7634 25342 7646 25394
rect 7698 25342 7710 25394
rect 7970 25342 7982 25394
rect 8034 25342 8046 25394
rect 10334 25330 10386 25342
rect 10670 25394 10722 25406
rect 10670 25330 10722 25342
rect 10894 25394 10946 25406
rect 10894 25330 10946 25342
rect 11230 25394 11282 25406
rect 11230 25330 11282 25342
rect 11678 25394 11730 25406
rect 11678 25330 11730 25342
rect 11902 25394 11954 25406
rect 11902 25330 11954 25342
rect 21646 25394 21698 25406
rect 21646 25330 21698 25342
rect 27806 25394 27858 25406
rect 27806 25330 27858 25342
rect 28030 25394 28082 25406
rect 37326 25394 37378 25406
rect 29810 25342 29822 25394
rect 29874 25342 29886 25394
rect 32946 25342 32958 25394
rect 33010 25342 33022 25394
rect 33170 25342 33182 25394
rect 33234 25342 33246 25394
rect 35858 25342 35870 25394
rect 35922 25342 35934 25394
rect 28030 25330 28082 25342
rect 37326 25330 37378 25342
rect 37774 25394 37826 25406
rect 37774 25330 37826 25342
rect 37886 25394 37938 25406
rect 37886 25330 37938 25342
rect 38334 25394 38386 25406
rect 38334 25330 38386 25342
rect 38782 25394 38834 25406
rect 38782 25330 38834 25342
rect 44270 25394 44322 25406
rect 50094 25394 50146 25406
rect 46498 25342 46510 25394
rect 46562 25342 46574 25394
rect 44270 25330 44322 25342
rect 50094 25330 50146 25342
rect 54238 25394 54290 25406
rect 56130 25342 56142 25394
rect 56194 25342 56206 25394
rect 54238 25330 54290 25342
rect 9998 25282 10050 25294
rect 9998 25218 10050 25230
rect 10446 25282 10498 25294
rect 10446 25218 10498 25230
rect 11118 25282 11170 25294
rect 20190 25282 20242 25294
rect 14018 25230 14030 25282
rect 14082 25230 14094 25282
rect 16706 25230 16718 25282
rect 16770 25230 16782 25282
rect 11118 25218 11170 25230
rect 20190 25218 20242 25230
rect 21422 25282 21474 25294
rect 21422 25218 21474 25230
rect 28702 25282 28754 25294
rect 36430 25282 36482 25294
rect 32722 25230 32734 25282
rect 32786 25230 32798 25282
rect 28702 25218 28754 25230
rect 36430 25218 36482 25230
rect 37102 25282 37154 25294
rect 37102 25218 37154 25230
rect 37550 25282 37602 25294
rect 37550 25218 37602 25230
rect 38894 25282 38946 25294
rect 38894 25218 38946 25230
rect 39118 25282 39170 25294
rect 39118 25218 39170 25230
rect 44158 25282 44210 25294
rect 44158 25218 44210 25230
rect 47182 25282 47234 25294
rect 47182 25218 47234 25230
rect 48190 25282 48242 25294
rect 48190 25218 48242 25230
rect 50206 25282 50258 25294
rect 50206 25218 50258 25230
rect 50430 25282 50482 25294
rect 50430 25218 50482 25230
rect 52110 25282 52162 25294
rect 52110 25218 52162 25230
rect 53118 25282 53170 25294
rect 53118 25218 53170 25230
rect 53342 25282 53394 25294
rect 53342 25218 53394 25230
rect 54126 25282 54178 25294
rect 54126 25218 54178 25230
rect 1344 25114 58731 25148
rect 1344 25062 15520 25114
rect 15572 25062 15624 25114
rect 15676 25062 15728 25114
rect 15780 25062 29827 25114
rect 29879 25062 29931 25114
rect 29983 25062 30035 25114
rect 30087 25062 44134 25114
rect 44186 25062 44238 25114
rect 44290 25062 44342 25114
rect 44394 25062 58441 25114
rect 58493 25062 58545 25114
rect 58597 25062 58649 25114
rect 58701 25062 58731 25114
rect 1344 25028 58731 25062
rect 2158 24946 2210 24958
rect 2158 24882 2210 24894
rect 3166 24946 3218 24958
rect 3166 24882 3218 24894
rect 4846 24946 4898 24958
rect 23662 24946 23714 24958
rect 22866 24894 22878 24946
rect 22930 24894 22942 24946
rect 4846 24882 4898 24894
rect 23662 24882 23714 24894
rect 23886 24946 23938 24958
rect 23886 24882 23938 24894
rect 24110 24946 24162 24958
rect 24110 24882 24162 24894
rect 27134 24946 27186 24958
rect 27134 24882 27186 24894
rect 32286 24946 32338 24958
rect 32286 24882 32338 24894
rect 42254 24946 42306 24958
rect 42254 24882 42306 24894
rect 42590 24946 42642 24958
rect 42590 24882 42642 24894
rect 3390 24834 3442 24846
rect 3390 24770 3442 24782
rect 4062 24834 4114 24846
rect 4062 24770 4114 24782
rect 4622 24834 4674 24846
rect 17502 24834 17554 24846
rect 25230 24834 25282 24846
rect 11106 24782 11118 24834
rect 11170 24782 11182 24834
rect 21410 24782 21422 24834
rect 21474 24782 21486 24834
rect 22978 24782 22990 24834
rect 23042 24782 23054 24834
rect 4622 24770 4674 24782
rect 17502 24770 17554 24782
rect 25230 24770 25282 24782
rect 29150 24834 29202 24846
rect 29150 24770 29202 24782
rect 30494 24834 30546 24846
rect 30494 24770 30546 24782
rect 34078 24834 34130 24846
rect 34078 24770 34130 24782
rect 36766 24834 36818 24846
rect 36766 24770 36818 24782
rect 36878 24834 36930 24846
rect 36878 24770 36930 24782
rect 38110 24834 38162 24846
rect 38110 24770 38162 24782
rect 38670 24834 38722 24846
rect 41918 24834 41970 24846
rect 39218 24782 39230 24834
rect 39282 24782 39294 24834
rect 38670 24770 38722 24782
rect 41918 24770 41970 24782
rect 42814 24834 42866 24846
rect 42814 24770 42866 24782
rect 44046 24834 44098 24846
rect 44046 24770 44098 24782
rect 45502 24834 45554 24846
rect 45502 24770 45554 24782
rect 45838 24834 45890 24846
rect 45838 24770 45890 24782
rect 50542 24834 50594 24846
rect 55358 24834 55410 24846
rect 51426 24782 51438 24834
rect 51490 24782 51502 24834
rect 53442 24782 53454 24834
rect 53506 24782 53518 24834
rect 50542 24770 50594 24782
rect 55358 24770 55410 24782
rect 56590 24834 56642 24846
rect 56590 24770 56642 24782
rect 2494 24722 2546 24734
rect 2494 24658 2546 24670
rect 3054 24722 3106 24734
rect 3054 24658 3106 24670
rect 3502 24722 3554 24734
rect 3502 24658 3554 24670
rect 3950 24722 4002 24734
rect 3950 24658 4002 24670
rect 4510 24722 4562 24734
rect 15934 24722 15986 24734
rect 23774 24722 23826 24734
rect 5730 24670 5742 24722
rect 5794 24670 5806 24722
rect 10322 24670 10334 24722
rect 10386 24670 10398 24722
rect 15474 24670 15486 24722
rect 15538 24670 15550 24722
rect 18274 24670 18286 24722
rect 18338 24670 18350 24722
rect 19618 24670 19630 24722
rect 19682 24670 19694 24722
rect 21634 24670 21646 24722
rect 21698 24670 21710 24722
rect 4510 24658 4562 24670
rect 15934 24658 15986 24670
rect 23774 24658 23826 24670
rect 25342 24722 25394 24734
rect 29262 24722 29314 24734
rect 31726 24722 31778 24734
rect 25666 24670 25678 24722
rect 25730 24670 25742 24722
rect 27570 24670 27582 24722
rect 27634 24670 27646 24722
rect 29810 24670 29822 24722
rect 29874 24670 29886 24722
rect 25342 24658 25394 24670
rect 29262 24658 29314 24670
rect 31726 24658 31778 24670
rect 32174 24722 32226 24734
rect 32174 24658 32226 24670
rect 32398 24722 32450 24734
rect 32398 24658 32450 24670
rect 33182 24722 33234 24734
rect 37102 24722 37154 24734
rect 33394 24670 33406 24722
rect 33458 24670 33470 24722
rect 34850 24670 34862 24722
rect 34914 24670 34926 24722
rect 35970 24670 35982 24722
rect 36034 24670 36046 24722
rect 33182 24658 33234 24670
rect 37102 24658 37154 24670
rect 38446 24722 38498 24734
rect 42142 24722 42194 24734
rect 39106 24670 39118 24722
rect 39170 24670 39182 24722
rect 40002 24670 40014 24722
rect 40066 24670 40078 24722
rect 38446 24658 38498 24670
rect 42142 24658 42194 24670
rect 42366 24722 42418 24734
rect 42366 24658 42418 24670
rect 42926 24722 42978 24734
rect 42926 24658 42978 24670
rect 43934 24722 43986 24734
rect 43934 24658 43986 24670
rect 44270 24722 44322 24734
rect 44270 24658 44322 24670
rect 44606 24722 44658 24734
rect 47854 24722 47906 24734
rect 50430 24722 50482 24734
rect 45042 24670 45054 24722
rect 45106 24670 45118 24722
rect 48626 24670 48638 24722
rect 48690 24670 48702 24722
rect 49410 24670 49422 24722
rect 49474 24670 49486 24722
rect 44606 24658 44658 24670
rect 47854 24658 47906 24670
rect 50430 24658 50482 24670
rect 50766 24722 50818 24734
rect 56814 24722 56866 24734
rect 51314 24670 51326 24722
rect 51378 24670 51390 24722
rect 51538 24670 51550 24722
rect 51602 24670 51614 24722
rect 52210 24670 52222 24722
rect 52274 24670 52286 24722
rect 54002 24670 54014 24722
rect 54066 24670 54078 24722
rect 54674 24670 54686 24722
rect 54738 24670 54750 24722
rect 56018 24670 56030 24722
rect 56082 24670 56094 24722
rect 57026 24670 57038 24722
rect 57090 24670 57102 24722
rect 50766 24658 50818 24670
rect 56814 24658 56866 24670
rect 15038 24610 15090 24622
rect 31502 24610 31554 24622
rect 6514 24558 6526 24610
rect 6578 24558 6590 24610
rect 8642 24558 8654 24610
rect 8706 24558 8718 24610
rect 13346 24558 13358 24610
rect 13410 24558 13422 24610
rect 19730 24558 19742 24610
rect 19794 24558 19806 24610
rect 27906 24558 27918 24610
rect 27970 24558 27982 24610
rect 30930 24558 30942 24610
rect 30994 24558 31006 24610
rect 15038 24546 15090 24558
rect 31502 24546 31554 24558
rect 34414 24610 34466 24622
rect 36318 24610 36370 24622
rect 36194 24558 36206 24610
rect 36258 24558 36270 24610
rect 34414 24546 34466 24558
rect 36318 24546 36370 24558
rect 37998 24610 38050 24622
rect 46398 24610 46450 24622
rect 38770 24558 38782 24610
rect 38834 24558 38846 24610
rect 39554 24558 39566 24610
rect 39618 24558 39630 24610
rect 37998 24546 38050 24558
rect 46398 24546 46450 24558
rect 47406 24610 47458 24622
rect 47406 24546 47458 24558
rect 47630 24610 47682 24622
rect 47630 24546 47682 24558
rect 48190 24610 48242 24622
rect 55806 24610 55858 24622
rect 48850 24558 48862 24610
rect 48914 24558 48926 24610
rect 49298 24558 49310 24610
rect 49362 24558 49374 24610
rect 48190 24546 48242 24558
rect 55806 24546 55858 24558
rect 58158 24610 58210 24622
rect 58158 24546 58210 24558
rect 4062 24498 4114 24510
rect 46062 24498 46114 24510
rect 28018 24446 28030 24498
rect 28082 24446 28094 24498
rect 4062 24434 4114 24446
rect 46062 24434 46114 24446
rect 55694 24498 55746 24510
rect 55694 24434 55746 24446
rect 1344 24330 58576 24364
rect 1344 24278 8367 24330
rect 8419 24278 8471 24330
rect 8523 24278 8575 24330
rect 8627 24278 22674 24330
rect 22726 24278 22778 24330
rect 22830 24278 22882 24330
rect 22934 24278 36981 24330
rect 37033 24278 37085 24330
rect 37137 24278 37189 24330
rect 37241 24278 51288 24330
rect 51340 24278 51392 24330
rect 51444 24278 51496 24330
rect 51548 24278 58576 24330
rect 1344 24244 58576 24278
rect 7534 24162 7586 24174
rect 7534 24098 7586 24110
rect 18510 24162 18562 24174
rect 42030 24162 42082 24174
rect 55246 24162 55298 24174
rect 32498 24110 32510 24162
rect 32562 24110 32574 24162
rect 47842 24110 47854 24162
rect 47906 24110 47918 24162
rect 51986 24110 51998 24162
rect 52050 24110 52062 24162
rect 18510 24098 18562 24110
rect 42030 24098 42082 24110
rect 55246 24098 55298 24110
rect 55582 24162 55634 24174
rect 55582 24098 55634 24110
rect 6638 24050 6690 24062
rect 6638 23986 6690 23998
rect 9438 24050 9490 24062
rect 9438 23986 9490 23998
rect 10222 24050 10274 24062
rect 17726 24050 17778 24062
rect 16370 23998 16382 24050
rect 16434 23998 16446 24050
rect 10222 23986 10274 23998
rect 17726 23986 17778 23998
rect 17950 24050 18002 24062
rect 17950 23986 18002 23998
rect 18286 24050 18338 24062
rect 18286 23986 18338 23998
rect 19630 24050 19682 24062
rect 30158 24050 30210 24062
rect 37550 24050 37602 24062
rect 40574 24050 40626 24062
rect 21410 23998 21422 24050
rect 21474 23998 21486 24050
rect 27010 23998 27022 24050
rect 27074 23998 27086 24050
rect 33618 23998 33630 24050
rect 33682 23998 33694 24050
rect 35522 23998 35534 24050
rect 35586 23998 35598 24050
rect 38434 23998 38446 24050
rect 38498 23998 38510 24050
rect 19630 23986 19682 23998
rect 30158 23986 30210 23998
rect 37550 23986 37602 23998
rect 40574 23986 40626 23998
rect 45278 24050 45330 24062
rect 45278 23986 45330 23998
rect 46510 24050 46562 24062
rect 53342 24050 53394 24062
rect 48514 23998 48526 24050
rect 48578 23998 48590 24050
rect 51314 23998 51326 24050
rect 51378 23998 51390 24050
rect 46510 23986 46562 23998
rect 53342 23986 53394 23998
rect 2046 23938 2098 23950
rect 2046 23874 2098 23886
rect 2382 23938 2434 23950
rect 2382 23874 2434 23886
rect 3054 23938 3106 23950
rect 3054 23874 3106 23886
rect 4062 23938 4114 23950
rect 4062 23874 4114 23886
rect 6414 23938 6466 23950
rect 6414 23874 6466 23886
rect 6862 23938 6914 23950
rect 6862 23874 6914 23886
rect 7646 23938 7698 23950
rect 7646 23874 7698 23886
rect 8206 23938 8258 23950
rect 8206 23874 8258 23886
rect 10894 23938 10946 23950
rect 19518 23938 19570 23950
rect 13458 23886 13470 23938
rect 13522 23886 13534 23938
rect 10894 23874 10946 23886
rect 19518 23874 19570 23886
rect 24334 23938 24386 23950
rect 24334 23874 24386 23886
rect 24670 23938 24722 23950
rect 24670 23874 24722 23886
rect 26126 23938 26178 23950
rect 27806 23938 27858 23950
rect 26786 23886 26798 23938
rect 26850 23886 26862 23938
rect 26126 23874 26178 23886
rect 27806 23874 27858 23886
rect 28478 23938 28530 23950
rect 28478 23874 28530 23886
rect 28590 23938 28642 23950
rect 28590 23874 28642 23886
rect 29262 23938 29314 23950
rect 32398 23938 32450 23950
rect 41246 23938 41298 23950
rect 29474 23886 29486 23938
rect 29538 23886 29550 23938
rect 30706 23886 30718 23938
rect 30770 23886 30782 23938
rect 32050 23886 32062 23938
rect 32114 23886 32126 23938
rect 32946 23886 32958 23938
rect 33010 23886 33022 23938
rect 34066 23886 34078 23938
rect 34130 23886 34142 23938
rect 35858 23886 35870 23938
rect 35922 23886 35934 23938
rect 37090 23886 37102 23938
rect 37154 23886 37166 23938
rect 39890 23886 39902 23938
rect 39954 23886 39966 23938
rect 29262 23874 29314 23886
rect 32398 23874 32450 23886
rect 41246 23874 41298 23886
rect 41694 23938 41746 23950
rect 46062 23938 46114 23950
rect 49086 23938 49138 23950
rect 42690 23886 42702 23938
rect 42754 23886 42766 23938
rect 48178 23886 48190 23938
rect 48242 23886 48254 23938
rect 41694 23874 41746 23886
rect 46062 23874 46114 23886
rect 49086 23874 49138 23886
rect 49422 23938 49474 23950
rect 49422 23874 49474 23886
rect 49758 23938 49810 23950
rect 49758 23874 49810 23886
rect 50430 23938 50482 23950
rect 52558 23938 52610 23950
rect 51650 23886 51662 23938
rect 51714 23886 51726 23938
rect 56802 23886 56814 23938
rect 56866 23886 56878 23938
rect 57586 23886 57598 23938
rect 57650 23886 57662 23938
rect 50430 23874 50482 23886
rect 52558 23874 52610 23886
rect 2606 23826 2658 23838
rect 2606 23762 2658 23774
rect 3278 23826 3330 23838
rect 3278 23762 3330 23774
rect 3390 23826 3442 23838
rect 3390 23762 3442 23774
rect 4398 23826 4450 23838
rect 4398 23762 4450 23774
rect 7086 23826 7138 23838
rect 7086 23762 7138 23774
rect 7870 23826 7922 23838
rect 7870 23762 7922 23774
rect 8094 23826 8146 23838
rect 11342 23826 11394 23838
rect 10546 23774 10558 23826
rect 10610 23774 10622 23826
rect 8094 23762 8146 23774
rect 11342 23762 11394 23774
rect 11454 23826 11506 23838
rect 11454 23762 11506 23774
rect 11902 23826 11954 23838
rect 11902 23762 11954 23774
rect 12014 23826 12066 23838
rect 12014 23762 12066 23774
rect 12574 23826 12626 23838
rect 19182 23826 19234 23838
rect 14242 23774 14254 23826
rect 14306 23774 14318 23826
rect 18834 23774 18846 23826
rect 18898 23774 18910 23826
rect 12574 23762 12626 23774
rect 19182 23762 19234 23774
rect 19742 23826 19794 23838
rect 25342 23826 25394 23838
rect 35198 23826 35250 23838
rect 40910 23826 40962 23838
rect 21746 23774 21758 23826
rect 21810 23774 21822 23826
rect 23314 23774 23326 23826
rect 23378 23774 23390 23826
rect 30482 23774 30494 23826
rect 30546 23774 30558 23826
rect 33058 23774 33070 23826
rect 33122 23774 33134 23826
rect 38994 23774 39006 23826
rect 39058 23774 39070 23826
rect 19742 23762 19794 23774
rect 25342 23762 25394 23774
rect 35198 23762 35250 23774
rect 40910 23762 40962 23774
rect 41470 23826 41522 23838
rect 41470 23762 41522 23774
rect 45726 23826 45778 23838
rect 45726 23762 45778 23774
rect 45838 23826 45890 23838
rect 45838 23762 45890 23774
rect 52894 23826 52946 23838
rect 58158 23826 58210 23838
rect 56242 23774 56254 23826
rect 56306 23774 56318 23826
rect 52894 23762 52946 23774
rect 58158 23762 58210 23774
rect 2158 23714 2210 23726
rect 2158 23650 2210 23662
rect 2718 23714 2770 23726
rect 2718 23650 2770 23662
rect 2942 23714 2994 23726
rect 2942 23650 2994 23662
rect 3726 23714 3778 23726
rect 3726 23650 3778 23662
rect 3950 23714 4002 23726
rect 3950 23650 4002 23662
rect 4510 23714 4562 23726
rect 4510 23650 4562 23662
rect 4734 23714 4786 23726
rect 4734 23650 4786 23662
rect 7534 23714 7586 23726
rect 7534 23650 7586 23662
rect 11118 23714 11170 23726
rect 11118 23650 11170 23662
rect 12238 23714 12290 23726
rect 24558 23714 24610 23726
rect 17378 23662 17390 23714
rect 17442 23662 17454 23714
rect 23202 23662 23214 23714
rect 23266 23662 23278 23714
rect 12238 23650 12290 23662
rect 24558 23650 24610 23662
rect 25230 23714 25282 23726
rect 25230 23650 25282 23662
rect 25790 23714 25842 23726
rect 25790 23650 25842 23662
rect 27582 23714 27634 23726
rect 27582 23650 27634 23662
rect 27694 23714 27746 23726
rect 27694 23650 27746 23662
rect 28030 23714 28082 23726
rect 28030 23650 28082 23662
rect 34638 23714 34690 23726
rect 34638 23650 34690 23662
rect 41022 23714 41074 23726
rect 43598 23714 43650 23726
rect 42914 23662 42926 23714
rect 42978 23662 42990 23714
rect 41022 23650 41074 23662
rect 43598 23650 43650 23662
rect 44942 23714 44994 23726
rect 44942 23650 44994 23662
rect 45166 23714 45218 23726
rect 45166 23650 45218 23662
rect 45390 23714 45442 23726
rect 47182 23714 47234 23726
rect 46834 23662 46846 23714
rect 46898 23662 46910 23714
rect 45390 23650 45442 23662
rect 47182 23650 47234 23662
rect 49310 23714 49362 23726
rect 49310 23650 49362 23662
rect 49870 23714 49922 23726
rect 49870 23650 49922 23662
rect 50094 23714 50146 23726
rect 50094 23650 50146 23662
rect 50542 23714 50594 23726
rect 50542 23650 50594 23662
rect 50766 23714 50818 23726
rect 50766 23650 50818 23662
rect 52782 23714 52834 23726
rect 52782 23650 52834 23662
rect 55358 23714 55410 23726
rect 55358 23650 55410 23662
rect 1344 23546 58731 23580
rect 1344 23494 15520 23546
rect 15572 23494 15624 23546
rect 15676 23494 15728 23546
rect 15780 23494 29827 23546
rect 29879 23494 29931 23546
rect 29983 23494 30035 23546
rect 30087 23494 44134 23546
rect 44186 23494 44238 23546
rect 44290 23494 44342 23546
rect 44394 23494 58441 23546
rect 58493 23494 58545 23546
rect 58597 23494 58649 23546
rect 58701 23494 58731 23546
rect 1344 23460 58731 23494
rect 14030 23378 14082 23390
rect 8418 23326 8430 23378
rect 8482 23326 8494 23378
rect 14030 23314 14082 23326
rect 15150 23378 15202 23390
rect 15150 23314 15202 23326
rect 15710 23378 15762 23390
rect 15710 23314 15762 23326
rect 16382 23378 16434 23390
rect 16382 23314 16434 23326
rect 20638 23378 20690 23390
rect 31390 23378 31442 23390
rect 28914 23326 28926 23378
rect 28978 23326 28990 23378
rect 20638 23314 20690 23326
rect 31390 23314 31442 23326
rect 32174 23378 32226 23390
rect 32174 23314 32226 23326
rect 32398 23378 32450 23390
rect 32398 23314 32450 23326
rect 33294 23378 33346 23390
rect 33294 23314 33346 23326
rect 33966 23378 34018 23390
rect 33966 23314 34018 23326
rect 35534 23378 35586 23390
rect 35534 23314 35586 23326
rect 35870 23378 35922 23390
rect 35870 23314 35922 23326
rect 37550 23378 37602 23390
rect 37550 23314 37602 23326
rect 42814 23378 42866 23390
rect 47630 23378 47682 23390
rect 43474 23326 43486 23378
rect 43538 23326 43550 23378
rect 44706 23326 44718 23378
rect 44770 23326 44782 23378
rect 42814 23314 42866 23326
rect 47630 23314 47682 23326
rect 47966 23378 48018 23390
rect 47966 23314 48018 23326
rect 50206 23378 50258 23390
rect 50978 23326 50990 23378
rect 51042 23326 51054 23378
rect 50206 23314 50258 23326
rect 23550 23266 23602 23278
rect 23550 23202 23602 23214
rect 25902 23266 25954 23278
rect 25902 23202 25954 23214
rect 26014 23266 26066 23278
rect 26014 23202 26066 23214
rect 27358 23266 27410 23278
rect 27358 23202 27410 23214
rect 27694 23266 27746 23278
rect 27694 23202 27746 23214
rect 28030 23266 28082 23278
rect 28030 23202 28082 23214
rect 28254 23266 28306 23278
rect 28254 23202 28306 23214
rect 30494 23266 30546 23278
rect 31614 23266 31666 23278
rect 31154 23214 31166 23266
rect 31218 23214 31230 23266
rect 30494 23202 30546 23214
rect 31614 23202 31666 23214
rect 31726 23266 31778 23278
rect 31726 23202 31778 23214
rect 33518 23266 33570 23278
rect 33518 23202 33570 23214
rect 34862 23266 34914 23278
rect 34862 23202 34914 23214
rect 35310 23266 35362 23278
rect 35310 23202 35362 23214
rect 35758 23266 35810 23278
rect 37774 23266 37826 23278
rect 36754 23214 36766 23266
rect 36818 23214 36830 23266
rect 35758 23202 35810 23214
rect 37774 23202 37826 23214
rect 37886 23266 37938 23278
rect 37886 23202 37938 23214
rect 39678 23266 39730 23278
rect 39678 23202 39730 23214
rect 41470 23266 41522 23278
rect 41470 23202 41522 23214
rect 45278 23266 45330 23278
rect 45278 23202 45330 23214
rect 47406 23266 47458 23278
rect 47406 23202 47458 23214
rect 50654 23266 50706 23278
rect 50654 23202 50706 23214
rect 51550 23266 51602 23278
rect 55010 23214 55022 23266
rect 55074 23214 55086 23266
rect 51550 23202 51602 23214
rect 8766 23154 8818 23166
rect 13694 23154 13746 23166
rect 1810 23102 1822 23154
rect 1874 23102 1886 23154
rect 5170 23102 5182 23154
rect 5234 23102 5246 23154
rect 9762 23102 9774 23154
rect 9826 23102 9838 23154
rect 8766 23090 8818 23102
rect 13694 23090 13746 23102
rect 14142 23154 14194 23166
rect 14142 23090 14194 23102
rect 14254 23154 14306 23166
rect 14254 23090 14306 23102
rect 14926 23154 14978 23166
rect 14926 23090 14978 23102
rect 15262 23154 15314 23166
rect 15262 23090 15314 23102
rect 15598 23154 15650 23166
rect 15598 23090 15650 23102
rect 15934 23154 15986 23166
rect 29486 23154 29538 23166
rect 17378 23102 17390 23154
rect 17442 23102 17454 23154
rect 20850 23102 20862 23154
rect 20914 23102 20926 23154
rect 24098 23102 24110 23154
rect 24162 23102 24174 23154
rect 26674 23102 26686 23154
rect 26738 23102 26750 23154
rect 15934 23090 15986 23102
rect 29486 23090 29538 23102
rect 30830 23154 30882 23166
rect 30830 23090 30882 23102
rect 32510 23154 32562 23166
rect 32510 23090 32562 23102
rect 32958 23154 33010 23166
rect 32958 23090 33010 23102
rect 34302 23154 34354 23166
rect 34302 23090 34354 23102
rect 35198 23154 35250 23166
rect 36430 23154 36482 23166
rect 43822 23154 43874 23166
rect 36082 23102 36094 23154
rect 36146 23102 36158 23154
rect 39218 23102 39230 23154
rect 39282 23102 39294 23154
rect 43250 23102 43262 23154
rect 43314 23102 43326 23154
rect 35198 23090 35250 23102
rect 36430 23090 36482 23102
rect 43822 23090 43874 23102
rect 45166 23154 45218 23166
rect 45166 23090 45218 23102
rect 45390 23154 45442 23166
rect 45390 23090 45442 23102
rect 47294 23154 47346 23166
rect 47294 23090 47346 23102
rect 48078 23154 48130 23166
rect 51326 23154 51378 23166
rect 49074 23102 49086 23154
rect 49138 23102 49150 23154
rect 54338 23102 54350 23154
rect 54402 23102 54414 23154
rect 54898 23102 54910 23154
rect 54962 23102 54974 23154
rect 56914 23102 56926 23154
rect 56978 23102 56990 23154
rect 48078 23090 48130 23102
rect 51326 23090 51378 23102
rect 13358 23042 13410 23054
rect 21982 23042 22034 23054
rect 25566 23042 25618 23054
rect 27806 23042 27858 23054
rect 37214 23042 37266 23054
rect 2482 22990 2494 23042
rect 2546 22990 2558 23042
rect 4610 22990 4622 23042
rect 4674 22990 4686 23042
rect 5954 22990 5966 23042
rect 6018 22990 6030 23042
rect 8082 22990 8094 23042
rect 8146 22990 8158 23042
rect 10546 22990 10558 23042
rect 10610 22990 10622 23042
rect 12674 22990 12686 23042
rect 12738 22990 12750 23042
rect 18162 22990 18174 23042
rect 18226 22990 18238 23042
rect 20290 22990 20302 23042
rect 20354 22990 20366 23042
rect 24434 22990 24446 23042
rect 24498 22990 24510 23042
rect 26898 22990 26910 23042
rect 26962 22990 26974 23042
rect 30258 22990 30270 23042
rect 30322 22990 30334 23042
rect 13358 22978 13410 22990
rect 21982 22978 22034 22990
rect 25566 22978 25618 22990
rect 27806 22978 27858 22990
rect 37214 22978 37266 22990
rect 38334 23042 38386 23054
rect 41582 23042 41634 23054
rect 38770 22990 38782 23042
rect 38834 22990 38846 23042
rect 38334 22978 38386 22990
rect 41582 22978 41634 22990
rect 46062 23042 46114 23054
rect 46062 22978 46114 22990
rect 46958 23042 47010 23054
rect 46958 22978 47010 22990
rect 48190 23042 48242 23054
rect 49758 23042 49810 23054
rect 48850 22990 48862 23042
rect 48914 22990 48926 23042
rect 48190 22978 48242 22990
rect 49758 22978 49810 22990
rect 52446 23042 52498 23054
rect 57598 23042 57650 23054
rect 54786 22990 54798 23042
rect 54850 22990 54862 23042
rect 56690 22990 56702 23042
rect 56754 22990 56766 23042
rect 52446 22978 52498 22990
rect 57598 22978 57650 22990
rect 25902 22930 25954 22942
rect 25902 22866 25954 22878
rect 29262 22930 29314 22942
rect 29262 22866 29314 22878
rect 33182 22930 33234 22942
rect 33182 22866 33234 22878
rect 41694 22930 41746 22942
rect 41694 22866 41746 22878
rect 44046 22930 44098 22942
rect 51886 22930 51938 22942
rect 44370 22878 44382 22930
rect 44434 22878 44446 22930
rect 44046 22866 44098 22878
rect 51886 22866 51938 22878
rect 52222 22930 52274 22942
rect 52222 22866 52274 22878
rect 1344 22762 58576 22796
rect 1344 22710 8367 22762
rect 8419 22710 8471 22762
rect 8523 22710 8575 22762
rect 8627 22710 22674 22762
rect 22726 22710 22778 22762
rect 22830 22710 22882 22762
rect 22934 22710 36981 22762
rect 37033 22710 37085 22762
rect 37137 22710 37189 22762
rect 37241 22710 51288 22762
rect 51340 22710 51392 22762
rect 51444 22710 51496 22762
rect 51548 22710 58576 22762
rect 1344 22676 58576 22710
rect 7758 22594 7810 22606
rect 7758 22530 7810 22542
rect 8094 22594 8146 22606
rect 37774 22594 37826 22606
rect 27234 22542 27246 22594
rect 27298 22542 27310 22594
rect 8094 22530 8146 22542
rect 37774 22530 37826 22542
rect 38222 22594 38274 22606
rect 38222 22530 38274 22542
rect 48526 22594 48578 22606
rect 55010 22542 55022 22594
rect 55074 22542 55086 22594
rect 56130 22542 56142 22594
rect 56194 22542 56206 22594
rect 48526 22530 48578 22542
rect 3054 22482 3106 22494
rect 3054 22418 3106 22430
rect 6078 22482 6130 22494
rect 6078 22418 6130 22430
rect 11006 22482 11058 22494
rect 11006 22418 11058 22430
rect 24110 22482 24162 22494
rect 24110 22418 24162 22430
rect 25006 22482 25058 22494
rect 25006 22418 25058 22430
rect 34750 22482 34802 22494
rect 34750 22418 34802 22430
rect 35646 22482 35698 22494
rect 35646 22418 35698 22430
rect 38782 22482 38834 22494
rect 38782 22418 38834 22430
rect 39902 22482 39954 22494
rect 39902 22418 39954 22430
rect 43262 22482 43314 22494
rect 54450 22430 54462 22482
rect 54514 22430 54526 22482
rect 55906 22430 55918 22482
rect 55970 22430 55982 22482
rect 43262 22418 43314 22430
rect 2942 22370 2994 22382
rect 2942 22306 2994 22318
rect 3278 22370 3330 22382
rect 3278 22306 3330 22318
rect 3502 22370 3554 22382
rect 3502 22306 3554 22318
rect 4510 22370 4562 22382
rect 4510 22306 4562 22318
rect 6302 22370 6354 22382
rect 6302 22306 6354 22318
rect 10894 22370 10946 22382
rect 10894 22306 10946 22318
rect 11118 22370 11170 22382
rect 13022 22370 13074 22382
rect 11666 22318 11678 22370
rect 11730 22318 11742 22370
rect 11118 22306 11170 22318
rect 13022 22306 13074 22318
rect 14030 22370 14082 22382
rect 14030 22306 14082 22318
rect 14702 22370 14754 22382
rect 14702 22306 14754 22318
rect 15038 22370 15090 22382
rect 15038 22306 15090 22318
rect 15262 22370 15314 22382
rect 15262 22306 15314 22318
rect 15710 22370 15762 22382
rect 15710 22306 15762 22318
rect 16270 22370 16322 22382
rect 16270 22306 16322 22318
rect 21534 22370 21586 22382
rect 21534 22306 21586 22318
rect 22430 22370 22482 22382
rect 25790 22370 25842 22382
rect 22866 22318 22878 22370
rect 22930 22318 22942 22370
rect 22430 22306 22482 22318
rect 25790 22306 25842 22318
rect 26126 22370 26178 22382
rect 28366 22370 28418 22382
rect 26338 22318 26350 22370
rect 26402 22318 26414 22370
rect 27346 22318 27358 22370
rect 27410 22318 27422 22370
rect 27570 22318 27582 22370
rect 27634 22318 27646 22370
rect 26126 22306 26178 22318
rect 28366 22306 28418 22318
rect 28590 22370 28642 22382
rect 31166 22370 31218 22382
rect 33406 22370 33458 22382
rect 36206 22370 36258 22382
rect 30146 22318 30158 22370
rect 30210 22318 30222 22370
rect 30818 22318 30830 22370
rect 30882 22318 30894 22370
rect 32834 22318 32846 22370
rect 32898 22318 32910 22370
rect 33954 22318 33966 22370
rect 34018 22318 34030 22370
rect 28590 22306 28642 22318
rect 31166 22306 31218 22318
rect 33406 22306 33458 22318
rect 36206 22306 36258 22318
rect 37326 22370 37378 22382
rect 37326 22306 37378 22318
rect 38334 22370 38386 22382
rect 44382 22370 44434 22382
rect 41682 22318 41694 22370
rect 41746 22318 41758 22370
rect 42578 22318 42590 22370
rect 42642 22318 42654 22370
rect 38334 22306 38386 22318
rect 44382 22306 44434 22318
rect 45166 22370 45218 22382
rect 45166 22306 45218 22318
rect 45502 22370 45554 22382
rect 45502 22306 45554 22318
rect 46510 22370 46562 22382
rect 46510 22306 46562 22318
rect 49870 22370 49922 22382
rect 49870 22306 49922 22318
rect 50430 22370 50482 22382
rect 50430 22306 50482 22318
rect 50654 22370 50706 22382
rect 51550 22370 51602 22382
rect 52894 22370 52946 22382
rect 50978 22318 50990 22370
rect 51042 22318 51054 22370
rect 51874 22318 51886 22370
rect 51938 22318 51950 22370
rect 50654 22306 50706 22318
rect 51550 22306 51602 22318
rect 52894 22306 52946 22318
rect 53230 22370 53282 22382
rect 57038 22370 57090 22382
rect 54226 22318 54238 22370
rect 54290 22318 54302 22370
rect 55794 22318 55806 22370
rect 55858 22318 55870 22370
rect 53230 22306 53282 22318
rect 57038 22306 57090 22318
rect 57262 22370 57314 22382
rect 57262 22306 57314 22318
rect 2606 22258 2658 22270
rect 2606 22194 2658 22206
rect 4174 22258 4226 22270
rect 4174 22194 4226 22206
rect 5966 22258 6018 22270
rect 5966 22194 6018 22206
rect 6526 22258 6578 22270
rect 8990 22258 9042 22270
rect 7074 22206 7086 22258
rect 7138 22206 7150 22258
rect 7410 22206 7422 22258
rect 7474 22206 7486 22258
rect 6526 22194 6578 22206
rect 8990 22194 9042 22206
rect 9326 22258 9378 22270
rect 9326 22194 9378 22206
rect 10558 22258 10610 22270
rect 10558 22194 10610 22206
rect 12686 22258 12738 22270
rect 12686 22194 12738 22206
rect 13694 22258 13746 22270
rect 14590 22258 14642 22270
rect 13694 22194 13746 22206
rect 14254 22202 14306 22214
rect 2270 22146 2322 22158
rect 2270 22082 2322 22094
rect 9774 22146 9826 22158
rect 9774 22082 9826 22094
rect 10334 22146 10386 22158
rect 12350 22146 12402 22158
rect 11442 22094 11454 22146
rect 11506 22094 11518 22146
rect 10334 22082 10386 22094
rect 12350 22082 12402 22094
rect 12798 22146 12850 22158
rect 12798 22082 12850 22094
rect 13806 22146 13858 22158
rect 14590 22194 14642 22206
rect 15934 22258 15986 22270
rect 15934 22194 15986 22206
rect 19406 22258 19458 22270
rect 23998 22258 24050 22270
rect 22082 22206 22094 22258
rect 22146 22206 22158 22258
rect 23090 22206 23102 22258
rect 23154 22206 23166 22258
rect 19406 22194 19458 22206
rect 23998 22194 24050 22206
rect 24894 22258 24946 22270
rect 24894 22194 24946 22206
rect 29038 22258 29090 22270
rect 31390 22258 31442 22270
rect 29362 22206 29374 22258
rect 29426 22206 29438 22258
rect 29922 22206 29934 22258
rect 29986 22206 29998 22258
rect 30594 22206 30606 22258
rect 30658 22206 30670 22258
rect 29038 22194 29090 22206
rect 31390 22194 31442 22206
rect 31502 22258 31554 22270
rect 33294 22258 33346 22270
rect 37662 22258 37714 22270
rect 32050 22206 32062 22258
rect 32114 22206 32126 22258
rect 32610 22206 32622 22258
rect 32674 22206 32686 22258
rect 36978 22206 36990 22258
rect 37042 22206 37054 22258
rect 31502 22194 31554 22206
rect 33294 22194 33346 22206
rect 37662 22194 37714 22206
rect 39454 22258 39506 22270
rect 39454 22194 39506 22206
rect 40462 22258 40514 22270
rect 45838 22258 45890 22270
rect 41346 22206 41358 22258
rect 41410 22206 41422 22258
rect 44818 22206 44830 22258
rect 44882 22206 44894 22258
rect 40462 22194 40514 22206
rect 45838 22194 45890 22206
rect 46174 22258 46226 22270
rect 46174 22194 46226 22206
rect 47406 22258 47458 22270
rect 48526 22258 48578 22270
rect 48066 22206 48078 22258
rect 48130 22206 48142 22258
rect 47406 22194 47458 22206
rect 48526 22194 48578 22206
rect 48638 22258 48690 22270
rect 48638 22194 48690 22206
rect 48974 22258 49026 22270
rect 48974 22194 49026 22206
rect 49310 22258 49362 22270
rect 49310 22194 49362 22206
rect 14254 22138 14306 22150
rect 14366 22146 14418 22158
rect 13806 22082 13858 22094
rect 14366 22082 14418 22094
rect 15038 22146 15090 22158
rect 15038 22082 15090 22094
rect 16158 22146 16210 22158
rect 16158 22082 16210 22094
rect 16718 22146 16770 22158
rect 16718 22082 16770 22094
rect 20302 22146 20354 22158
rect 20302 22082 20354 22094
rect 21646 22146 21698 22158
rect 21646 22082 21698 22094
rect 21870 22146 21922 22158
rect 21870 22082 21922 22094
rect 24222 22146 24274 22158
rect 24222 22082 24274 22094
rect 24446 22146 24498 22158
rect 24446 22082 24498 22094
rect 25118 22146 25170 22158
rect 25118 22082 25170 22094
rect 25342 22146 25394 22158
rect 25342 22082 25394 22094
rect 25902 22146 25954 22158
rect 35310 22146 35362 22158
rect 28018 22094 28030 22146
rect 28082 22094 28094 22146
rect 32274 22094 32286 22146
rect 32338 22094 32350 22146
rect 25902 22082 25954 22094
rect 35310 22082 35362 22094
rect 38222 22146 38274 22158
rect 38222 22082 38274 22094
rect 39118 22146 39170 22158
rect 39118 22082 39170 22094
rect 39342 22146 39394 22158
rect 39342 22082 39394 22094
rect 40574 22146 40626 22158
rect 40574 22082 40626 22094
rect 40798 22146 40850 22158
rect 40798 22082 40850 22094
rect 46286 22146 46338 22158
rect 47742 22146 47794 22158
rect 47058 22094 47070 22146
rect 47122 22094 47134 22146
rect 46286 22082 46338 22094
rect 47742 22082 47794 22094
rect 49982 22146 50034 22158
rect 49982 22082 50034 22094
rect 50206 22146 50258 22158
rect 50206 22082 50258 22094
rect 51326 22146 51378 22158
rect 51326 22082 51378 22094
rect 51438 22146 51490 22158
rect 57586 22094 57598 22146
rect 57650 22094 57662 22146
rect 51438 22082 51490 22094
rect 1344 21978 58731 22012
rect 1344 21926 15520 21978
rect 15572 21926 15624 21978
rect 15676 21926 15728 21978
rect 15780 21926 29827 21978
rect 29879 21926 29931 21978
rect 29983 21926 30035 21978
rect 30087 21926 44134 21978
rect 44186 21926 44238 21978
rect 44290 21926 44342 21978
rect 44394 21926 58441 21978
rect 58493 21926 58545 21978
rect 58597 21926 58649 21978
rect 58701 21926 58731 21978
rect 1344 21892 58731 21926
rect 1934 21810 1986 21822
rect 3166 21810 3218 21822
rect 2818 21758 2830 21810
rect 2882 21758 2894 21810
rect 1934 21746 1986 21758
rect 3166 21746 3218 21758
rect 4846 21810 4898 21822
rect 4846 21746 4898 21758
rect 9998 21810 10050 21822
rect 15262 21810 15314 21822
rect 14690 21758 14702 21810
rect 14754 21758 14766 21810
rect 9998 21746 10050 21758
rect 15262 21746 15314 21758
rect 18398 21810 18450 21822
rect 18398 21746 18450 21758
rect 18958 21810 19010 21822
rect 18958 21746 19010 21758
rect 22766 21810 22818 21822
rect 22766 21746 22818 21758
rect 22990 21810 23042 21822
rect 22990 21746 23042 21758
rect 25790 21810 25842 21822
rect 25790 21746 25842 21758
rect 25902 21810 25954 21822
rect 25902 21746 25954 21758
rect 26126 21810 26178 21822
rect 26126 21746 26178 21758
rect 31614 21810 31666 21822
rect 31614 21746 31666 21758
rect 32398 21810 32450 21822
rect 32398 21746 32450 21758
rect 33630 21810 33682 21822
rect 33630 21746 33682 21758
rect 33854 21810 33906 21822
rect 38110 21810 38162 21822
rect 41246 21810 41298 21822
rect 34402 21758 34414 21810
rect 34466 21758 34478 21810
rect 37762 21758 37774 21810
rect 37826 21758 37838 21810
rect 39778 21758 39790 21810
rect 39842 21758 39854 21810
rect 33854 21746 33906 21758
rect 38110 21746 38162 21758
rect 41246 21746 41298 21758
rect 46174 21810 46226 21822
rect 46174 21746 46226 21758
rect 46846 21810 46898 21822
rect 46846 21746 46898 21758
rect 51326 21810 51378 21822
rect 54350 21810 54402 21822
rect 53666 21758 53678 21810
rect 53730 21758 53742 21810
rect 51326 21746 51378 21758
rect 54350 21746 54402 21758
rect 55694 21810 55746 21822
rect 57922 21758 57934 21810
rect 57986 21758 57998 21810
rect 55694 21746 55746 21758
rect 2494 21698 2546 21710
rect 2146 21646 2158 21698
rect 2210 21646 2222 21698
rect 2494 21634 2546 21646
rect 8654 21698 8706 21710
rect 8654 21634 8706 21646
rect 10110 21698 10162 21710
rect 10110 21634 10162 21646
rect 14030 21698 14082 21710
rect 14030 21634 14082 21646
rect 14366 21698 14418 21710
rect 14366 21634 14418 21646
rect 15486 21698 15538 21710
rect 15486 21634 15538 21646
rect 15598 21698 15650 21710
rect 15598 21634 15650 21646
rect 15934 21698 15986 21710
rect 15934 21634 15986 21646
rect 16046 21698 16098 21710
rect 16046 21634 16098 21646
rect 17502 21698 17554 21710
rect 17502 21634 17554 21646
rect 18062 21698 18114 21710
rect 18062 21634 18114 21646
rect 18510 21698 18562 21710
rect 18510 21634 18562 21646
rect 19070 21698 19122 21710
rect 36878 21698 36930 21710
rect 35410 21646 35422 21698
rect 35474 21646 35486 21698
rect 36082 21646 36094 21698
rect 36146 21646 36158 21698
rect 19070 21634 19122 21646
rect 36878 21634 36930 21646
rect 38446 21698 38498 21710
rect 44382 21698 44434 21710
rect 43810 21646 43822 21698
rect 43874 21646 43886 21698
rect 38446 21634 38498 21646
rect 44382 21634 44434 21646
rect 47406 21698 47458 21710
rect 47406 21634 47458 21646
rect 47518 21698 47570 21710
rect 47518 21634 47570 21646
rect 47966 21698 48018 21710
rect 47966 21634 48018 21646
rect 48078 21698 48130 21710
rect 50990 21698 51042 21710
rect 50642 21646 50654 21698
rect 50706 21646 50718 21698
rect 48078 21634 48130 21646
rect 50990 21634 51042 21646
rect 51102 21698 51154 21710
rect 54462 21698 54514 21710
rect 51986 21646 51998 21698
rect 52050 21646 52062 21698
rect 51102 21634 51154 21646
rect 54462 21634 54514 21646
rect 55918 21698 55970 21710
rect 57250 21646 57262 21698
rect 57314 21646 57326 21698
rect 55918 21634 55970 21646
rect 8206 21586 8258 21598
rect 16606 21586 16658 21598
rect 23438 21586 23490 21598
rect 4162 21534 4174 21586
rect 4226 21534 4238 21586
rect 4610 21534 4622 21586
rect 4674 21534 4686 21586
rect 10434 21534 10446 21586
rect 10498 21534 10510 21586
rect 14914 21534 14926 21586
rect 14978 21534 14990 21586
rect 19506 21534 19518 21586
rect 19570 21534 19582 21586
rect 8206 21522 8258 21534
rect 16606 21522 16658 21534
rect 23438 21522 23490 21534
rect 26238 21586 26290 21598
rect 31950 21586 32002 21598
rect 27234 21534 27246 21586
rect 27298 21534 27310 21586
rect 28130 21534 28142 21586
rect 28194 21534 28206 21586
rect 28578 21534 28590 21586
rect 28642 21534 28654 21586
rect 29698 21534 29710 21586
rect 29762 21534 29774 21586
rect 26238 21522 26290 21534
rect 31950 21522 32002 21534
rect 32174 21586 32226 21598
rect 32174 21522 32226 21534
rect 32510 21586 32562 21598
rect 35086 21586 35138 21598
rect 36766 21586 36818 21598
rect 33058 21534 33070 21586
rect 33122 21534 33134 21586
rect 33394 21534 33406 21586
rect 33458 21534 33470 21586
rect 34626 21534 34638 21586
rect 34690 21534 34702 21586
rect 36194 21534 36206 21586
rect 36258 21534 36270 21586
rect 32510 21522 32562 21534
rect 35086 21522 35138 21534
rect 36766 21522 36818 21534
rect 37102 21586 37154 21598
rect 40126 21586 40178 21598
rect 39106 21534 39118 21586
rect 39170 21534 39182 21586
rect 37102 21522 37154 21534
rect 40126 21522 40178 21534
rect 41022 21586 41074 21598
rect 41022 21522 41074 21534
rect 41358 21586 41410 21598
rect 41358 21522 41410 21534
rect 41582 21586 41634 21598
rect 44158 21586 44210 21598
rect 42354 21534 42366 21586
rect 42418 21534 42430 21586
rect 42914 21534 42926 21586
rect 42978 21534 42990 21586
rect 41582 21522 41634 21534
rect 44158 21522 44210 21534
rect 44494 21586 44546 21598
rect 44494 21522 44546 21534
rect 45166 21586 45218 21598
rect 45166 21522 45218 21534
rect 45838 21586 45890 21598
rect 45838 21522 45890 21534
rect 45950 21586 46002 21598
rect 45950 21522 46002 21534
rect 46286 21586 46338 21598
rect 46286 21522 46338 21534
rect 46734 21586 46786 21598
rect 46734 21522 46786 21534
rect 48302 21586 48354 21598
rect 49746 21534 49758 21586
rect 49810 21534 49822 21586
rect 50418 21534 50430 21586
rect 50482 21534 50494 21586
rect 52210 21534 52222 21586
rect 52274 21534 52286 21586
rect 53106 21534 53118 21586
rect 53170 21534 53182 21586
rect 57362 21534 57374 21586
rect 57426 21534 57438 21586
rect 57810 21534 57822 21586
rect 57874 21534 57886 21586
rect 48302 21522 48354 21534
rect 22878 21474 22930 21486
rect 4050 21422 4062 21474
rect 4114 21422 4126 21474
rect 7746 21422 7758 21474
rect 7810 21422 7822 21474
rect 11218 21422 11230 21474
rect 11282 21422 11294 21474
rect 13346 21422 13358 21474
rect 13410 21422 13422 21474
rect 20290 21422 20302 21474
rect 20354 21422 20366 21474
rect 22418 21422 22430 21474
rect 22482 21422 22494 21474
rect 22878 21410 22930 21422
rect 23774 21474 23826 21486
rect 37438 21474 37490 21486
rect 45390 21474 45442 21486
rect 26786 21422 26798 21474
rect 26850 21422 26862 21474
rect 30258 21422 30270 21474
rect 30322 21422 30334 21474
rect 33618 21422 33630 21474
rect 33682 21422 33694 21474
rect 36306 21422 36318 21474
rect 36370 21422 36382 21474
rect 39330 21422 39342 21474
rect 39394 21422 39406 21474
rect 44818 21422 44830 21474
rect 44882 21422 44894 21474
rect 23774 21410 23826 21422
rect 37438 21410 37490 21422
rect 45390 21410 45442 21422
rect 46062 21474 46114 21486
rect 48850 21422 48862 21474
rect 48914 21422 48926 21474
rect 55570 21422 55582 21474
rect 55634 21422 55646 21474
rect 46062 21410 46114 21422
rect 3838 21362 3890 21374
rect 3838 21298 3890 21310
rect 8542 21362 8594 21374
rect 8542 21298 8594 21310
rect 8878 21362 8930 21374
rect 8878 21298 8930 21310
rect 9998 21362 10050 21374
rect 9998 21298 10050 21310
rect 16046 21362 16098 21374
rect 16046 21298 16098 21310
rect 18398 21362 18450 21374
rect 18398 21298 18450 21310
rect 18958 21362 19010 21374
rect 18958 21298 19010 21310
rect 46846 21362 46898 21374
rect 46846 21298 46898 21310
rect 47518 21362 47570 21374
rect 47518 21298 47570 21310
rect 54238 21362 54290 21374
rect 54238 21298 54290 21310
rect 1344 21194 58576 21228
rect 1344 21142 8367 21194
rect 8419 21142 8471 21194
rect 8523 21142 8575 21194
rect 8627 21142 22674 21194
rect 22726 21142 22778 21194
rect 22830 21142 22882 21194
rect 22934 21142 36981 21194
rect 37033 21142 37085 21194
rect 37137 21142 37189 21194
rect 37241 21142 51288 21194
rect 51340 21142 51392 21194
rect 51444 21142 51496 21194
rect 51548 21142 58576 21194
rect 1344 21108 58576 21142
rect 9102 21026 9154 21038
rect 9102 20962 9154 20974
rect 9438 21026 9490 21038
rect 9438 20962 9490 20974
rect 16270 21026 16322 21038
rect 16270 20962 16322 20974
rect 20302 21026 20354 21038
rect 20302 20962 20354 20974
rect 8878 20914 8930 20926
rect 4610 20862 4622 20914
rect 4674 20862 4686 20914
rect 8530 20862 8542 20914
rect 8594 20862 8606 20914
rect 8878 20850 8930 20862
rect 10670 20914 10722 20926
rect 32062 20914 32114 20926
rect 17378 20862 17390 20914
rect 17442 20862 17454 20914
rect 19506 20862 19518 20914
rect 19570 20862 19582 20914
rect 21858 20862 21870 20914
rect 21922 20862 21934 20914
rect 26450 20862 26462 20914
rect 26514 20862 26526 20914
rect 10670 20850 10722 20862
rect 32062 20850 32114 20862
rect 32622 20914 32674 20926
rect 34974 20914 35026 20926
rect 41470 20914 41522 20926
rect 33842 20862 33854 20914
rect 33906 20862 33918 20914
rect 37426 20862 37438 20914
rect 37490 20862 37502 20914
rect 32622 20850 32674 20862
rect 34974 20850 35026 20862
rect 41470 20850 41522 20862
rect 46398 20914 46450 20926
rect 46398 20850 46450 20862
rect 48526 20914 48578 20926
rect 48526 20850 48578 20862
rect 51550 20914 51602 20926
rect 51550 20850 51602 20862
rect 53454 20914 53506 20926
rect 53890 20862 53902 20914
rect 53954 20862 53966 20914
rect 57026 20862 57038 20914
rect 57090 20862 57102 20914
rect 58034 20862 58046 20914
rect 58098 20862 58110 20914
rect 53454 20850 53506 20862
rect 1810 20762 1822 20814
rect 1874 20762 1886 20814
rect 10894 20802 10946 20814
rect 5618 20750 5630 20802
rect 5682 20750 5694 20802
rect 10894 20738 10946 20750
rect 11342 20802 11394 20814
rect 11342 20738 11394 20750
rect 11454 20802 11506 20814
rect 14814 20802 14866 20814
rect 14130 20750 14142 20802
rect 14194 20750 14206 20802
rect 11454 20738 11506 20750
rect 14814 20738 14866 20750
rect 15038 20802 15090 20814
rect 15038 20738 15090 20750
rect 15374 20802 15426 20814
rect 32734 20802 32786 20814
rect 16258 20750 16270 20802
rect 16322 20750 16334 20802
rect 16594 20750 16606 20802
rect 16658 20750 16670 20802
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 20626 20750 20638 20802
rect 20690 20750 20702 20802
rect 21970 20750 21982 20802
rect 22034 20750 22046 20802
rect 28466 20750 28478 20802
rect 28530 20750 28542 20802
rect 29138 20750 29150 20802
rect 29202 20750 29214 20802
rect 30258 20750 30270 20802
rect 30322 20750 30334 20802
rect 30482 20750 30494 20802
rect 30546 20750 30558 20802
rect 31826 20750 31838 20802
rect 31890 20750 31902 20802
rect 15374 20738 15426 20750
rect 32734 20738 32786 20750
rect 33182 20802 33234 20814
rect 36094 20802 36146 20814
rect 36430 20802 36482 20814
rect 40574 20802 40626 20814
rect 47182 20802 47234 20814
rect 49310 20802 49362 20814
rect 33506 20750 33518 20802
rect 33570 20750 33582 20802
rect 36306 20750 36318 20802
rect 36370 20750 36382 20802
rect 37314 20750 37326 20802
rect 37378 20750 37390 20802
rect 38098 20750 38110 20802
rect 38162 20750 38174 20802
rect 39442 20750 39454 20802
rect 39506 20750 39518 20802
rect 41234 20750 41246 20802
rect 41298 20750 41310 20802
rect 41906 20750 41918 20802
rect 41970 20750 41982 20802
rect 43922 20750 43934 20802
rect 43986 20750 43998 20802
rect 46050 20750 46062 20802
rect 46114 20750 46126 20802
rect 47842 20750 47854 20802
rect 47906 20750 47918 20802
rect 33182 20738 33234 20750
rect 36094 20738 36146 20750
rect 36430 20738 36482 20750
rect 40574 20738 40626 20750
rect 47182 20738 47234 20750
rect 49310 20738 49362 20750
rect 49646 20802 49698 20814
rect 49646 20738 49698 20750
rect 50318 20802 50370 20814
rect 50318 20738 50370 20750
rect 50654 20802 50706 20814
rect 50654 20738 50706 20750
rect 50878 20802 50930 20814
rect 50878 20738 50930 20750
rect 53118 20802 53170 20814
rect 55806 20802 55858 20814
rect 54114 20750 54126 20802
rect 54178 20750 54190 20802
rect 56914 20750 56926 20802
rect 56978 20750 56990 20802
rect 53118 20738 53170 20750
rect 55806 20738 55858 20750
rect 15934 20690 15986 20702
rect 2482 20638 2494 20690
rect 2546 20638 2558 20690
rect 6402 20638 6414 20690
rect 6466 20638 6478 20690
rect 12226 20638 12238 20690
rect 12290 20638 12302 20690
rect 15934 20626 15986 20638
rect 19854 20690 19906 20702
rect 19854 20626 19906 20638
rect 22654 20690 22706 20702
rect 32174 20690 32226 20702
rect 29250 20638 29262 20690
rect 29314 20638 29326 20690
rect 22654 20626 22706 20638
rect 32174 20626 32226 20638
rect 35422 20690 35474 20702
rect 40350 20690 40402 20702
rect 40002 20638 40014 20690
rect 40066 20638 40078 20690
rect 35422 20626 35474 20638
rect 40350 20626 40402 20638
rect 40910 20690 40962 20702
rect 40910 20626 40962 20638
rect 41582 20690 41634 20702
rect 46622 20690 46674 20702
rect 42018 20638 42030 20690
rect 42082 20638 42094 20690
rect 44146 20638 44158 20690
rect 44210 20638 44222 20690
rect 44930 20638 44942 20690
rect 44994 20638 45006 20690
rect 41582 20626 41634 20638
rect 46622 20626 46674 20638
rect 46734 20690 46786 20702
rect 46734 20626 46786 20638
rect 47630 20690 47682 20702
rect 47630 20626 47682 20638
rect 50990 20690 51042 20702
rect 50990 20626 51042 20638
rect 52894 20690 52946 20702
rect 52894 20626 52946 20638
rect 54798 20690 54850 20702
rect 54798 20626 54850 20638
rect 55358 20690 55410 20702
rect 55358 20626 55410 20638
rect 55470 20690 55522 20702
rect 55470 20626 55522 20638
rect 56142 20690 56194 20702
rect 56142 20626 56194 20638
rect 5070 20578 5122 20590
rect 5070 20514 5122 20526
rect 11230 20578 11282 20590
rect 11230 20514 11282 20526
rect 11902 20578 11954 20590
rect 11902 20514 11954 20526
rect 12686 20578 12738 20590
rect 12686 20514 12738 20526
rect 13694 20578 13746 20590
rect 13694 20514 13746 20526
rect 14366 20578 14418 20590
rect 14366 20514 14418 20526
rect 15038 20578 15090 20590
rect 32510 20578 32562 20590
rect 20178 20526 20190 20578
rect 20242 20526 20254 20578
rect 15038 20514 15090 20526
rect 32510 20514 32562 20526
rect 34414 20578 34466 20590
rect 34414 20514 34466 20526
rect 40798 20578 40850 20590
rect 40798 20514 40850 20526
rect 47406 20578 47458 20590
rect 47406 20514 47458 20526
rect 49198 20578 49250 20590
rect 49198 20514 49250 20526
rect 49422 20578 49474 20590
rect 49422 20514 49474 20526
rect 49534 20578 49586 20590
rect 49534 20514 49586 20526
rect 50430 20578 50482 20590
rect 50430 20514 50482 20526
rect 51214 20578 51266 20590
rect 51214 20514 51266 20526
rect 51998 20578 52050 20590
rect 51998 20514 52050 20526
rect 55694 20578 55746 20590
rect 55694 20514 55746 20526
rect 56030 20578 56082 20590
rect 56030 20514 56082 20526
rect 1344 20410 58731 20444
rect 1344 20358 15520 20410
rect 15572 20358 15624 20410
rect 15676 20358 15728 20410
rect 15780 20358 29827 20410
rect 29879 20358 29931 20410
rect 29983 20358 30035 20410
rect 30087 20358 44134 20410
rect 44186 20358 44238 20410
rect 44290 20358 44342 20410
rect 44394 20358 58441 20410
rect 58493 20358 58545 20410
rect 58597 20358 58649 20410
rect 58701 20358 58731 20410
rect 1344 20324 58731 20358
rect 1934 20242 1986 20254
rect 1934 20178 1986 20190
rect 3278 20242 3330 20254
rect 3278 20178 3330 20190
rect 18510 20242 18562 20254
rect 31054 20242 31106 20254
rect 19282 20190 19294 20242
rect 19346 20190 19358 20242
rect 30482 20190 30494 20242
rect 30546 20190 30558 20242
rect 18510 20178 18562 20190
rect 31054 20178 31106 20190
rect 40798 20242 40850 20254
rect 40798 20178 40850 20190
rect 50878 20242 50930 20254
rect 50878 20178 50930 20190
rect 51326 20242 51378 20254
rect 51326 20178 51378 20190
rect 54126 20242 54178 20254
rect 54126 20178 54178 20190
rect 3166 20130 3218 20142
rect 5630 20130 5682 20142
rect 11678 20130 11730 20142
rect 17502 20130 17554 20142
rect 2258 20078 2270 20130
rect 2322 20078 2334 20130
rect 4610 20078 4622 20130
rect 4674 20078 4686 20130
rect 4946 20078 4958 20130
rect 5010 20078 5022 20130
rect 8642 20078 8654 20130
rect 8706 20078 8718 20130
rect 14690 20078 14702 20130
rect 14754 20078 14766 20130
rect 3166 20066 3218 20078
rect 5630 20066 5682 20078
rect 11678 20066 11730 20078
rect 17502 20066 17554 20078
rect 17726 20130 17778 20142
rect 17726 20066 17778 20078
rect 18174 20130 18226 20142
rect 18174 20066 18226 20078
rect 19742 20130 19794 20142
rect 24670 20130 24722 20142
rect 31390 20130 31442 20142
rect 35982 20130 36034 20142
rect 21746 20078 21758 20130
rect 21810 20078 21822 20130
rect 24322 20078 24334 20130
rect 24386 20078 24398 20130
rect 26002 20078 26014 20130
rect 26066 20078 26078 20130
rect 34402 20078 34414 20130
rect 34466 20078 34478 20130
rect 19742 20066 19794 20078
rect 24670 20066 24722 20078
rect 31390 20066 31442 20078
rect 35982 20066 36034 20078
rect 37326 20130 37378 20142
rect 37326 20066 37378 20078
rect 38670 20130 38722 20142
rect 38670 20066 38722 20078
rect 39230 20130 39282 20142
rect 39230 20066 39282 20078
rect 41022 20130 41074 20142
rect 41022 20066 41074 20078
rect 42366 20130 42418 20142
rect 50318 20130 50370 20142
rect 47842 20078 47854 20130
rect 47906 20078 47918 20130
rect 42366 20066 42418 20078
rect 50318 20066 50370 20078
rect 53006 20130 53058 20142
rect 53006 20066 53058 20078
rect 53902 20130 53954 20142
rect 53902 20066 53954 20078
rect 55694 20130 55746 20142
rect 55694 20066 55746 20078
rect 55918 20130 55970 20142
rect 55918 20066 55970 20078
rect 3502 20018 3554 20030
rect 5294 20018 5346 20030
rect 3714 19966 3726 20018
rect 3778 19966 3790 20018
rect 3502 19954 3554 19966
rect 5294 19954 5346 19966
rect 8094 20018 8146 20030
rect 8094 19954 8146 19966
rect 8318 20018 8370 20030
rect 8318 19954 8370 19966
rect 10782 20018 10834 20030
rect 10782 19954 10834 19966
rect 11454 20018 11506 20030
rect 19406 20018 19458 20030
rect 22990 20018 23042 20030
rect 28702 20018 28754 20030
rect 30158 20018 30210 20030
rect 12450 19966 12462 20018
rect 12514 19966 12526 20018
rect 13906 19966 13918 20018
rect 13970 19966 13982 20018
rect 18946 19966 18958 20018
rect 19010 19966 19022 20018
rect 22306 19966 22318 20018
rect 22370 19966 22382 20018
rect 23314 19966 23326 20018
rect 23378 19966 23390 20018
rect 25218 19966 25230 20018
rect 25282 19966 25294 20018
rect 29362 19966 29374 20018
rect 29426 19966 29438 20018
rect 11454 19954 11506 19966
rect 19406 19954 19458 19966
rect 22990 19954 23042 19966
rect 28702 19954 28754 19966
rect 30158 19954 30210 19966
rect 33182 20018 33234 20030
rect 36430 20018 36482 20030
rect 37662 20018 37714 20030
rect 34626 19966 34638 20018
rect 34690 19966 34702 20018
rect 35298 19966 35310 20018
rect 35362 19966 35374 20018
rect 36642 19966 36654 20018
rect 36706 19966 36718 20018
rect 33182 19954 33234 19966
rect 36430 19954 36482 19966
rect 37662 19954 37714 19966
rect 38222 20018 38274 20030
rect 38222 19954 38274 19966
rect 38446 20018 38498 20030
rect 38446 19954 38498 19966
rect 38782 20018 38834 20030
rect 38782 19954 38834 19966
rect 39678 20018 39730 20030
rect 39678 19954 39730 19966
rect 41134 20018 41186 20030
rect 41134 19954 41186 19966
rect 42030 20018 42082 20030
rect 48750 20018 48802 20030
rect 43810 19966 43822 20018
rect 43874 19966 43886 20018
rect 44482 19966 44494 20018
rect 44546 19966 44558 20018
rect 46610 19966 46622 20018
rect 46674 19966 46686 20018
rect 48066 19966 48078 20018
rect 48130 19966 48142 20018
rect 42030 19954 42082 19966
rect 48750 19954 48802 19966
rect 48974 20018 49026 20030
rect 48974 19954 49026 19966
rect 49086 20018 49138 20030
rect 49086 19954 49138 19966
rect 49534 20018 49586 20030
rect 49534 19954 49586 19966
rect 49758 20018 49810 20030
rect 49758 19954 49810 19966
rect 50206 20018 50258 20030
rect 50206 19954 50258 19966
rect 50542 20018 50594 20030
rect 50542 19954 50594 19966
rect 52446 20018 52498 20030
rect 52446 19954 52498 19966
rect 52894 20018 52946 20030
rect 52894 19954 52946 19966
rect 53118 20018 53170 20030
rect 53118 19954 53170 19966
rect 56030 20018 56082 20030
rect 56030 19954 56082 19966
rect 56702 20018 56754 20030
rect 57026 19966 57038 20018
rect 57090 19966 57102 20018
rect 56702 19954 56754 19966
rect 2606 19906 2658 19918
rect 2606 19842 2658 19854
rect 6190 19906 6242 19918
rect 6190 19842 6242 19854
rect 6638 19906 6690 19918
rect 6638 19842 6690 19854
rect 7198 19906 7250 19918
rect 7198 19842 7250 19854
rect 9886 19906 9938 19918
rect 9886 19842 9938 19854
rect 10334 19906 10386 19918
rect 10334 19842 10386 19854
rect 10558 19906 10610 19918
rect 10558 19842 10610 19854
rect 11118 19906 11170 19918
rect 12910 19906 12962 19918
rect 11778 19854 11790 19906
rect 11842 19854 11854 19906
rect 11118 19842 11170 19854
rect 12910 19842 12962 19854
rect 13694 19906 13746 19918
rect 20190 19906 20242 19918
rect 16818 19854 16830 19906
rect 16882 19854 16894 19906
rect 13694 19842 13746 19854
rect 20190 19842 20242 19854
rect 20974 19906 21026 19918
rect 28590 19906 28642 19918
rect 28130 19854 28142 19906
rect 28194 19854 28206 19906
rect 20974 19842 21026 19854
rect 28590 19842 28642 19854
rect 29934 19906 29986 19918
rect 29934 19842 29986 19854
rect 32510 19906 32562 19918
rect 32510 19842 32562 19854
rect 40126 19906 40178 19918
rect 51774 19906 51826 19918
rect 56590 19906 56642 19918
rect 41794 19854 41806 19906
rect 41858 19854 41870 19906
rect 43362 19854 43374 19906
rect 43426 19854 43438 19906
rect 44706 19854 44718 19906
rect 44770 19854 44782 19906
rect 46050 19854 46062 19906
rect 46114 19854 46126 19906
rect 54226 19854 54238 19906
rect 54290 19854 54302 19906
rect 40126 19842 40178 19854
rect 51774 19842 51826 19854
rect 56590 19842 56642 19854
rect 2718 19794 2770 19806
rect 17838 19794 17890 19806
rect 32286 19794 32338 19806
rect 3714 19742 3726 19794
rect 3778 19742 3790 19794
rect 6850 19742 6862 19794
rect 6914 19791 6926 19794
rect 7186 19791 7198 19794
rect 6914 19745 7198 19791
rect 6914 19742 6926 19745
rect 7186 19742 7198 19745
rect 7250 19742 7262 19794
rect 8866 19742 8878 19794
rect 8930 19791 8942 19794
rect 9090 19791 9102 19794
rect 8930 19745 9102 19791
rect 8930 19742 8942 19745
rect 9090 19742 9102 19745
rect 9154 19742 9166 19794
rect 19170 19742 19182 19794
rect 19234 19742 19246 19794
rect 31938 19742 31950 19794
rect 32002 19742 32014 19794
rect 2718 19730 2770 19742
rect 17838 19730 17890 19742
rect 32286 19730 32338 19742
rect 33070 19794 33122 19806
rect 50754 19742 50766 19794
rect 50818 19791 50830 19794
rect 51762 19791 51774 19794
rect 50818 19745 51774 19791
rect 50818 19742 50830 19745
rect 51762 19742 51774 19745
rect 51826 19742 51838 19794
rect 33070 19730 33122 19742
rect 1344 19626 58576 19660
rect 1344 19574 8367 19626
rect 8419 19574 8471 19626
rect 8523 19574 8575 19626
rect 8627 19574 22674 19626
rect 22726 19574 22778 19626
rect 22830 19574 22882 19626
rect 22934 19574 36981 19626
rect 37033 19574 37085 19626
rect 37137 19574 37189 19626
rect 37241 19574 51288 19626
rect 51340 19574 51392 19626
rect 51444 19574 51496 19626
rect 51548 19574 58576 19626
rect 1344 19540 58576 19574
rect 8542 19458 8594 19470
rect 8542 19394 8594 19406
rect 8990 19458 9042 19470
rect 21646 19458 21698 19470
rect 11442 19406 11454 19458
rect 11506 19406 11518 19458
rect 16818 19406 16830 19458
rect 16882 19455 16894 19458
rect 17378 19455 17390 19458
rect 16882 19409 17390 19455
rect 16882 19406 16894 19409
rect 17378 19406 17390 19409
rect 17442 19406 17454 19458
rect 8990 19394 9042 19406
rect 21646 19394 21698 19406
rect 23438 19458 23490 19470
rect 34414 19458 34466 19470
rect 52110 19458 52162 19470
rect 53566 19458 53618 19470
rect 32722 19406 32734 19458
rect 32786 19406 32798 19458
rect 43922 19406 43934 19458
rect 43986 19406 43998 19458
rect 53218 19406 53230 19458
rect 53282 19406 53294 19458
rect 23438 19394 23490 19406
rect 34414 19394 34466 19406
rect 52110 19394 52162 19406
rect 53566 19394 53618 19406
rect 53902 19458 53954 19470
rect 57474 19406 57486 19458
rect 57538 19406 57550 19458
rect 53902 19394 53954 19406
rect 9998 19346 10050 19358
rect 16830 19346 16882 19358
rect 4610 19294 4622 19346
rect 4674 19294 4686 19346
rect 7186 19294 7198 19346
rect 7250 19294 7262 19346
rect 11666 19294 11678 19346
rect 11730 19294 11742 19346
rect 9998 19282 10050 19294
rect 16830 19282 16882 19294
rect 19854 19346 19906 19358
rect 23998 19346 24050 19358
rect 22754 19294 22766 19346
rect 22818 19294 22830 19346
rect 19854 19282 19906 19294
rect 23998 19282 24050 19294
rect 24446 19346 24498 19358
rect 24446 19282 24498 19294
rect 24894 19346 24946 19358
rect 28590 19346 28642 19358
rect 25442 19294 25454 19346
rect 25506 19294 25518 19346
rect 24894 19282 24946 19294
rect 28590 19282 28642 19294
rect 29262 19346 29314 19358
rect 29262 19282 29314 19294
rect 30270 19346 30322 19358
rect 30270 19282 30322 19294
rect 30606 19346 30658 19358
rect 31950 19346 32002 19358
rect 34078 19346 34130 19358
rect 31490 19294 31502 19346
rect 31554 19294 31566 19346
rect 32834 19294 32846 19346
rect 32898 19294 32910 19346
rect 30606 19282 30658 19294
rect 31950 19282 32002 19294
rect 34078 19282 34130 19294
rect 35982 19346 36034 19358
rect 40686 19346 40738 19358
rect 45166 19346 45218 19358
rect 37986 19294 37998 19346
rect 38050 19294 38062 19346
rect 40114 19294 40126 19346
rect 40178 19294 40190 19346
rect 42018 19294 42030 19346
rect 42082 19294 42094 19346
rect 35982 19282 36034 19294
rect 40686 19282 40738 19294
rect 45166 19282 45218 19294
rect 50206 19346 50258 19358
rect 50206 19282 50258 19294
rect 51550 19346 51602 19358
rect 51550 19282 51602 19294
rect 52670 19346 52722 19358
rect 56254 19346 56306 19358
rect 55010 19294 55022 19346
rect 55074 19294 55086 19346
rect 56914 19294 56926 19346
rect 56978 19294 56990 19346
rect 52670 19282 52722 19294
rect 56254 19282 56306 19294
rect 5742 19234 5794 19246
rect 1698 19182 1710 19234
rect 1762 19182 1774 19234
rect 5742 19170 5794 19182
rect 6526 19234 6578 19246
rect 9214 19234 9266 19246
rect 6850 19182 6862 19234
rect 6914 19182 6926 19234
rect 8082 19182 8094 19234
rect 8146 19182 8158 19234
rect 6526 19170 6578 19182
rect 9214 19170 9266 19182
rect 9438 19234 9490 19246
rect 9438 19170 9490 19182
rect 10670 19234 10722 19246
rect 10670 19170 10722 19182
rect 11118 19234 11170 19246
rect 13470 19234 13522 19246
rect 11554 19182 11566 19234
rect 11618 19182 11630 19234
rect 12562 19182 12574 19234
rect 12626 19182 12638 19234
rect 11118 19170 11170 19182
rect 13470 19170 13522 19182
rect 13806 19234 13858 19246
rect 13806 19170 13858 19182
rect 14030 19234 14082 19246
rect 14030 19170 14082 19182
rect 17278 19234 17330 19246
rect 19518 19234 19570 19246
rect 19058 19182 19070 19234
rect 19122 19182 19134 19234
rect 17278 19170 17330 19182
rect 19518 19170 19570 19182
rect 20078 19234 20130 19246
rect 23774 19234 23826 19246
rect 26462 19234 26514 19246
rect 28478 19234 28530 19246
rect 22866 19182 22878 19234
rect 22930 19182 22942 19234
rect 25778 19182 25790 19234
rect 25842 19182 25854 19234
rect 28130 19182 28142 19234
rect 28194 19182 28206 19234
rect 20078 19170 20130 19182
rect 23774 19170 23826 19182
rect 26462 19170 26514 19182
rect 28478 19170 28530 19182
rect 29038 19234 29090 19246
rect 35758 19234 35810 19246
rect 31266 19182 31278 19234
rect 31330 19182 31342 19234
rect 33058 19182 33070 19234
rect 33122 19182 33134 19234
rect 33842 19182 33854 19234
rect 33906 19182 33918 19234
rect 35298 19182 35310 19234
rect 35362 19182 35374 19234
rect 29038 19170 29090 19182
rect 35758 19170 35810 19182
rect 36206 19234 36258 19246
rect 47854 19234 47906 19246
rect 37202 19182 37214 19234
rect 37266 19182 37278 19234
rect 41122 19182 41134 19234
rect 41186 19182 41198 19234
rect 42242 19182 42254 19234
rect 42306 19182 42318 19234
rect 43250 19182 43262 19234
rect 43314 19182 43326 19234
rect 36206 19170 36258 19182
rect 47854 19170 47906 19182
rect 48190 19234 48242 19246
rect 50766 19234 50818 19246
rect 48850 19182 48862 19234
rect 48914 19182 48926 19234
rect 49522 19182 49534 19234
rect 49586 19182 49598 19234
rect 48190 19170 48242 19182
rect 50766 19170 50818 19182
rect 51774 19234 51826 19246
rect 51774 19170 51826 19182
rect 52894 19234 52946 19246
rect 55470 19234 55522 19246
rect 55122 19182 55134 19234
rect 55186 19182 55198 19234
rect 55682 19182 55694 19234
rect 55746 19182 55758 19234
rect 56802 19182 56814 19234
rect 56866 19182 56878 19234
rect 52894 19170 52946 19182
rect 55470 19170 55522 19182
rect 6078 19122 6130 19134
rect 7534 19122 7586 19134
rect 2482 19070 2494 19122
rect 2546 19070 2558 19122
rect 6290 19070 6302 19122
rect 6354 19070 6366 19122
rect 6078 19058 6130 19070
rect 7534 19058 7586 19070
rect 8318 19122 8370 19134
rect 8318 19058 8370 19070
rect 9886 19122 9938 19134
rect 9886 19058 9938 19070
rect 10334 19122 10386 19134
rect 10334 19058 10386 19070
rect 10446 19122 10498 19134
rect 14590 19122 14642 19134
rect 12786 19070 12798 19122
rect 12850 19070 12862 19122
rect 10446 19058 10498 19070
rect 14590 19058 14642 19070
rect 14702 19122 14754 19134
rect 14702 19058 14754 19070
rect 15822 19122 15874 19134
rect 15822 19058 15874 19070
rect 17614 19122 17666 19134
rect 17614 19058 17666 19070
rect 26910 19122 26962 19134
rect 26910 19058 26962 19070
rect 29486 19122 29538 19134
rect 29486 19058 29538 19070
rect 29710 19122 29762 19134
rect 29710 19058 29762 19070
rect 34638 19122 34690 19134
rect 34638 19058 34690 19070
rect 36430 19122 36482 19134
rect 36430 19058 36482 19070
rect 46286 19122 46338 19134
rect 46286 19058 46338 19070
rect 46622 19122 46674 19134
rect 46622 19058 46674 19070
rect 46958 19122 47010 19134
rect 46958 19058 47010 19070
rect 47294 19122 47346 19134
rect 47294 19058 47346 19070
rect 47406 19122 47458 19134
rect 47406 19058 47458 19070
rect 47966 19122 48018 19134
rect 50878 19122 50930 19134
rect 49746 19070 49758 19122
rect 49810 19070 49822 19122
rect 47966 19058 48018 19070
rect 50878 19058 50930 19070
rect 53790 19122 53842 19134
rect 53790 19058 53842 19070
rect 54798 19122 54850 19134
rect 54798 19058 54850 19070
rect 5070 19010 5122 19022
rect 7310 19010 7362 19022
rect 6402 18958 6414 19010
rect 6466 18958 6478 19010
rect 5070 18946 5122 18958
rect 7310 18946 7362 18958
rect 13918 19010 13970 19022
rect 13918 18946 13970 18958
rect 14366 19010 14418 19022
rect 14366 18946 14418 18958
rect 15486 19010 15538 19022
rect 15486 18946 15538 18958
rect 15934 19010 15986 19022
rect 15934 18946 15986 18958
rect 16158 19010 16210 19022
rect 16158 18946 16210 18958
rect 17726 19010 17778 19022
rect 17726 18946 17778 18958
rect 17950 19010 18002 19022
rect 17950 18946 18002 18958
rect 18734 19010 18786 19022
rect 26126 19010 26178 19022
rect 20402 18958 20414 19010
rect 20466 18958 20478 19010
rect 18734 18946 18786 18958
rect 26126 18946 26178 18958
rect 26350 19010 26402 19022
rect 26350 18946 26402 18958
rect 35534 19010 35586 19022
rect 45726 19010 45778 19022
rect 47630 19010 47682 19022
rect 51102 19010 51154 19022
rect 41346 18958 41358 19010
rect 41410 18958 41422 19010
rect 45938 18958 45950 19010
rect 46002 18958 46014 19010
rect 49074 18958 49086 19010
rect 49138 18958 49150 19010
rect 35534 18946 35586 18958
rect 45726 18946 45778 18958
rect 47630 18946 47682 18958
rect 51102 18946 51154 18958
rect 1344 18842 58731 18876
rect 1344 18790 15520 18842
rect 15572 18790 15624 18842
rect 15676 18790 15728 18842
rect 15780 18790 29827 18842
rect 29879 18790 29931 18842
rect 29983 18790 30035 18842
rect 30087 18790 44134 18842
rect 44186 18790 44238 18842
rect 44290 18790 44342 18842
rect 44394 18790 58441 18842
rect 58493 18790 58545 18842
rect 58597 18790 58649 18842
rect 58701 18790 58731 18842
rect 1344 18756 58731 18790
rect 2046 18674 2098 18686
rect 3502 18674 3554 18686
rect 8654 18674 8706 18686
rect 3042 18622 3054 18674
rect 3106 18622 3118 18674
rect 4498 18622 4510 18674
rect 4562 18622 4574 18674
rect 2046 18610 2098 18622
rect 3502 18610 3554 18622
rect 8654 18610 8706 18622
rect 12126 18674 12178 18686
rect 12126 18610 12178 18622
rect 13694 18674 13746 18686
rect 13694 18610 13746 18622
rect 24446 18674 24498 18686
rect 24446 18610 24498 18622
rect 24670 18674 24722 18686
rect 33294 18674 33346 18686
rect 30034 18622 30046 18674
rect 30098 18622 30110 18674
rect 24670 18610 24722 18622
rect 33294 18610 33346 18622
rect 33966 18674 34018 18686
rect 33966 18610 34018 18622
rect 34190 18674 34242 18686
rect 34190 18610 34242 18622
rect 36318 18674 36370 18686
rect 36318 18610 36370 18622
rect 37774 18674 37826 18686
rect 37774 18610 37826 18622
rect 38782 18674 38834 18686
rect 42702 18674 42754 18686
rect 41458 18622 41470 18674
rect 41522 18622 41534 18674
rect 38782 18610 38834 18622
rect 42702 18610 42754 18622
rect 47854 18674 47906 18686
rect 47854 18610 47906 18622
rect 50542 18674 50594 18686
rect 50542 18610 50594 18622
rect 51102 18674 51154 18686
rect 51102 18610 51154 18622
rect 3390 18562 3442 18574
rect 5854 18562 5906 18574
rect 8542 18562 8594 18574
rect 3602 18510 3614 18562
rect 3666 18510 3678 18562
rect 5170 18510 5182 18562
rect 5234 18510 5246 18562
rect 6850 18510 6862 18562
rect 6914 18510 6926 18562
rect 3390 18498 3442 18510
rect 5854 18498 5906 18510
rect 8542 18498 8594 18510
rect 13022 18562 13074 18574
rect 13022 18498 13074 18510
rect 13470 18562 13522 18574
rect 21198 18562 21250 18574
rect 14690 18510 14702 18562
rect 14754 18510 14766 18562
rect 19730 18510 19742 18562
rect 19794 18510 19806 18562
rect 13470 18498 13522 18510
rect 21198 18498 21250 18510
rect 22766 18562 22818 18574
rect 22766 18498 22818 18510
rect 26686 18562 26738 18574
rect 26686 18498 26738 18510
rect 28590 18562 28642 18574
rect 28590 18498 28642 18510
rect 30942 18562 30994 18574
rect 30942 18498 30994 18510
rect 31054 18562 31106 18574
rect 31054 18498 31106 18510
rect 31502 18562 31554 18574
rect 31502 18498 31554 18510
rect 34862 18562 34914 18574
rect 34862 18498 34914 18510
rect 34974 18562 35026 18574
rect 34974 18498 35026 18510
rect 37886 18562 37938 18574
rect 49982 18562 50034 18574
rect 46498 18510 46510 18562
rect 46562 18510 46574 18562
rect 47170 18510 47182 18562
rect 47234 18510 47246 18562
rect 37886 18498 37938 18510
rect 49982 18498 50034 18510
rect 50430 18562 50482 18574
rect 51986 18510 51998 18562
rect 52050 18510 52062 18562
rect 50430 18498 50482 18510
rect 4846 18450 4898 18462
rect 1810 18398 1822 18450
rect 1874 18398 1886 18450
rect 2818 18398 2830 18450
rect 2882 18398 2894 18450
rect 4162 18398 4174 18450
rect 4226 18398 4238 18450
rect 4846 18386 4898 18398
rect 5518 18450 5570 18462
rect 5518 18386 5570 18398
rect 6190 18450 6242 18462
rect 6190 18386 6242 18398
rect 6526 18450 6578 18462
rect 6526 18386 6578 18398
rect 7646 18450 7698 18462
rect 7646 18386 7698 18398
rect 8206 18450 8258 18462
rect 10334 18450 10386 18462
rect 8866 18398 8878 18450
rect 8930 18398 8942 18450
rect 10210 18398 10222 18450
rect 10274 18398 10286 18450
rect 8206 18386 8258 18398
rect 10334 18386 10386 18398
rect 11230 18450 11282 18462
rect 11230 18386 11282 18398
rect 11678 18450 11730 18462
rect 11678 18386 11730 18398
rect 12686 18450 12738 18462
rect 12686 18386 12738 18398
rect 13358 18450 13410 18462
rect 17950 18450 18002 18462
rect 18846 18450 18898 18462
rect 21086 18450 21138 18462
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 18498 18398 18510 18450
rect 18562 18398 18574 18450
rect 19282 18398 19294 18450
rect 19346 18398 19358 18450
rect 20402 18398 20414 18450
rect 20466 18398 20478 18450
rect 13358 18386 13410 18398
rect 17950 18386 18002 18398
rect 18846 18386 18898 18398
rect 21086 18386 21138 18398
rect 21422 18450 21474 18462
rect 23102 18450 23154 18462
rect 22194 18398 22206 18450
rect 22258 18398 22270 18450
rect 21422 18386 21474 18398
rect 23102 18386 23154 18398
rect 23662 18450 23714 18462
rect 23662 18386 23714 18398
rect 24110 18450 24162 18462
rect 24110 18386 24162 18398
rect 24782 18450 24834 18462
rect 26126 18450 26178 18462
rect 25890 18398 25902 18450
rect 25954 18398 25966 18450
rect 24782 18386 24834 18398
rect 26126 18386 26178 18398
rect 26462 18450 26514 18462
rect 26462 18386 26514 18398
rect 26798 18450 26850 18462
rect 29150 18450 29202 18462
rect 27906 18398 27918 18450
rect 27970 18398 27982 18450
rect 28354 18398 28366 18450
rect 28418 18398 28430 18450
rect 26798 18386 26850 18398
rect 29150 18386 29202 18398
rect 29262 18450 29314 18462
rect 29262 18386 29314 18398
rect 29374 18450 29426 18462
rect 29374 18386 29426 18398
rect 29822 18450 29874 18462
rect 29822 18386 29874 18398
rect 31278 18450 31330 18462
rect 32398 18450 32450 18462
rect 32162 18398 32174 18450
rect 32226 18398 32238 18450
rect 31278 18386 31330 18398
rect 32398 18386 32450 18398
rect 33070 18450 33122 18462
rect 33070 18386 33122 18398
rect 33182 18450 33234 18462
rect 33854 18450 33906 18462
rect 34638 18450 34690 18462
rect 33618 18398 33630 18450
rect 33682 18398 33694 18450
rect 34402 18398 34414 18450
rect 34466 18398 34478 18450
rect 33182 18386 33234 18398
rect 33854 18386 33906 18398
rect 34638 18386 34690 18398
rect 36766 18450 36818 18462
rect 36766 18386 36818 18398
rect 37102 18450 37154 18462
rect 37102 18386 37154 18398
rect 37326 18450 37378 18462
rect 37326 18386 37378 18398
rect 37550 18450 37602 18462
rect 37550 18386 37602 18398
rect 40462 18450 40514 18462
rect 40462 18386 40514 18398
rect 41806 18450 41858 18462
rect 41806 18386 41858 18398
rect 42030 18450 42082 18462
rect 42030 18386 42082 18398
rect 42366 18450 42418 18462
rect 44382 18450 44434 18462
rect 43810 18398 43822 18450
rect 43874 18398 43886 18450
rect 42366 18386 42418 18398
rect 44382 18386 44434 18398
rect 44718 18450 44770 18462
rect 46846 18450 46898 18462
rect 46274 18398 46286 18450
rect 46338 18398 46350 18450
rect 44718 18386 44770 18398
rect 46846 18386 46898 18398
rect 47518 18450 47570 18462
rect 47518 18386 47570 18398
rect 48974 18450 49026 18462
rect 48974 18386 49026 18398
rect 49870 18450 49922 18462
rect 49870 18386 49922 18398
rect 50206 18450 50258 18462
rect 50206 18386 50258 18398
rect 50766 18450 50818 18462
rect 56030 18450 56082 18462
rect 52994 18398 53006 18450
rect 53058 18398 53070 18450
rect 55122 18398 55134 18450
rect 55186 18398 55198 18450
rect 57138 18398 57150 18450
rect 57202 18398 57214 18450
rect 50766 18386 50818 18398
rect 56030 18386 56082 18398
rect 7310 18338 7362 18350
rect 17614 18338 17666 18350
rect 25230 18338 25282 18350
rect 10658 18286 10670 18338
rect 10722 18286 10734 18338
rect 16818 18286 16830 18338
rect 16882 18286 16894 18338
rect 19618 18286 19630 18338
rect 19682 18286 19694 18338
rect 21970 18286 21982 18338
rect 22034 18286 22046 18338
rect 7310 18274 7362 18286
rect 17614 18274 17666 18286
rect 25230 18274 25282 18286
rect 30382 18338 30434 18350
rect 30382 18274 30434 18286
rect 30606 18338 30658 18350
rect 30606 18274 30658 18286
rect 35534 18338 35586 18350
rect 35534 18274 35586 18286
rect 35870 18338 35922 18350
rect 35870 18274 35922 18286
rect 37214 18338 37266 18350
rect 37214 18274 37266 18286
rect 38334 18338 38386 18350
rect 38334 18274 38386 18286
rect 41022 18338 41074 18350
rect 41022 18274 41074 18286
rect 44158 18338 44210 18350
rect 45726 18338 45778 18350
rect 45154 18286 45166 18338
rect 45218 18286 45230 18338
rect 44158 18274 44210 18286
rect 45726 18274 45778 18286
rect 49534 18338 49586 18350
rect 53678 18338 53730 18350
rect 51538 18286 51550 18338
rect 51602 18286 51614 18338
rect 55570 18286 55582 18338
rect 55634 18286 55646 18338
rect 56802 18286 56814 18338
rect 56866 18286 56878 18338
rect 49534 18274 49586 18286
rect 53678 18274 53730 18286
rect 11454 18226 11506 18238
rect 3938 18174 3950 18226
rect 4002 18174 4014 18226
rect 9762 18174 9774 18226
rect 9826 18174 9838 18226
rect 40786 18174 40798 18226
rect 40850 18223 40862 18226
rect 41010 18223 41022 18226
rect 40850 18177 41022 18223
rect 40850 18174 40862 18177
rect 41010 18174 41022 18177
rect 41074 18174 41086 18226
rect 56690 18174 56702 18226
rect 56754 18174 56766 18226
rect 11454 18162 11506 18174
rect 1344 18058 58576 18092
rect 1344 18006 8367 18058
rect 8419 18006 8471 18058
rect 8523 18006 8575 18058
rect 8627 18006 22674 18058
rect 22726 18006 22778 18058
rect 22830 18006 22882 18058
rect 22934 18006 36981 18058
rect 37033 18006 37085 18058
rect 37137 18006 37189 18058
rect 37241 18006 51288 18058
rect 51340 18006 51392 18058
rect 51444 18006 51496 18058
rect 51548 18006 58576 18058
rect 1344 17972 58576 18006
rect 10334 17890 10386 17902
rect 10334 17826 10386 17838
rect 10558 17890 10610 17902
rect 10558 17826 10610 17838
rect 16606 17890 16658 17902
rect 16606 17826 16658 17838
rect 30718 17890 30770 17902
rect 35310 17890 35362 17902
rect 34962 17838 34974 17890
rect 35026 17838 35038 17890
rect 30718 17826 30770 17838
rect 35310 17826 35362 17838
rect 35758 17890 35810 17902
rect 35758 17826 35810 17838
rect 50542 17890 50594 17902
rect 55582 17890 55634 17902
rect 53330 17838 53342 17890
rect 53394 17838 53406 17890
rect 50542 17826 50594 17838
rect 55582 17826 55634 17838
rect 55918 17890 55970 17902
rect 55918 17826 55970 17838
rect 4062 17778 4114 17790
rect 12910 17778 12962 17790
rect 17278 17778 17330 17790
rect 11890 17726 11902 17778
rect 11954 17726 11966 17778
rect 16146 17726 16158 17778
rect 16210 17726 16222 17778
rect 4062 17714 4114 17726
rect 12910 17714 12962 17726
rect 17278 17714 17330 17726
rect 18622 17778 18674 17790
rect 18622 17714 18674 17726
rect 20190 17778 20242 17790
rect 20190 17714 20242 17726
rect 28030 17778 28082 17790
rect 32286 17778 32338 17790
rect 30034 17726 30046 17778
rect 30098 17726 30110 17778
rect 28030 17714 28082 17726
rect 32286 17714 32338 17726
rect 33966 17778 34018 17790
rect 33966 17714 34018 17726
rect 37102 17778 37154 17790
rect 49310 17778 49362 17790
rect 40338 17726 40350 17778
rect 40402 17726 40414 17778
rect 41458 17726 41470 17778
rect 41522 17726 41534 17778
rect 43922 17726 43934 17778
rect 43986 17726 43998 17778
rect 37102 17714 37154 17726
rect 49310 17714 49362 17726
rect 51774 17778 51826 17790
rect 51774 17714 51826 17726
rect 55246 17778 55298 17790
rect 57822 17778 57874 17790
rect 56690 17726 56702 17778
rect 56754 17726 56766 17778
rect 55246 17714 55298 17726
rect 57822 17714 57874 17726
rect 1710 17666 1762 17678
rect 6414 17666 6466 17678
rect 2594 17614 2606 17666
rect 2658 17614 2670 17666
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 5842 17614 5854 17666
rect 5906 17614 5918 17666
rect 1710 17602 1762 17614
rect 6414 17602 6466 17614
rect 7086 17666 7138 17678
rect 8542 17666 8594 17678
rect 10110 17666 10162 17678
rect 12574 17666 12626 17678
rect 7522 17614 7534 17666
rect 7586 17614 7598 17666
rect 9650 17614 9662 17666
rect 9714 17614 9726 17666
rect 11778 17614 11790 17666
rect 11842 17614 11854 17666
rect 12114 17614 12126 17666
rect 12178 17614 12190 17666
rect 7086 17602 7138 17614
rect 8542 17602 8594 17614
rect 10110 17602 10162 17614
rect 12574 17602 12626 17614
rect 13470 17666 13522 17678
rect 13470 17602 13522 17614
rect 14030 17666 14082 17678
rect 14030 17602 14082 17614
rect 14478 17666 14530 17678
rect 14478 17602 14530 17614
rect 14926 17666 14978 17678
rect 14926 17602 14978 17614
rect 17726 17666 17778 17678
rect 19518 17666 19570 17678
rect 19282 17614 19294 17666
rect 19346 17614 19358 17666
rect 17726 17602 17778 17614
rect 19518 17602 19570 17614
rect 20526 17666 20578 17678
rect 20526 17602 20578 17614
rect 20862 17666 20914 17678
rect 27918 17666 27970 17678
rect 26562 17614 26574 17666
rect 26626 17614 26638 17666
rect 27346 17614 27358 17666
rect 27410 17614 27422 17666
rect 20862 17602 20914 17614
rect 27918 17602 27970 17614
rect 29150 17666 29202 17678
rect 31278 17666 31330 17678
rect 29586 17614 29598 17666
rect 29650 17614 29662 17666
rect 30818 17614 30830 17666
rect 30882 17614 30894 17666
rect 29150 17602 29202 17614
rect 31278 17602 31330 17614
rect 31614 17666 31666 17678
rect 33182 17666 33234 17678
rect 32722 17614 32734 17666
rect 32786 17614 32798 17666
rect 31614 17602 31666 17614
rect 33182 17602 33234 17614
rect 34750 17666 34802 17678
rect 34750 17602 34802 17614
rect 35534 17666 35586 17678
rect 45614 17666 45666 17678
rect 36306 17614 36318 17666
rect 36370 17614 36382 17666
rect 37538 17614 37550 17666
rect 37602 17614 37614 17666
rect 38210 17614 38222 17666
rect 38274 17614 38286 17666
rect 42914 17614 42926 17666
rect 42978 17614 42990 17666
rect 35534 17602 35586 17614
rect 45614 17602 45666 17614
rect 45950 17666 46002 17678
rect 45950 17602 46002 17614
rect 48750 17666 48802 17678
rect 48750 17602 48802 17614
rect 49534 17666 49586 17678
rect 49534 17602 49586 17614
rect 50766 17666 50818 17678
rect 50766 17602 50818 17614
rect 51102 17666 51154 17678
rect 54910 17666 54962 17678
rect 53106 17614 53118 17666
rect 53170 17614 53182 17666
rect 53330 17614 53342 17666
rect 53394 17614 53406 17666
rect 54450 17614 54462 17666
rect 54514 17614 54526 17666
rect 55570 17614 55582 17666
rect 55634 17614 55646 17666
rect 56914 17614 56926 17666
rect 56978 17614 56990 17666
rect 51102 17602 51154 17614
rect 54910 17602 54962 17614
rect 2046 17554 2098 17566
rect 2046 17490 2098 17502
rect 2382 17554 2434 17566
rect 2382 17490 2434 17502
rect 3950 17554 4002 17566
rect 3950 17490 4002 17502
rect 4958 17554 5010 17566
rect 13582 17554 13634 17566
rect 9426 17502 9438 17554
rect 9490 17502 9502 17554
rect 4958 17490 5010 17502
rect 13582 17490 13634 17502
rect 14702 17554 14754 17566
rect 14702 17490 14754 17502
rect 15150 17554 15202 17566
rect 15150 17490 15202 17502
rect 15262 17554 15314 17566
rect 15262 17490 15314 17502
rect 15822 17554 15874 17566
rect 15822 17490 15874 17502
rect 16046 17554 16098 17566
rect 16046 17490 16098 17502
rect 16494 17554 16546 17566
rect 16494 17490 16546 17502
rect 16606 17554 16658 17566
rect 16606 17490 16658 17502
rect 20638 17554 20690 17566
rect 30606 17554 30658 17566
rect 21522 17502 21534 17554
rect 21586 17502 21598 17554
rect 20638 17490 20690 17502
rect 30606 17490 30658 17502
rect 34190 17554 34242 17566
rect 46510 17554 46562 17566
rect 49086 17554 49138 17566
rect 42018 17502 42030 17554
rect 42082 17502 42094 17554
rect 44818 17502 44830 17554
rect 44882 17502 44894 17554
rect 47842 17502 47854 17554
rect 47906 17502 47918 17554
rect 34190 17490 34242 17502
rect 46510 17490 46562 17502
rect 49086 17490 49138 17502
rect 54686 17554 54738 17566
rect 54686 17490 54738 17502
rect 56254 17554 56306 17566
rect 56254 17490 56306 17502
rect 57710 17554 57762 17566
rect 57710 17490 57762 17502
rect 3166 17442 3218 17454
rect 3166 17378 3218 17390
rect 3726 17442 3778 17454
rect 3726 17378 3778 17390
rect 4622 17442 4674 17454
rect 9102 17442 9154 17454
rect 5618 17390 5630 17442
rect 5682 17390 5694 17442
rect 7746 17390 7758 17442
rect 7810 17390 7822 17442
rect 4622 17378 4674 17390
rect 9102 17378 9154 17390
rect 11006 17442 11058 17454
rect 11006 17378 11058 17390
rect 13806 17442 13858 17454
rect 13806 17378 13858 17390
rect 14366 17442 14418 17454
rect 14366 17378 14418 17390
rect 17838 17442 17890 17454
rect 17838 17378 17890 17390
rect 18062 17442 18114 17454
rect 18062 17378 18114 17390
rect 31054 17442 31106 17454
rect 31054 17378 31106 17390
rect 31502 17442 31554 17454
rect 31502 17378 31554 17390
rect 34414 17442 34466 17454
rect 34414 17378 34466 17390
rect 34638 17442 34690 17454
rect 34638 17378 34690 17390
rect 35870 17442 35922 17454
rect 35870 17378 35922 17390
rect 36094 17442 36146 17454
rect 36094 17378 36146 17390
rect 45166 17442 45218 17454
rect 45166 17378 45218 17390
rect 45726 17442 45778 17454
rect 45726 17378 45778 17390
rect 46846 17442 46898 17454
rect 46846 17378 46898 17390
rect 47518 17442 47570 17454
rect 47518 17378 47570 17390
rect 48414 17442 48466 17454
rect 48414 17378 48466 17390
rect 48862 17442 48914 17454
rect 51214 17442 51266 17454
rect 49858 17390 49870 17442
rect 49922 17390 49934 17442
rect 50194 17390 50206 17442
rect 50258 17390 50270 17442
rect 48862 17378 48914 17390
rect 51214 17378 51266 17390
rect 51438 17442 51490 17454
rect 51438 17378 51490 17390
rect 57934 17442 57986 17454
rect 57934 17378 57986 17390
rect 1344 17274 58731 17308
rect 1344 17222 15520 17274
rect 15572 17222 15624 17274
rect 15676 17222 15728 17274
rect 15780 17222 29827 17274
rect 29879 17222 29931 17274
rect 29983 17222 30035 17274
rect 30087 17222 44134 17274
rect 44186 17222 44238 17274
rect 44290 17222 44342 17274
rect 44394 17222 58441 17274
rect 58493 17222 58545 17274
rect 58597 17222 58649 17274
rect 58701 17222 58731 17274
rect 1344 17188 58731 17222
rect 2046 17106 2098 17118
rect 2046 17042 2098 17054
rect 6414 17106 6466 17118
rect 6414 17042 6466 17054
rect 11454 17106 11506 17118
rect 11454 17042 11506 17054
rect 12798 17106 12850 17118
rect 12798 17042 12850 17054
rect 13022 17106 13074 17118
rect 13022 17042 13074 17054
rect 13358 17106 13410 17118
rect 13358 17042 13410 17054
rect 14030 17106 14082 17118
rect 20862 17106 20914 17118
rect 14354 17054 14366 17106
rect 14418 17054 14430 17106
rect 14030 17042 14082 17054
rect 20862 17042 20914 17054
rect 24222 17106 24274 17118
rect 24222 17042 24274 17054
rect 24446 17106 24498 17118
rect 24446 17042 24498 17054
rect 30270 17106 30322 17118
rect 30270 17042 30322 17054
rect 31390 17106 31442 17118
rect 33630 17106 33682 17118
rect 35086 17106 35138 17118
rect 32162 17054 32174 17106
rect 32226 17054 32238 17106
rect 33058 17054 33070 17106
rect 33122 17054 33134 17106
rect 34738 17054 34750 17106
rect 34802 17054 34814 17106
rect 31390 17042 31442 17054
rect 33630 17042 33682 17054
rect 35086 17042 35138 17054
rect 35646 17106 35698 17118
rect 35646 17042 35698 17054
rect 42366 17106 42418 17118
rect 42366 17042 42418 17054
rect 43150 17106 43202 17118
rect 43150 17042 43202 17054
rect 45278 17106 45330 17118
rect 47742 17106 47794 17118
rect 45938 17054 45950 17106
rect 46002 17054 46014 17106
rect 45278 17042 45330 17054
rect 47742 17042 47794 17054
rect 50430 17106 50482 17118
rect 50430 17042 50482 17054
rect 55918 17106 55970 17118
rect 55918 17042 55970 17054
rect 2382 16994 2434 17006
rect 2382 16930 2434 16942
rect 2718 16994 2770 17006
rect 8318 16994 8370 17006
rect 3826 16942 3838 16994
rect 3890 16942 3902 16994
rect 2718 16930 2770 16942
rect 8318 16930 8370 16942
rect 9550 16994 9602 17006
rect 9550 16930 9602 16942
rect 10894 16994 10946 17006
rect 10894 16930 10946 16942
rect 12686 16994 12738 17006
rect 12686 16930 12738 16942
rect 15262 16994 15314 17006
rect 15262 16930 15314 16942
rect 15710 16994 15762 17006
rect 15710 16930 15762 16942
rect 16830 16994 16882 17006
rect 20974 16994 21026 17006
rect 18162 16942 18174 16994
rect 18226 16942 18238 16994
rect 16830 16930 16882 16942
rect 20974 16930 21026 16942
rect 21310 16994 21362 17006
rect 21310 16930 21362 16942
rect 29038 16994 29090 17006
rect 29038 16930 29090 16942
rect 30494 16994 30546 17006
rect 30494 16930 30546 16942
rect 30606 16994 30658 17006
rect 30606 16930 30658 16942
rect 31726 16994 31778 17006
rect 31726 16930 31778 16942
rect 33406 16994 33458 17006
rect 33406 16930 33458 16942
rect 33854 16994 33906 17006
rect 33854 16930 33906 16942
rect 35982 16994 36034 17006
rect 35982 16930 36034 16942
rect 41246 16994 41298 17006
rect 41246 16930 41298 16942
rect 43038 16994 43090 17006
rect 43038 16930 43090 16942
rect 43598 16994 43650 17006
rect 43598 16930 43650 16942
rect 43934 16994 43986 17006
rect 46958 16994 47010 17006
rect 45602 16942 45614 16994
rect 45666 16942 45678 16994
rect 43934 16930 43986 16942
rect 46958 16930 47010 16942
rect 47294 16994 47346 17006
rect 47294 16930 47346 16942
rect 1710 16882 1762 16894
rect 12014 16882 12066 16894
rect 3042 16830 3054 16882
rect 3106 16830 3118 16882
rect 7746 16830 7758 16882
rect 7810 16830 7822 16882
rect 8530 16830 8542 16882
rect 8594 16830 8606 16882
rect 8754 16830 8766 16882
rect 8818 16830 8830 16882
rect 1710 16818 1762 16830
rect 12014 16818 12066 16830
rect 13470 16882 13522 16894
rect 13470 16818 13522 16830
rect 14702 16882 14754 16894
rect 14702 16818 14754 16830
rect 15038 16882 15090 16894
rect 20638 16882 20690 16894
rect 22206 16882 22258 16894
rect 16258 16830 16270 16882
rect 16322 16830 16334 16882
rect 16594 16830 16606 16882
rect 16658 16830 16670 16882
rect 17490 16830 17502 16882
rect 17554 16830 17566 16882
rect 21746 16830 21758 16882
rect 21810 16830 21822 16882
rect 15038 16818 15090 16830
rect 20638 16818 20690 16830
rect 22206 16818 22258 16830
rect 22654 16882 22706 16894
rect 24782 16882 24834 16894
rect 33966 16882 34018 16894
rect 23090 16830 23102 16882
rect 23154 16830 23166 16882
rect 25666 16830 25678 16882
rect 25730 16830 25742 16882
rect 27346 16830 27358 16882
rect 27410 16830 27422 16882
rect 28354 16830 28366 16882
rect 28418 16830 28430 16882
rect 29474 16830 29486 16882
rect 29538 16830 29550 16882
rect 32386 16830 32398 16882
rect 32450 16830 32462 16882
rect 22654 16818 22706 16830
rect 24782 16818 24834 16830
rect 33966 16818 34018 16830
rect 34414 16882 34466 16894
rect 34414 16818 34466 16830
rect 35870 16882 35922 16894
rect 35870 16818 35922 16830
rect 36206 16882 36258 16894
rect 36206 16818 36258 16830
rect 36430 16882 36482 16894
rect 36430 16818 36482 16830
rect 36654 16882 36706 16894
rect 36654 16818 36706 16830
rect 36878 16882 36930 16894
rect 36878 16818 36930 16830
rect 37102 16882 37154 16894
rect 41134 16882 41186 16894
rect 37426 16830 37438 16882
rect 37490 16830 37502 16882
rect 38098 16830 38110 16882
rect 38162 16830 38174 16882
rect 37102 16818 37154 16830
rect 41134 16818 41186 16830
rect 41470 16882 41522 16894
rect 41470 16818 41522 16830
rect 42702 16882 42754 16894
rect 42702 16818 42754 16830
rect 43374 16882 43426 16894
rect 47630 16882 47682 16894
rect 46162 16830 46174 16882
rect 46226 16830 46238 16882
rect 43374 16818 43426 16830
rect 47630 16818 47682 16830
rect 48974 16882 49026 16894
rect 48974 16818 49026 16830
rect 49198 16882 49250 16894
rect 49198 16818 49250 16830
rect 49646 16882 49698 16894
rect 55134 16882 55186 16894
rect 51202 16830 51214 16882
rect 51266 16830 51278 16882
rect 52770 16830 52782 16882
rect 52834 16830 52846 16882
rect 54674 16830 54686 16882
rect 54738 16830 54750 16882
rect 49646 16818 49698 16830
rect 55134 16818 55186 16830
rect 56814 16882 56866 16894
rect 57138 16830 57150 16882
rect 57202 16830 57214 16882
rect 56814 16818 56866 16830
rect 6974 16770 7026 16782
rect 9774 16770 9826 16782
rect 5954 16718 5966 16770
rect 6018 16718 6030 16770
rect 7634 16718 7646 16770
rect 7698 16718 7710 16770
rect 6974 16706 7026 16718
rect 9774 16706 9826 16718
rect 11006 16770 11058 16782
rect 11006 16706 11058 16718
rect 11118 16770 11170 16782
rect 11118 16706 11170 16718
rect 15150 16770 15202 16782
rect 15150 16706 15202 16718
rect 16718 16770 16770 16782
rect 24558 16770 24610 16782
rect 20290 16718 20302 16770
rect 20354 16718 20366 16770
rect 23426 16718 23438 16770
rect 23490 16718 23502 16770
rect 16718 16706 16770 16718
rect 24558 16706 24610 16718
rect 25342 16770 25394 16782
rect 49086 16770 49138 16782
rect 25554 16718 25566 16770
rect 25618 16718 25630 16770
rect 27794 16718 27806 16770
rect 27858 16718 27870 16770
rect 29922 16718 29934 16770
rect 29986 16718 29998 16770
rect 40226 16718 40238 16770
rect 40290 16718 40302 16770
rect 25342 16706 25394 16718
rect 49086 16706 49138 16718
rect 49982 16770 50034 16782
rect 51886 16770 51938 16782
rect 53566 16770 53618 16782
rect 55694 16770 55746 16782
rect 51426 16718 51438 16770
rect 51490 16718 51502 16770
rect 53106 16718 53118 16770
rect 53170 16718 53182 16770
rect 54338 16718 54350 16770
rect 54402 16718 54414 16770
rect 56018 16718 56030 16770
rect 56082 16718 56094 16770
rect 49982 16706 50034 16718
rect 51886 16706 51938 16718
rect 53566 16706 53618 16718
rect 55694 16706 55746 16718
rect 8206 16658 8258 16670
rect 8206 16594 8258 16606
rect 10110 16658 10162 16670
rect 10110 16594 10162 16606
rect 13358 16658 13410 16670
rect 47742 16658 47794 16670
rect 16258 16606 16270 16658
rect 16322 16606 16334 16658
rect 27346 16606 27358 16658
rect 27410 16606 27422 16658
rect 56914 16606 56926 16658
rect 56978 16606 56990 16658
rect 13358 16594 13410 16606
rect 47742 16594 47794 16606
rect 1344 16490 58576 16524
rect 1344 16438 8367 16490
rect 8419 16438 8471 16490
rect 8523 16438 8575 16490
rect 8627 16438 22674 16490
rect 22726 16438 22778 16490
rect 22830 16438 22882 16490
rect 22934 16438 36981 16490
rect 37033 16438 37085 16490
rect 37137 16438 37189 16490
rect 37241 16438 51288 16490
rect 51340 16438 51392 16490
rect 51444 16438 51496 16490
rect 51548 16438 58576 16490
rect 1344 16404 58576 16438
rect 12686 16322 12738 16334
rect 28366 16322 28418 16334
rect 49870 16322 49922 16334
rect 55582 16322 55634 16334
rect 24770 16270 24782 16322
rect 24834 16270 24846 16322
rect 27346 16270 27358 16322
rect 27410 16270 27422 16322
rect 42354 16270 42366 16322
rect 42418 16270 42430 16322
rect 48962 16270 48974 16322
rect 49026 16270 49038 16322
rect 50978 16270 50990 16322
rect 51042 16319 51054 16322
rect 51314 16319 51326 16322
rect 51042 16273 51326 16319
rect 51042 16270 51054 16273
rect 51314 16270 51326 16273
rect 51378 16270 51390 16322
rect 12686 16258 12738 16270
rect 28366 16258 28418 16270
rect 49870 16258 49922 16270
rect 55582 16258 55634 16270
rect 9774 16210 9826 16222
rect 2482 16158 2494 16210
rect 2546 16158 2558 16210
rect 4610 16158 4622 16210
rect 4674 16158 4686 16210
rect 6962 16158 6974 16210
rect 7026 16158 7038 16210
rect 9774 16146 9826 16158
rect 14366 16210 14418 16222
rect 19630 16210 19682 16222
rect 29374 16210 29426 16222
rect 15586 16158 15598 16210
rect 15650 16158 15662 16210
rect 17714 16158 17726 16210
rect 17778 16158 17790 16210
rect 21746 16158 21758 16210
rect 21810 16158 21822 16210
rect 25106 16158 25118 16210
rect 25170 16158 25182 16210
rect 27570 16158 27582 16210
rect 27634 16158 27646 16210
rect 14366 16146 14418 16158
rect 19630 16146 19682 16158
rect 29374 16146 29426 16158
rect 31278 16210 31330 16222
rect 31278 16146 31330 16158
rect 34414 16210 34466 16222
rect 34414 16146 34466 16158
rect 34974 16210 35026 16222
rect 34974 16146 35026 16158
rect 35310 16210 35362 16222
rect 35310 16146 35362 16158
rect 38110 16210 38162 16222
rect 38110 16146 38162 16158
rect 38894 16210 38946 16222
rect 44158 16210 44210 16222
rect 42466 16158 42478 16210
rect 42530 16158 42542 16210
rect 43250 16158 43262 16210
rect 43314 16158 43326 16210
rect 38894 16146 38946 16158
rect 44158 16146 44210 16158
rect 48414 16210 48466 16222
rect 48414 16146 48466 16158
rect 49310 16210 49362 16222
rect 49310 16146 49362 16158
rect 50878 16210 50930 16222
rect 50878 16146 50930 16158
rect 51326 16210 51378 16222
rect 51326 16146 51378 16158
rect 51774 16210 51826 16222
rect 52994 16158 53006 16210
rect 53058 16158 53070 16210
rect 56018 16158 56030 16210
rect 56082 16158 56094 16210
rect 51774 16146 51826 16158
rect 6302 16098 6354 16110
rect 8542 16098 8594 16110
rect 1810 16046 1822 16098
rect 1874 16046 1886 16098
rect 7186 16046 7198 16098
rect 7250 16046 7262 16098
rect 6302 16034 6354 16046
rect 8542 16034 8594 16046
rect 8990 16098 9042 16110
rect 11342 16098 11394 16110
rect 12574 16098 12626 16110
rect 18286 16098 18338 16110
rect 10770 16046 10782 16098
rect 10834 16046 10846 16098
rect 12002 16046 12014 16098
rect 12066 16046 12078 16098
rect 14914 16046 14926 16098
rect 14978 16046 14990 16098
rect 8990 16034 9042 16046
rect 11342 16034 11394 16046
rect 12574 16034 12626 16046
rect 18286 16034 18338 16046
rect 20526 16098 20578 16110
rect 20526 16034 20578 16046
rect 20862 16098 20914 16110
rect 28254 16098 28306 16110
rect 23314 16046 23326 16098
rect 23378 16046 23390 16098
rect 25330 16046 25342 16098
rect 25394 16046 25406 16098
rect 27682 16046 27694 16098
rect 27746 16046 27758 16098
rect 20862 16034 20914 16046
rect 28254 16034 28306 16046
rect 29710 16098 29762 16110
rect 29710 16034 29762 16046
rect 30046 16098 30098 16110
rect 30046 16034 30098 16046
rect 30382 16098 30434 16110
rect 32286 16098 32338 16110
rect 36206 16098 36258 16110
rect 30818 16046 30830 16098
rect 30882 16046 30894 16098
rect 33170 16046 33182 16098
rect 33234 16046 33246 16098
rect 30382 16034 30434 16046
rect 32286 16034 32338 16046
rect 36206 16034 36258 16046
rect 36990 16098 37042 16110
rect 36990 16034 37042 16046
rect 37662 16098 37714 16110
rect 37662 16034 37714 16046
rect 39902 16098 39954 16110
rect 39902 16034 39954 16046
rect 40462 16098 40514 16110
rect 45278 16098 45330 16110
rect 46174 16098 46226 16110
rect 42242 16046 42254 16098
rect 42306 16046 42318 16098
rect 43474 16046 43486 16098
rect 43538 16046 43550 16098
rect 45714 16046 45726 16098
rect 45778 16046 45790 16098
rect 40462 16034 40514 16046
rect 45278 16034 45330 16046
rect 46174 16034 46226 16046
rect 46510 16098 46562 16110
rect 46510 16034 46562 16046
rect 47070 16098 47122 16110
rect 47070 16034 47122 16046
rect 47854 16098 47906 16110
rect 47854 16034 47906 16046
rect 48190 16098 48242 16110
rect 48190 16034 48242 16046
rect 48638 16098 48690 16110
rect 48638 16034 48690 16046
rect 49534 16098 49586 16110
rect 49534 16034 49586 16046
rect 50094 16098 50146 16110
rect 55570 16046 55582 16098
rect 55634 16046 55646 16098
rect 50094 16034 50146 16046
rect 5070 15986 5122 15998
rect 5070 15922 5122 15934
rect 8094 15986 8146 15998
rect 8094 15922 8146 15934
rect 8766 15986 8818 15998
rect 8766 15922 8818 15934
rect 9214 15986 9266 15998
rect 9214 15922 9266 15934
rect 9326 15986 9378 15998
rect 9326 15922 9378 15934
rect 10558 15986 10610 15998
rect 10558 15922 10610 15934
rect 12238 15986 12290 15998
rect 12238 15922 12290 15934
rect 12686 15986 12738 15998
rect 12686 15922 12738 15934
rect 18398 15986 18450 15998
rect 26014 15986 26066 15998
rect 22194 15934 22206 15986
rect 22258 15934 22270 15986
rect 18398 15922 18450 15934
rect 26014 15922 26066 15934
rect 31726 15986 31778 15998
rect 31726 15922 31778 15934
rect 32062 15986 32114 15998
rect 32062 15922 32114 15934
rect 32622 15986 32674 15998
rect 32622 15922 32674 15934
rect 36542 15986 36594 15998
rect 36542 15922 36594 15934
rect 37214 15986 37266 15998
rect 46286 15986 46338 15998
rect 39554 15934 39566 15986
rect 39618 15934 39630 15986
rect 41010 15934 41022 15986
rect 41074 15934 41086 15986
rect 45490 15934 45502 15986
rect 45554 15934 45566 15986
rect 37214 15922 37266 15934
rect 46286 15922 46338 15934
rect 46734 15986 46786 15998
rect 46734 15922 46786 15934
rect 46846 15986 46898 15998
rect 46846 15922 46898 15934
rect 47966 15986 48018 15998
rect 47966 15922 48018 15934
rect 50318 15986 50370 15998
rect 50318 15922 50370 15934
rect 50430 15986 50482 15998
rect 50430 15922 50482 15934
rect 52670 15986 52722 15998
rect 52670 15922 52722 15934
rect 52894 15986 52946 15998
rect 52894 15922 52946 15934
rect 55246 15986 55298 15998
rect 56242 15934 56254 15986
rect 56306 15934 56318 15986
rect 57922 15934 57934 15986
rect 57986 15934 57998 15986
rect 55246 15922 55298 15934
rect 6078 15874 6130 15886
rect 6078 15810 6130 15822
rect 8318 15874 8370 15886
rect 8318 15810 8370 15822
rect 8878 15874 8930 15886
rect 8878 15810 8930 15822
rect 10222 15874 10274 15886
rect 10222 15810 10274 15822
rect 11454 15874 11506 15886
rect 11454 15810 11506 15822
rect 11678 15874 11730 15886
rect 11678 15810 11730 15822
rect 13918 15874 13970 15886
rect 13918 15810 13970 15822
rect 18622 15874 18674 15886
rect 18622 15810 18674 15822
rect 18958 15874 19010 15886
rect 18958 15810 19010 15822
rect 20078 15874 20130 15886
rect 20078 15810 20130 15822
rect 20638 15874 20690 15886
rect 26126 15874 26178 15886
rect 23538 15822 23550 15874
rect 23602 15822 23614 15874
rect 20638 15810 20690 15822
rect 26126 15810 26178 15822
rect 26350 15874 26402 15886
rect 26350 15810 26402 15822
rect 28366 15874 28418 15886
rect 28366 15810 28418 15822
rect 29822 15874 29874 15886
rect 29822 15810 29874 15822
rect 31950 15874 32002 15886
rect 31950 15810 32002 15822
rect 32510 15874 32562 15886
rect 33630 15874 33682 15886
rect 35758 15874 35810 15886
rect 32946 15822 32958 15874
rect 33010 15822 33022 15874
rect 33954 15822 33966 15874
rect 34018 15822 34030 15874
rect 32510 15810 32562 15822
rect 33630 15810 33682 15822
rect 35758 15810 35810 15822
rect 36318 15874 36370 15886
rect 36318 15810 36370 15822
rect 37438 15874 37490 15886
rect 37438 15810 37490 15822
rect 38446 15874 38498 15886
rect 38446 15810 38498 15822
rect 41358 15874 41410 15886
rect 41358 15810 41410 15822
rect 47406 15874 47458 15886
rect 57810 15822 57822 15874
rect 57874 15822 57886 15874
rect 47406 15810 47458 15822
rect 1344 15706 58731 15740
rect 1344 15654 15520 15706
rect 15572 15654 15624 15706
rect 15676 15654 15728 15706
rect 15780 15654 29827 15706
rect 29879 15654 29931 15706
rect 29983 15654 30035 15706
rect 30087 15654 44134 15706
rect 44186 15654 44238 15706
rect 44290 15654 44342 15706
rect 44394 15654 58441 15706
rect 58493 15654 58545 15706
rect 58597 15654 58649 15706
rect 58701 15654 58731 15706
rect 1344 15620 58731 15654
rect 5742 15538 5794 15550
rect 5742 15474 5794 15486
rect 11454 15538 11506 15550
rect 11454 15474 11506 15486
rect 15486 15538 15538 15550
rect 15486 15474 15538 15486
rect 15934 15538 15986 15550
rect 15934 15474 15986 15486
rect 16382 15538 16434 15550
rect 16382 15474 16434 15486
rect 17614 15538 17666 15550
rect 17614 15474 17666 15486
rect 18062 15538 18114 15550
rect 18062 15474 18114 15486
rect 20414 15538 20466 15550
rect 20414 15474 20466 15486
rect 21982 15538 22034 15550
rect 21982 15474 22034 15486
rect 22206 15538 22258 15550
rect 22206 15474 22258 15486
rect 25342 15538 25394 15550
rect 25342 15474 25394 15486
rect 28702 15538 28754 15550
rect 28702 15474 28754 15486
rect 28926 15538 28978 15550
rect 28926 15474 28978 15486
rect 30718 15538 30770 15550
rect 30718 15474 30770 15486
rect 33742 15538 33794 15550
rect 33742 15474 33794 15486
rect 41022 15538 41074 15550
rect 41022 15474 41074 15486
rect 42366 15538 42418 15550
rect 42366 15474 42418 15486
rect 43150 15538 43202 15550
rect 43150 15474 43202 15486
rect 43710 15538 43762 15550
rect 43710 15474 43762 15486
rect 44606 15538 44658 15550
rect 44606 15474 44658 15486
rect 47406 15538 47458 15550
rect 47406 15474 47458 15486
rect 48078 15538 48130 15550
rect 48078 15474 48130 15486
rect 56926 15538 56978 15550
rect 56926 15474 56978 15486
rect 57486 15538 57538 15550
rect 57486 15474 57538 15486
rect 5518 15426 5570 15438
rect 5518 15362 5570 15374
rect 6526 15426 6578 15438
rect 9886 15426 9938 15438
rect 7410 15374 7422 15426
rect 7474 15374 7486 15426
rect 6526 15362 6578 15374
rect 9886 15362 9938 15374
rect 10558 15426 10610 15438
rect 10558 15362 10610 15374
rect 20750 15426 20802 15438
rect 20750 15362 20802 15374
rect 22318 15426 22370 15438
rect 22318 15362 22370 15374
rect 23662 15426 23714 15438
rect 23662 15362 23714 15374
rect 26910 15426 26962 15438
rect 26910 15362 26962 15374
rect 27246 15426 27298 15438
rect 27246 15362 27298 15374
rect 27358 15426 27410 15438
rect 27358 15362 27410 15374
rect 27582 15426 27634 15438
rect 27582 15362 27634 15374
rect 28030 15426 28082 15438
rect 28030 15362 28082 15374
rect 30270 15426 30322 15438
rect 30270 15362 30322 15374
rect 35310 15426 35362 15438
rect 35310 15362 35362 15374
rect 35982 15426 36034 15438
rect 35982 15362 36034 15374
rect 36318 15426 36370 15438
rect 40910 15426 40962 15438
rect 37426 15374 37438 15426
rect 37490 15374 37502 15426
rect 36318 15362 36370 15374
rect 40910 15362 40962 15374
rect 41470 15426 41522 15438
rect 42926 15426 42978 15438
rect 41794 15374 41806 15426
rect 41858 15374 41870 15426
rect 41470 15362 41522 15374
rect 42926 15362 42978 15374
rect 43822 15426 43874 15438
rect 43822 15362 43874 15374
rect 44270 15426 44322 15438
rect 44270 15362 44322 15374
rect 48190 15426 48242 15438
rect 52446 15426 52498 15438
rect 49186 15374 49198 15426
rect 49250 15374 49262 15426
rect 50642 15374 50654 15426
rect 50706 15374 50718 15426
rect 48190 15362 48242 15374
rect 52446 15362 52498 15374
rect 55806 15426 55858 15438
rect 55806 15362 55858 15374
rect 56030 15426 56082 15438
rect 56030 15362 56082 15374
rect 56702 15426 56754 15438
rect 56702 15362 56754 15374
rect 57710 15426 57762 15438
rect 57710 15362 57762 15374
rect 15038 15314 15090 15326
rect 23102 15314 23154 15326
rect 1810 15262 1822 15314
rect 1874 15262 1886 15314
rect 5954 15262 5966 15314
rect 6018 15262 6030 15314
rect 6738 15262 6750 15314
rect 6802 15262 6814 15314
rect 7858 15262 7870 15314
rect 7922 15262 7934 15314
rect 10098 15262 10110 15314
rect 10162 15262 10174 15314
rect 10770 15262 10782 15314
rect 10834 15262 10846 15314
rect 14578 15262 14590 15314
rect 14642 15262 14654 15314
rect 21410 15262 21422 15314
rect 21474 15262 21486 15314
rect 22754 15262 22766 15314
rect 22818 15262 22830 15314
rect 15038 15250 15090 15262
rect 23102 15250 23154 15262
rect 23214 15314 23266 15326
rect 23214 15250 23266 15262
rect 23326 15314 23378 15326
rect 24558 15314 24610 15326
rect 24098 15262 24110 15314
rect 24162 15262 24174 15314
rect 23326 15250 23378 15262
rect 24558 15250 24610 15262
rect 25454 15314 25506 15326
rect 25454 15250 25506 15262
rect 26014 15314 26066 15326
rect 27918 15314 27970 15326
rect 26450 15262 26462 15314
rect 26514 15262 26526 15314
rect 26014 15250 26066 15262
rect 27918 15250 27970 15262
rect 28254 15314 28306 15326
rect 29374 15314 29426 15326
rect 32286 15314 32338 15326
rect 28466 15262 28478 15314
rect 28530 15262 28542 15314
rect 29586 15262 29598 15314
rect 29650 15262 29662 15314
rect 28254 15250 28306 15262
rect 29374 15250 29426 15262
rect 32286 15250 32338 15262
rect 33630 15314 33682 15326
rect 41246 15314 41298 15326
rect 34402 15262 34414 15314
rect 34466 15262 34478 15314
rect 36754 15262 36766 15314
rect 36818 15262 36830 15314
rect 33630 15250 33682 15262
rect 41246 15250 41298 15262
rect 42142 15314 42194 15326
rect 42142 15250 42194 15262
rect 44942 15314 44994 15326
rect 44942 15250 44994 15262
rect 45166 15314 45218 15326
rect 45166 15250 45218 15262
rect 46062 15314 46114 15326
rect 46062 15250 46114 15262
rect 46398 15314 46450 15326
rect 46398 15250 46450 15262
rect 46622 15314 46674 15326
rect 51538 15262 51550 15314
rect 51602 15262 51614 15314
rect 52994 15262 53006 15314
rect 53058 15262 53070 15314
rect 54786 15262 54798 15314
rect 54850 15262 54862 15314
rect 46622 15250 46674 15262
rect 5182 15202 5234 15214
rect 8990 15202 9042 15214
rect 16830 15202 16882 15214
rect 2482 15150 2494 15202
rect 2546 15150 2558 15202
rect 4610 15150 4622 15202
rect 4674 15150 4686 15202
rect 7970 15150 7982 15202
rect 8034 15150 8046 15202
rect 13794 15150 13806 15202
rect 13858 15150 13870 15202
rect 5182 15138 5234 15150
rect 8990 15138 9042 15150
rect 5854 15090 5906 15102
rect 11666 15094 11678 15146
rect 11730 15094 11742 15146
rect 16830 15138 16882 15150
rect 19070 15202 19122 15214
rect 43598 15202 43650 15214
rect 50990 15202 51042 15214
rect 57598 15202 57650 15214
rect 21522 15150 21534 15202
rect 21586 15150 21598 15202
rect 34514 15150 34526 15202
rect 34578 15150 34590 15202
rect 39554 15150 39566 15202
rect 39618 15150 39630 15202
rect 43250 15150 43262 15202
rect 43314 15150 43326 15202
rect 48850 15150 48862 15202
rect 48914 15150 48926 15202
rect 51650 15150 51662 15202
rect 51714 15150 51726 15202
rect 53218 15150 53230 15202
rect 53282 15150 53294 15202
rect 55122 15150 55134 15202
rect 55186 15150 55198 15202
rect 55682 15150 55694 15202
rect 55746 15150 55758 15202
rect 57026 15150 57038 15202
rect 57090 15150 57102 15202
rect 19070 15138 19122 15150
rect 43598 15138 43650 15150
rect 50990 15138 51042 15150
rect 57598 15138 57650 15150
rect 25342 15090 25394 15102
rect 14802 15038 14814 15090
rect 14866 15087 14878 15090
rect 15586 15087 15598 15090
rect 14866 15041 15598 15087
rect 14866 15038 14878 15041
rect 15586 15038 15598 15041
rect 15650 15038 15662 15090
rect 5854 15026 5906 15038
rect 25342 15026 25394 15038
rect 28590 15090 28642 15102
rect 28590 15026 28642 15038
rect 33742 15090 33794 15102
rect 33742 15026 33794 15038
rect 42478 15090 42530 15102
rect 48078 15090 48130 15102
rect 45490 15038 45502 15090
rect 45554 15038 45566 15090
rect 46946 15038 46958 15090
rect 47010 15038 47022 15090
rect 53778 15038 53790 15090
rect 53842 15038 53854 15090
rect 54674 15038 54686 15090
rect 54738 15038 54750 15090
rect 42478 15026 42530 15038
rect 48078 15026 48130 15038
rect 1344 14922 58576 14956
rect 1344 14870 8367 14922
rect 8419 14870 8471 14922
rect 8523 14870 8575 14922
rect 8627 14870 22674 14922
rect 22726 14870 22778 14922
rect 22830 14870 22882 14922
rect 22934 14870 36981 14922
rect 37033 14870 37085 14922
rect 37137 14870 37189 14922
rect 37241 14870 51288 14922
rect 51340 14870 51392 14922
rect 51444 14870 51496 14922
rect 51548 14870 58576 14922
rect 1344 14836 58576 14870
rect 4174 14754 4226 14766
rect 4174 14690 4226 14702
rect 4510 14754 4562 14766
rect 28366 14754 28418 14766
rect 6850 14702 6862 14754
rect 6914 14751 6926 14754
rect 7298 14751 7310 14754
rect 6914 14705 7310 14751
rect 6914 14702 6926 14705
rect 7298 14702 7310 14705
rect 7362 14702 7374 14754
rect 4510 14690 4562 14702
rect 28366 14690 28418 14702
rect 55022 14754 55074 14766
rect 55022 14690 55074 14702
rect 3166 14642 3218 14654
rect 3166 14578 3218 14590
rect 3502 14642 3554 14654
rect 3502 14578 3554 14590
rect 4958 14642 5010 14654
rect 4958 14578 5010 14590
rect 6862 14642 6914 14654
rect 6862 14578 6914 14590
rect 7310 14642 7362 14654
rect 12350 14642 12402 14654
rect 8418 14590 8430 14642
rect 8482 14590 8494 14642
rect 7310 14578 7362 14590
rect 12350 14578 12402 14590
rect 14590 14642 14642 14654
rect 14590 14578 14642 14590
rect 17054 14642 17106 14654
rect 24894 14642 24946 14654
rect 18386 14590 18398 14642
rect 18450 14590 18462 14642
rect 20514 14590 20526 14642
rect 20578 14590 20590 14642
rect 17054 14578 17106 14590
rect 24894 14578 24946 14590
rect 25342 14642 25394 14654
rect 25342 14578 25394 14590
rect 27358 14642 27410 14654
rect 49422 14642 49474 14654
rect 33618 14590 33630 14642
rect 33682 14590 33694 14642
rect 35634 14590 35646 14642
rect 35698 14590 35710 14642
rect 44930 14590 44942 14642
rect 44994 14590 45006 14642
rect 27358 14578 27410 14590
rect 49422 14578 49474 14590
rect 49870 14642 49922 14654
rect 49870 14578 49922 14590
rect 50654 14642 50706 14654
rect 50654 14578 50706 14590
rect 50990 14642 51042 14654
rect 50990 14578 51042 14590
rect 52782 14642 52834 14654
rect 56130 14590 56142 14642
rect 56194 14590 56206 14642
rect 52782 14578 52834 14590
rect 3390 14530 3442 14542
rect 4846 14530 4898 14542
rect 10670 14530 10722 14542
rect 1810 14478 1822 14530
rect 1874 14478 1886 14530
rect 3826 14478 3838 14530
rect 3890 14478 3902 14530
rect 4162 14478 4174 14530
rect 4226 14478 4238 14530
rect 7634 14478 7646 14530
rect 7698 14478 7710 14530
rect 8754 14478 8766 14530
rect 8818 14478 8830 14530
rect 9874 14478 9886 14530
rect 9938 14478 9950 14530
rect 3390 14466 3442 14478
rect 4846 14466 4898 14478
rect 10670 14466 10722 14478
rect 11230 14530 11282 14542
rect 11230 14466 11282 14478
rect 12126 14530 12178 14542
rect 12126 14466 12178 14478
rect 12798 14530 12850 14542
rect 12798 14466 12850 14478
rect 15598 14530 15650 14542
rect 21310 14530 21362 14542
rect 22206 14530 22258 14542
rect 16594 14478 16606 14530
rect 16658 14478 16670 14530
rect 17714 14478 17726 14530
rect 17778 14478 17790 14530
rect 21746 14478 21758 14530
rect 21810 14478 21822 14530
rect 15598 14466 15650 14478
rect 21310 14466 21362 14478
rect 22206 14466 22258 14478
rect 22654 14530 22706 14542
rect 25454 14530 25506 14542
rect 24210 14478 24222 14530
rect 24274 14478 24286 14530
rect 24658 14478 24670 14530
rect 24722 14478 24734 14530
rect 22654 14466 22706 14478
rect 25454 14466 25506 14478
rect 25902 14530 25954 14542
rect 25902 14466 25954 14478
rect 28254 14530 28306 14542
rect 28254 14466 28306 14478
rect 29374 14530 29426 14542
rect 29374 14466 29426 14478
rect 32958 14530 33010 14542
rect 37102 14530 37154 14542
rect 40350 14530 40402 14542
rect 44270 14530 44322 14542
rect 35522 14478 35534 14530
rect 35586 14478 35598 14530
rect 38658 14478 38670 14530
rect 38722 14478 38734 14530
rect 40002 14478 40014 14530
rect 40066 14478 40078 14530
rect 40898 14478 40910 14530
rect 40962 14478 40974 14530
rect 41122 14478 41134 14530
rect 41186 14478 41198 14530
rect 41794 14478 41806 14530
rect 41858 14478 41870 14530
rect 32958 14466 33010 14478
rect 37102 14466 37154 14478
rect 40350 14466 40402 14478
rect 44270 14466 44322 14478
rect 45390 14530 45442 14542
rect 48750 14530 48802 14542
rect 46162 14478 46174 14530
rect 46226 14478 46238 14530
rect 46834 14478 46846 14530
rect 46898 14478 46910 14530
rect 47282 14478 47294 14530
rect 47346 14478 47358 14530
rect 45390 14466 45442 14478
rect 48750 14466 48802 14478
rect 51326 14530 51378 14542
rect 51326 14466 51378 14478
rect 51774 14530 51826 14542
rect 51774 14466 51826 14478
rect 51998 14530 52050 14542
rect 51998 14466 52050 14478
rect 52558 14530 52610 14542
rect 52558 14466 52610 14478
rect 52894 14530 52946 14542
rect 52894 14466 52946 14478
rect 53118 14530 53170 14542
rect 55794 14478 55806 14530
rect 55858 14478 55870 14530
rect 57586 14478 57598 14530
rect 57650 14478 57662 14530
rect 53118 14466 53170 14478
rect 2382 14418 2434 14430
rect 2382 14354 2434 14366
rect 2718 14418 2770 14430
rect 2718 14354 2770 14366
rect 3054 14418 3106 14430
rect 3054 14354 3106 14366
rect 10782 14418 10834 14430
rect 10782 14354 10834 14366
rect 11006 14418 11058 14430
rect 11006 14354 11058 14366
rect 12574 14418 12626 14430
rect 12574 14354 12626 14366
rect 14142 14418 14194 14430
rect 14142 14354 14194 14366
rect 15038 14418 15090 14430
rect 15038 14354 15090 14366
rect 15262 14418 15314 14430
rect 15262 14354 15314 14366
rect 15934 14418 15986 14430
rect 15934 14354 15986 14366
rect 16270 14418 16322 14430
rect 16270 14354 16322 14366
rect 22766 14418 22818 14430
rect 22766 14354 22818 14366
rect 23550 14418 23602 14430
rect 27918 14418 27970 14430
rect 26786 14366 26798 14418
rect 26850 14366 26862 14418
rect 23550 14354 23602 14366
rect 27918 14354 27970 14366
rect 29150 14418 29202 14430
rect 29150 14354 29202 14366
rect 29710 14418 29762 14430
rect 29710 14354 29762 14366
rect 30270 14418 30322 14430
rect 30270 14354 30322 14366
rect 31726 14418 31778 14430
rect 31726 14354 31778 14366
rect 32062 14418 32114 14430
rect 32062 14354 32114 14366
rect 34862 14418 34914 14430
rect 34862 14354 34914 14366
rect 34974 14418 35026 14430
rect 34974 14354 35026 14366
rect 36430 14418 36482 14430
rect 39230 14418 39282 14430
rect 38882 14366 38894 14418
rect 38946 14366 38958 14418
rect 36430 14354 36482 14366
rect 39230 14354 39282 14366
rect 39342 14418 39394 14430
rect 39342 14354 39394 14366
rect 39790 14418 39842 14430
rect 39790 14354 39842 14366
rect 40238 14418 40290 14430
rect 46286 14418 46338 14430
rect 40786 14366 40798 14418
rect 40850 14366 40862 14418
rect 43922 14366 43934 14418
rect 43986 14366 43998 14418
rect 40238 14354 40290 14366
rect 46286 14354 46338 14366
rect 48078 14418 48130 14430
rect 48078 14354 48130 14366
rect 48302 14418 48354 14430
rect 54686 14418 54738 14430
rect 51090 14366 51102 14418
rect 51154 14366 51166 14418
rect 56130 14366 56142 14418
rect 56194 14366 56206 14418
rect 48302 14354 48354 14366
rect 54686 14354 54738 14366
rect 2046 14306 2098 14318
rect 2046 14242 2098 14254
rect 6078 14306 6130 14318
rect 6078 14242 6130 14254
rect 6414 14306 6466 14318
rect 13694 14306 13746 14318
rect 11554 14254 11566 14306
rect 11618 14254 11630 14306
rect 6414 14242 6466 14254
rect 13694 14242 13746 14254
rect 15150 14306 15202 14318
rect 15150 14242 15202 14254
rect 16382 14306 16434 14318
rect 16382 14242 16434 14254
rect 22990 14306 23042 14318
rect 22990 14242 23042 14254
rect 23214 14306 23266 14318
rect 23214 14242 23266 14254
rect 23438 14306 23490 14318
rect 23438 14242 23490 14254
rect 25230 14306 25282 14318
rect 25230 14242 25282 14254
rect 26462 14306 26514 14318
rect 26462 14242 26514 14254
rect 28366 14306 28418 14318
rect 28366 14242 28418 14254
rect 29262 14306 29314 14318
rect 29262 14242 29314 14254
rect 29934 14306 29986 14318
rect 29934 14242 29986 14254
rect 30158 14306 30210 14318
rect 30158 14242 30210 14254
rect 32510 14306 32562 14318
rect 32510 14242 32562 14254
rect 33070 14306 33122 14318
rect 33070 14242 33122 14254
rect 33294 14306 33346 14318
rect 33294 14242 33346 14254
rect 34078 14306 34130 14318
rect 34078 14242 34130 14254
rect 34638 14306 34690 14318
rect 34638 14242 34690 14254
rect 39566 14306 39618 14318
rect 39566 14242 39618 14254
rect 47406 14306 47458 14318
rect 47406 14242 47458 14254
rect 48190 14306 48242 14318
rect 48190 14242 48242 14254
rect 48862 14306 48914 14318
rect 48862 14242 48914 14254
rect 49086 14306 49138 14318
rect 49086 14242 49138 14254
rect 54910 14306 54962 14318
rect 54910 14242 54962 14254
rect 1344 14138 58731 14172
rect 1344 14086 15520 14138
rect 15572 14086 15624 14138
rect 15676 14086 15728 14138
rect 15780 14086 29827 14138
rect 29879 14086 29931 14138
rect 29983 14086 30035 14138
rect 30087 14086 44134 14138
rect 44186 14086 44238 14138
rect 44290 14086 44342 14138
rect 44394 14086 58441 14138
rect 58493 14086 58545 14138
rect 58597 14086 58649 14138
rect 58701 14086 58731 14138
rect 1344 14052 58731 14086
rect 3502 13970 3554 13982
rect 3502 13906 3554 13918
rect 7646 13970 7698 13982
rect 7646 13906 7698 13918
rect 8766 13970 8818 13982
rect 8766 13906 8818 13918
rect 14030 13970 14082 13982
rect 14030 13906 14082 13918
rect 15598 13970 15650 13982
rect 24782 13970 24834 13982
rect 27358 13970 27410 13982
rect 30718 13970 30770 13982
rect 16482 13918 16494 13970
rect 16546 13918 16558 13970
rect 25218 13918 25230 13970
rect 25282 13918 25294 13970
rect 28018 13918 28030 13970
rect 28082 13918 28094 13970
rect 15598 13906 15650 13918
rect 24782 13906 24834 13918
rect 27358 13906 27410 13918
rect 30718 13906 30770 13918
rect 33182 13970 33234 13982
rect 33182 13906 33234 13918
rect 35086 13970 35138 13982
rect 35086 13906 35138 13918
rect 35646 13970 35698 13982
rect 55918 13970 55970 13982
rect 37314 13918 37326 13970
rect 37378 13918 37390 13970
rect 40338 13918 40350 13970
rect 40402 13918 40414 13970
rect 49746 13918 49758 13970
rect 49810 13918 49822 13970
rect 53890 13918 53902 13970
rect 53954 13918 53966 13970
rect 35646 13906 35698 13918
rect 55918 13906 55970 13918
rect 2382 13858 2434 13870
rect 2382 13794 2434 13806
rect 2718 13858 2770 13870
rect 2718 13794 2770 13806
rect 2942 13858 2994 13870
rect 2942 13794 2994 13806
rect 3726 13858 3778 13870
rect 3726 13794 3778 13806
rect 7310 13858 7362 13870
rect 8990 13858 9042 13870
rect 8306 13806 8318 13858
rect 8370 13806 8382 13858
rect 7310 13794 7362 13806
rect 8990 13794 9042 13806
rect 11790 13858 11842 13870
rect 11790 13794 11842 13806
rect 12462 13858 12514 13870
rect 12462 13794 12514 13806
rect 13358 13858 13410 13870
rect 13358 13794 13410 13806
rect 13470 13858 13522 13870
rect 23886 13858 23938 13870
rect 30942 13858 30994 13870
rect 14354 13806 14366 13858
rect 14418 13806 14430 13858
rect 21634 13806 21646 13858
rect 21698 13806 21710 13858
rect 29474 13806 29486 13858
rect 29538 13806 29550 13858
rect 13470 13794 13522 13806
rect 23886 13794 23938 13806
rect 30942 13794 30994 13806
rect 31502 13858 31554 13870
rect 33070 13858 33122 13870
rect 53006 13858 53058 13870
rect 31938 13806 31950 13858
rect 32002 13806 32014 13858
rect 36418 13806 36430 13858
rect 36482 13806 36494 13858
rect 41234 13806 41246 13858
rect 41298 13806 41310 13858
rect 43474 13806 43486 13858
rect 43538 13806 43550 13858
rect 46274 13806 46286 13858
rect 46338 13806 46350 13858
rect 47282 13806 47294 13858
rect 47346 13806 47358 13858
rect 48738 13806 48750 13858
rect 48802 13806 48814 13858
rect 51090 13806 51102 13858
rect 51154 13806 51166 13858
rect 31502 13794 31554 13806
rect 33070 13794 33122 13806
rect 53006 13794 53058 13806
rect 56030 13858 56082 13870
rect 56030 13794 56082 13806
rect 6750 13746 6802 13758
rect 2034 13694 2046 13746
rect 2098 13694 2110 13746
rect 4722 13694 4734 13746
rect 4786 13694 4798 13746
rect 6290 13694 6302 13746
rect 6354 13694 6366 13746
rect 6750 13682 6802 13694
rect 7982 13746 8034 13758
rect 7982 13682 8034 13694
rect 9550 13746 9602 13758
rect 12126 13746 12178 13758
rect 10546 13694 10558 13746
rect 10610 13694 10622 13746
rect 9550 13682 9602 13694
rect 12126 13682 12178 13694
rect 12798 13746 12850 13758
rect 12798 13682 12850 13694
rect 12910 13746 12962 13758
rect 12910 13682 12962 13694
rect 13694 13746 13746 13758
rect 15374 13746 15426 13758
rect 16830 13746 16882 13758
rect 18174 13746 18226 13758
rect 25566 13746 25618 13758
rect 14690 13694 14702 13746
rect 14754 13694 14766 13746
rect 16034 13694 16046 13746
rect 16098 13694 16110 13746
rect 16594 13694 16606 13746
rect 16658 13694 16670 13746
rect 17378 13694 17390 13746
rect 17442 13694 17454 13746
rect 17938 13694 17950 13746
rect 18002 13694 18014 13746
rect 21410 13694 21422 13746
rect 21474 13694 21486 13746
rect 22082 13694 22094 13746
rect 22146 13694 22158 13746
rect 23426 13694 23438 13746
rect 23490 13694 23502 13746
rect 13694 13682 13746 13694
rect 15374 13682 15426 13694
rect 16830 13682 16882 13694
rect 18174 13682 18226 13694
rect 25566 13682 25618 13694
rect 25902 13746 25954 13758
rect 25902 13682 25954 13694
rect 26462 13746 26514 13758
rect 31614 13746 31666 13758
rect 28578 13694 28590 13746
rect 28642 13694 28654 13746
rect 30482 13694 30494 13746
rect 30546 13694 30558 13746
rect 26462 13682 26514 13694
rect 31614 13682 31666 13694
rect 33294 13746 33346 13758
rect 33294 13682 33346 13694
rect 33742 13746 33794 13758
rect 53566 13746 53618 13758
rect 55358 13746 55410 13758
rect 36754 13694 36766 13746
rect 36818 13694 36830 13746
rect 37314 13694 37326 13746
rect 37378 13694 37390 13746
rect 42466 13694 42478 13746
rect 42530 13694 42542 13746
rect 44594 13694 44606 13746
rect 44658 13694 44670 13746
rect 47842 13694 47854 13746
rect 47906 13694 47918 13746
rect 49074 13694 49086 13746
rect 49138 13694 49150 13746
rect 49634 13694 49646 13746
rect 49698 13694 49710 13746
rect 51650 13694 51662 13746
rect 51714 13694 51726 13746
rect 52322 13694 52334 13746
rect 52386 13694 52398 13746
rect 54898 13694 54910 13746
rect 54962 13694 54974 13746
rect 56690 13694 56702 13746
rect 56754 13694 56766 13746
rect 57250 13694 57262 13746
rect 57314 13694 57326 13746
rect 57586 13694 57598 13746
rect 57650 13694 57662 13746
rect 33742 13682 33794 13694
rect 53566 13682 53618 13694
rect 55358 13682 55410 13694
rect 8878 13634 8930 13646
rect 11566 13634 11618 13646
rect 2146 13582 2158 13634
rect 2210 13582 2222 13634
rect 3938 13582 3950 13634
rect 4002 13631 4014 13634
rect 4162 13631 4174 13634
rect 4002 13585 4174 13631
rect 4002 13582 4014 13585
rect 4162 13582 4174 13585
rect 4226 13582 4238 13634
rect 10098 13582 10110 13634
rect 10162 13582 10174 13634
rect 10658 13582 10670 13634
rect 10722 13582 10734 13634
rect 8878 13570 8930 13582
rect 11566 13570 11618 13582
rect 12574 13634 12626 13646
rect 12574 13570 12626 13582
rect 14926 13634 14978 13646
rect 14926 13570 14978 13582
rect 18062 13634 18114 13646
rect 18062 13570 18114 13582
rect 18622 13634 18674 13646
rect 18622 13570 18674 13582
rect 19070 13634 19122 13646
rect 19070 13570 19122 13582
rect 19742 13634 19794 13646
rect 19742 13570 19794 13582
rect 20190 13634 20242 13646
rect 20190 13570 20242 13582
rect 20638 13634 20690 13646
rect 20638 13570 20690 13582
rect 20974 13634 21026 13646
rect 27022 13634 27074 13646
rect 32286 13634 32338 13646
rect 22418 13582 22430 13634
rect 22482 13582 22494 13634
rect 23090 13582 23102 13634
rect 23154 13582 23166 13634
rect 30034 13582 30046 13634
rect 30098 13582 30110 13634
rect 20974 13570 21026 13582
rect 27022 13570 27074 13582
rect 32286 13570 32338 13582
rect 32510 13634 32562 13646
rect 32510 13570 32562 13582
rect 33966 13634 34018 13646
rect 33966 13570 34018 13582
rect 34190 13634 34242 13646
rect 34190 13570 34242 13582
rect 34526 13634 34578 13646
rect 34526 13570 34578 13582
rect 39790 13634 39842 13646
rect 50318 13634 50370 13646
rect 41122 13582 41134 13634
rect 41186 13582 41198 13634
rect 46050 13582 46062 13634
rect 46114 13582 46126 13634
rect 39790 13570 39842 13582
rect 50318 13570 50370 13582
rect 53342 13634 53394 13646
rect 54674 13582 54686 13634
rect 54738 13582 54750 13634
rect 57810 13582 57822 13634
rect 57874 13582 57886 13634
rect 53342 13570 53394 13582
rect 3054 13522 3106 13534
rect 3054 13458 3106 13470
rect 3390 13522 3442 13534
rect 9774 13522 9826 13534
rect 6514 13470 6526 13522
rect 6578 13470 6590 13522
rect 3390 13458 3442 13470
rect 9774 13458 9826 13470
rect 10894 13522 10946 13534
rect 10894 13458 10946 13470
rect 15038 13522 15090 13534
rect 15038 13458 15090 13470
rect 15710 13522 15762 13534
rect 30606 13522 30658 13534
rect 16258 13470 16270 13522
rect 16322 13470 16334 13522
rect 17602 13470 17614 13522
rect 17666 13470 17678 13522
rect 19170 13470 19182 13522
rect 19234 13519 19246 13522
rect 19954 13519 19966 13522
rect 19234 13473 19966 13519
rect 19234 13470 19246 13473
rect 19954 13470 19966 13473
rect 20018 13470 20030 13522
rect 15710 13458 15762 13470
rect 30606 13458 30658 13470
rect 31502 13522 31554 13534
rect 31502 13458 31554 13470
rect 40014 13522 40066 13534
rect 40014 13458 40066 13470
rect 55918 13522 55970 13534
rect 55918 13458 55970 13470
rect 1344 13354 58576 13388
rect 1344 13302 8367 13354
rect 8419 13302 8471 13354
rect 8523 13302 8575 13354
rect 8627 13302 22674 13354
rect 22726 13302 22778 13354
rect 22830 13302 22882 13354
rect 22934 13302 36981 13354
rect 37033 13302 37085 13354
rect 37137 13302 37189 13354
rect 37241 13302 51288 13354
rect 51340 13302 51392 13354
rect 51444 13302 51496 13354
rect 51548 13302 58576 13354
rect 1344 13268 58576 13302
rect 41358 13186 41410 13198
rect 15250 13134 15262 13186
rect 15314 13134 15326 13186
rect 40226 13134 40238 13186
rect 40290 13134 40302 13186
rect 41358 13122 41410 13134
rect 41694 13186 41746 13198
rect 41694 13122 41746 13134
rect 50766 13186 50818 13198
rect 50766 13122 50818 13134
rect 5070 13074 5122 13086
rect 5070 13010 5122 13022
rect 6526 13074 6578 13086
rect 22766 13074 22818 13086
rect 9538 13022 9550 13074
rect 9602 13022 9614 13074
rect 17154 13022 17166 13074
rect 17218 13022 17230 13074
rect 19282 13022 19294 13074
rect 19346 13022 19358 13074
rect 6526 13010 6578 13022
rect 22766 13010 22818 13022
rect 24894 13074 24946 13086
rect 24894 13010 24946 13022
rect 31054 13074 31106 13086
rect 41134 13074 41186 13086
rect 34850 13022 34862 13074
rect 34914 13022 34926 13074
rect 39330 13022 39342 13074
rect 39394 13022 39406 13074
rect 39890 13022 39902 13074
rect 39954 13022 39966 13074
rect 31054 13010 31106 13022
rect 41134 13010 41186 13022
rect 43598 13074 43650 13086
rect 52110 13074 52162 13086
rect 45490 13022 45502 13074
rect 45554 13022 45566 13074
rect 48962 13022 48974 13074
rect 49026 13022 49038 13074
rect 49858 13022 49870 13074
rect 49922 13022 49934 13074
rect 55458 13022 55470 13074
rect 55522 13022 55534 13074
rect 58034 13022 58046 13074
rect 58098 13022 58110 13074
rect 43598 13010 43650 13022
rect 52110 13010 52162 13022
rect 15822 12962 15874 12974
rect 20302 12962 20354 12974
rect 3490 12910 3502 12962
rect 3554 12910 3566 12962
rect 4386 12910 4398 12962
rect 4450 12910 4462 12962
rect 4834 12910 4846 12962
rect 4898 12910 4910 12962
rect 8082 12910 8094 12962
rect 8146 12910 8158 12962
rect 12450 12910 12462 12962
rect 12514 12910 12526 12962
rect 15250 12910 15262 12962
rect 15314 12910 15326 12962
rect 16370 12910 16382 12962
rect 16434 12910 16446 12962
rect 15822 12898 15874 12910
rect 20302 12898 20354 12910
rect 23550 12962 23602 12974
rect 23550 12898 23602 12910
rect 24446 12962 24498 12974
rect 24446 12898 24498 12910
rect 24670 12962 24722 12974
rect 26014 12962 26066 12974
rect 26462 12962 26514 12974
rect 25666 12910 25678 12962
rect 25730 12910 25742 12962
rect 26226 12910 26238 12962
rect 26290 12910 26302 12962
rect 24670 12898 24722 12910
rect 26014 12898 26066 12910
rect 26462 12898 26514 12910
rect 26686 12962 26738 12974
rect 26686 12898 26738 12910
rect 29150 12962 29202 12974
rect 29150 12898 29202 12910
rect 29374 12962 29426 12974
rect 29374 12898 29426 12910
rect 29934 12962 29986 12974
rect 29934 12898 29986 12910
rect 30270 12962 30322 12974
rect 30270 12898 30322 12910
rect 31166 12962 31218 12974
rect 37886 12962 37938 12974
rect 44270 12962 44322 12974
rect 46846 12962 46898 12974
rect 49534 12962 49586 12974
rect 51214 12962 51266 12974
rect 32722 12910 32734 12962
rect 32786 12910 32798 12962
rect 33618 12910 33630 12962
rect 33682 12910 33694 12962
rect 34962 12910 34974 12962
rect 35026 12910 35038 12962
rect 37426 12910 37438 12962
rect 37490 12910 37502 12962
rect 38546 12910 38558 12962
rect 38610 12910 38622 12962
rect 40226 12910 40238 12962
rect 40290 12910 40302 12962
rect 45266 12910 45278 12962
rect 45330 12910 45342 12962
rect 46274 12910 46286 12962
rect 46338 12910 46350 12962
rect 47506 12910 47518 12962
rect 47570 12910 47582 12962
rect 50194 12910 50206 12962
rect 50258 12910 50270 12962
rect 50418 12910 50430 12962
rect 50482 12910 50494 12962
rect 51426 12910 51438 12962
rect 51490 12910 51502 12962
rect 56578 12910 56590 12962
rect 56642 12910 56654 12962
rect 31166 12898 31218 12910
rect 37886 12898 37938 12910
rect 44270 12898 44322 12910
rect 46846 12898 46898 12910
rect 49534 12898 49586 12910
rect 51214 12898 51266 12910
rect 2046 12850 2098 12862
rect 2046 12786 2098 12798
rect 2382 12850 2434 12862
rect 2382 12786 2434 12798
rect 3726 12850 3778 12862
rect 3726 12786 3778 12798
rect 5742 12850 5794 12862
rect 8542 12850 8594 12862
rect 6626 12798 6638 12850
rect 6690 12798 6702 12850
rect 5742 12786 5794 12798
rect 8542 12786 8594 12798
rect 8878 12850 8930 12862
rect 8878 12786 8930 12798
rect 9214 12850 9266 12862
rect 13470 12850 13522 12862
rect 11666 12798 11678 12850
rect 11730 12798 11742 12850
rect 9214 12786 9266 12798
rect 13470 12786 13522 12798
rect 13806 12850 13858 12862
rect 19966 12850 20018 12862
rect 15586 12798 15598 12850
rect 15650 12798 15662 12850
rect 13806 12786 13858 12798
rect 19966 12786 20018 12798
rect 25118 12850 25170 12862
rect 25118 12786 25170 12798
rect 25342 12850 25394 12862
rect 25342 12786 25394 12798
rect 26910 12850 26962 12862
rect 26910 12786 26962 12798
rect 27022 12850 27074 12862
rect 27022 12786 27074 12798
rect 27470 12850 27522 12862
rect 27470 12786 27522 12798
rect 30158 12850 30210 12862
rect 30158 12786 30210 12798
rect 30942 12850 30994 12862
rect 35646 12850 35698 12862
rect 49758 12850 49810 12862
rect 32386 12798 32398 12850
rect 32450 12798 32462 12850
rect 45154 12798 45166 12850
rect 45218 12798 45230 12850
rect 48626 12798 48638 12850
rect 48690 12798 48702 12850
rect 30942 12786 30994 12798
rect 35646 12786 35698 12798
rect 49758 12786 49810 12798
rect 50654 12850 50706 12862
rect 57362 12798 57374 12850
rect 57426 12798 57438 12850
rect 50654 12786 50706 12798
rect 2718 12738 2770 12750
rect 5630 12738 5682 12750
rect 3042 12686 3054 12738
rect 3106 12686 3118 12738
rect 2718 12674 2770 12686
rect 5630 12674 5682 12686
rect 13022 12738 13074 12750
rect 13022 12674 13074 12686
rect 14254 12738 14306 12750
rect 14254 12674 14306 12686
rect 14814 12738 14866 12750
rect 14814 12674 14866 12686
rect 15038 12738 15090 12750
rect 15038 12674 15090 12686
rect 20078 12738 20130 12750
rect 20078 12674 20130 12686
rect 20862 12738 20914 12750
rect 20862 12674 20914 12686
rect 21758 12738 21810 12750
rect 21758 12674 21810 12686
rect 22206 12738 22258 12750
rect 22206 12674 22258 12686
rect 22990 12738 23042 12750
rect 22990 12674 23042 12686
rect 23886 12738 23938 12750
rect 23886 12674 23938 12686
rect 25678 12738 25730 12750
rect 25678 12674 25730 12686
rect 27358 12738 27410 12750
rect 27358 12674 27410 12686
rect 28030 12738 28082 12750
rect 28030 12674 28082 12686
rect 29262 12738 29314 12750
rect 29262 12674 29314 12686
rect 29598 12738 29650 12750
rect 29598 12674 29650 12686
rect 30718 12738 30770 12750
rect 33954 12686 33966 12738
rect 34018 12686 34030 12738
rect 43922 12686 43934 12738
rect 43986 12686 43998 12738
rect 46162 12686 46174 12738
rect 46226 12686 46238 12738
rect 30718 12674 30770 12686
rect 1344 12570 58731 12604
rect 1344 12518 15520 12570
rect 15572 12518 15624 12570
rect 15676 12518 15728 12570
rect 15780 12518 29827 12570
rect 29879 12518 29931 12570
rect 29983 12518 30035 12570
rect 30087 12518 44134 12570
rect 44186 12518 44238 12570
rect 44290 12518 44342 12570
rect 44394 12518 58441 12570
rect 58493 12518 58545 12570
rect 58597 12518 58649 12570
rect 58701 12518 58731 12570
rect 1344 12484 58731 12518
rect 5518 12402 5570 12414
rect 5518 12338 5570 12350
rect 7870 12402 7922 12414
rect 7870 12338 7922 12350
rect 8094 12402 8146 12414
rect 8094 12338 8146 12350
rect 10782 12402 10834 12414
rect 10782 12338 10834 12350
rect 11230 12402 11282 12414
rect 11230 12338 11282 12350
rect 17390 12402 17442 12414
rect 28254 12402 28306 12414
rect 23986 12350 23998 12402
rect 24050 12350 24062 12402
rect 17390 12338 17442 12350
rect 28254 12338 28306 12350
rect 28926 12402 28978 12414
rect 28926 12338 28978 12350
rect 32062 12402 32114 12414
rect 32062 12338 32114 12350
rect 32286 12402 32338 12414
rect 33630 12402 33682 12414
rect 40014 12402 40066 12414
rect 45614 12402 45666 12414
rect 33394 12350 33406 12402
rect 33458 12350 33470 12402
rect 37314 12350 37326 12402
rect 37378 12350 37390 12402
rect 44034 12350 44046 12402
rect 44098 12350 44110 12402
rect 32286 12338 32338 12350
rect 33630 12338 33682 12350
rect 40014 12338 40066 12350
rect 45614 12338 45666 12350
rect 47182 12402 47234 12414
rect 47182 12338 47234 12350
rect 47854 12402 47906 12414
rect 47854 12338 47906 12350
rect 48302 12402 48354 12414
rect 48302 12338 48354 12350
rect 48862 12402 48914 12414
rect 48862 12338 48914 12350
rect 55470 12402 55522 12414
rect 55470 12338 55522 12350
rect 56702 12402 56754 12414
rect 56702 12338 56754 12350
rect 57598 12402 57650 12414
rect 57598 12338 57650 12350
rect 5182 12290 5234 12302
rect 5182 12226 5234 12238
rect 7758 12290 7810 12302
rect 7758 12226 7810 12238
rect 8318 12290 8370 12302
rect 8318 12226 8370 12238
rect 9550 12290 9602 12302
rect 9550 12226 9602 12238
rect 9886 12290 9938 12302
rect 15598 12290 15650 12302
rect 10434 12238 10446 12290
rect 10498 12238 10510 12290
rect 12338 12238 12350 12290
rect 12402 12238 12414 12290
rect 9886 12226 9938 12238
rect 15598 12226 15650 12238
rect 15822 12290 15874 12302
rect 15822 12226 15874 12238
rect 18174 12290 18226 12302
rect 22430 12290 22482 12302
rect 19842 12238 19854 12290
rect 19906 12238 19918 12290
rect 18174 12226 18226 12238
rect 22430 12226 22482 12238
rect 24558 12290 24610 12302
rect 31278 12290 31330 12302
rect 27122 12238 27134 12290
rect 27186 12238 27198 12290
rect 29922 12238 29934 12290
rect 29986 12238 29998 12290
rect 24558 12226 24610 12238
rect 31278 12226 31330 12238
rect 33854 12290 33906 12302
rect 33854 12226 33906 12238
rect 36990 12290 37042 12302
rect 36990 12226 37042 12238
rect 39342 12290 39394 12302
rect 39342 12226 39394 12238
rect 39566 12290 39618 12302
rect 39566 12226 39618 12238
rect 40126 12290 40178 12302
rect 40126 12226 40178 12238
rect 44382 12290 44434 12302
rect 44382 12226 44434 12238
rect 44718 12290 44770 12302
rect 56590 12290 56642 12302
rect 52322 12238 52334 12290
rect 52386 12238 52398 12290
rect 44718 12226 44770 12238
rect 56590 12226 56642 12238
rect 56814 12290 56866 12302
rect 56814 12226 56866 12238
rect 57262 12290 57314 12302
rect 57262 12226 57314 12238
rect 57374 12290 57426 12302
rect 57374 12226 57426 12238
rect 6302 12178 6354 12190
rect 6974 12178 7026 12190
rect 1922 12126 1934 12178
rect 1986 12126 1998 12178
rect 6626 12126 6638 12178
rect 6690 12126 6702 12178
rect 6302 12114 6354 12126
rect 6974 12114 7026 12126
rect 7198 12178 7250 12190
rect 17838 12178 17890 12190
rect 22542 12178 22594 12190
rect 23550 12178 23602 12190
rect 7522 12126 7534 12178
rect 7586 12126 7598 12178
rect 11554 12126 11566 12178
rect 11618 12126 11630 12178
rect 16482 12126 16494 12178
rect 16546 12126 16558 12178
rect 17378 12126 17390 12178
rect 17442 12126 17454 12178
rect 19058 12126 19070 12178
rect 19122 12126 19134 12178
rect 22978 12126 22990 12178
rect 23042 12126 23054 12178
rect 23426 12126 23438 12178
rect 23490 12126 23502 12178
rect 7198 12114 7250 12126
rect 17838 12114 17890 12126
rect 22542 12114 22594 12126
rect 23550 12114 23602 12126
rect 23662 12178 23714 12190
rect 23662 12114 23714 12126
rect 24334 12178 24386 12190
rect 27918 12178 27970 12190
rect 25554 12126 25566 12178
rect 25618 12126 25630 12178
rect 26226 12126 26238 12178
rect 26290 12126 26302 12178
rect 27234 12126 27246 12178
rect 27298 12126 27310 12178
rect 24334 12114 24386 12126
rect 27918 12114 27970 12126
rect 28254 12178 28306 12190
rect 28254 12114 28306 12126
rect 28478 12178 28530 12190
rect 28478 12114 28530 12126
rect 30942 12178 30994 12190
rect 30942 12114 30994 12126
rect 31390 12178 31442 12190
rect 31390 12114 31442 12126
rect 31950 12178 32002 12190
rect 33966 12178 34018 12190
rect 37662 12178 37714 12190
rect 33170 12126 33182 12178
rect 33234 12126 33246 12178
rect 36306 12126 36318 12178
rect 36370 12126 36382 12178
rect 36754 12126 36766 12178
rect 36818 12126 36830 12178
rect 31950 12114 32002 12126
rect 33966 12114 34018 12126
rect 37662 12114 37714 12126
rect 39230 12178 39282 12190
rect 39230 12114 39282 12126
rect 39678 12178 39730 12190
rect 39678 12114 39730 12126
rect 40350 12178 40402 12190
rect 45838 12178 45890 12190
rect 41122 12126 41134 12178
rect 41186 12126 41198 12178
rect 42466 12126 42478 12178
rect 42530 12126 42542 12178
rect 43810 12126 43822 12178
rect 43874 12126 43886 12178
rect 45042 12126 45054 12178
rect 45106 12126 45118 12178
rect 45378 12126 45390 12178
rect 45442 12126 45454 12178
rect 40350 12114 40402 12126
rect 45838 12114 45890 12126
rect 46174 12178 46226 12190
rect 46174 12114 46226 12126
rect 46398 12178 46450 12190
rect 46398 12114 46450 12126
rect 46622 12178 46674 12190
rect 46622 12114 46674 12126
rect 47294 12178 47346 12190
rect 49410 12126 49422 12178
rect 49474 12126 49486 12178
rect 50754 12126 50766 12178
rect 50818 12126 50830 12178
rect 53554 12126 53566 12178
rect 53618 12126 53630 12178
rect 47294 12114 47346 12126
rect 6078 12066 6130 12078
rect 2706 12014 2718 12066
rect 2770 12014 2782 12066
rect 4834 11987 4846 12039
rect 4898 11987 4910 12039
rect 6078 12002 6130 12014
rect 7086 12066 7138 12078
rect 7086 12002 7138 12014
rect 9102 12066 9154 12078
rect 9102 12002 9154 12014
rect 14478 12066 14530 12078
rect 18846 12066 18898 12078
rect 31054 12066 31106 12078
rect 16594 12014 16606 12066
rect 16658 12014 16670 12066
rect 21970 12014 21982 12066
rect 22034 12014 22046 12066
rect 25330 12014 25342 12066
rect 25394 12014 25406 12066
rect 26114 12014 26126 12066
rect 26178 12014 26190 12066
rect 27570 12014 27582 12066
rect 27634 12014 27646 12066
rect 14478 12002 14530 12014
rect 18846 12002 18898 12014
rect 31054 12002 31106 12014
rect 34414 12066 34466 12078
rect 34414 12002 34466 12014
rect 34862 12066 34914 12078
rect 34862 12002 34914 12014
rect 37886 12066 37938 12078
rect 45726 12066 45778 12078
rect 41010 12014 41022 12066
rect 41074 12014 41086 12066
rect 37886 12002 37938 12014
rect 45726 12002 45778 12014
rect 46286 12066 46338 12078
rect 49746 12014 49758 12066
rect 49810 12014 49822 12066
rect 51538 12014 51550 12066
rect 51602 12014 51614 12066
rect 52098 12014 52110 12066
rect 52162 12014 52174 12066
rect 55570 12014 55582 12066
rect 55634 12014 55646 12066
rect 46286 12002 46338 12014
rect 23214 11954 23266 11966
rect 47182 11954 47234 11966
rect 17602 11902 17614 11954
rect 17666 11902 17678 11954
rect 42690 11902 42702 11954
rect 42754 11902 42766 11954
rect 23214 11890 23266 11902
rect 47182 11890 47234 11902
rect 54910 11954 54962 11966
rect 54910 11890 54962 11902
rect 55246 11954 55298 11966
rect 55246 11890 55298 11902
rect 1344 11786 58576 11820
rect 1344 11734 8367 11786
rect 8419 11734 8471 11786
rect 8523 11734 8575 11786
rect 8627 11734 22674 11786
rect 22726 11734 22778 11786
rect 22830 11734 22882 11786
rect 22934 11734 36981 11786
rect 37033 11734 37085 11786
rect 37137 11734 37189 11786
rect 37241 11734 51288 11786
rect 51340 11734 51392 11786
rect 51444 11734 51496 11786
rect 51548 11734 58576 11786
rect 1344 11700 58576 11734
rect 2046 11618 2098 11630
rect 2046 11554 2098 11566
rect 3166 11618 3218 11630
rect 7646 11618 7698 11630
rect 10670 11618 10722 11630
rect 4162 11566 4174 11618
rect 4226 11566 4238 11618
rect 9202 11566 9214 11618
rect 9266 11566 9278 11618
rect 3166 11554 3218 11566
rect 7646 11554 7698 11566
rect 10670 11554 10722 11566
rect 18622 11618 18674 11630
rect 18622 11554 18674 11566
rect 20750 11618 20802 11630
rect 40910 11618 40962 11630
rect 30258 11566 30270 11618
rect 30322 11566 30334 11618
rect 35746 11566 35758 11618
rect 35810 11566 35822 11618
rect 20750 11554 20802 11566
rect 40910 11554 40962 11566
rect 41246 11618 41298 11630
rect 51550 11618 51602 11630
rect 45714 11566 45726 11618
rect 45778 11566 45790 11618
rect 41246 11554 41298 11566
rect 51550 11554 51602 11566
rect 11902 11506 11954 11518
rect 19070 11506 19122 11518
rect 27022 11506 27074 11518
rect 7970 11454 7982 11506
rect 8034 11454 8046 11506
rect 12674 11454 12686 11506
rect 12738 11454 12750 11506
rect 15026 11454 15038 11506
rect 15090 11454 15102 11506
rect 17154 11454 17166 11506
rect 17218 11454 17230 11506
rect 20514 11454 20526 11506
rect 20578 11454 20590 11506
rect 11902 11442 11954 11454
rect 19070 11442 19122 11454
rect 27022 11442 27074 11454
rect 27806 11506 27858 11518
rect 27806 11442 27858 11454
rect 31054 11506 31106 11518
rect 39230 11506 39282 11518
rect 33506 11454 33518 11506
rect 33570 11454 33582 11506
rect 35858 11454 35870 11506
rect 35922 11454 35934 11506
rect 37090 11454 37102 11506
rect 37154 11454 37166 11506
rect 31054 11442 31106 11454
rect 39230 11442 39282 11454
rect 39566 11506 39618 11518
rect 43486 11506 43538 11518
rect 47966 11506 48018 11518
rect 57934 11506 57986 11518
rect 39890 11454 39902 11506
rect 39954 11454 39966 11506
rect 46722 11454 46734 11506
rect 46786 11454 46798 11506
rect 50978 11454 50990 11506
rect 51042 11454 51054 11506
rect 39566 11442 39618 11454
rect 43486 11442 43538 11454
rect 47966 11442 48018 11454
rect 57934 11442 57986 11454
rect 2494 11394 2546 11406
rect 3614 11394 3666 11406
rect 4734 11394 4786 11406
rect 9438 11394 9490 11406
rect 1922 11342 1934 11394
rect 1986 11342 1998 11394
rect 3042 11342 3054 11394
rect 3106 11342 3118 11394
rect 3378 11342 3390 11394
rect 3442 11342 3454 11394
rect 4050 11342 4062 11394
rect 4114 11342 4126 11394
rect 5842 11342 5854 11394
rect 5906 11342 5918 11394
rect 6738 11342 6750 11394
rect 6802 11342 6814 11394
rect 8306 11342 8318 11394
rect 8370 11342 8382 11394
rect 9202 11342 9214 11394
rect 9266 11342 9278 11394
rect 2494 11330 2546 11342
rect 3614 11330 3666 11342
rect 4734 11330 4786 11342
rect 9438 11330 9490 11342
rect 10222 11394 10274 11406
rect 10222 11330 10274 11342
rect 10558 11394 10610 11406
rect 17838 11394 17890 11406
rect 10882 11342 10894 11394
rect 10946 11342 10958 11394
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 12338 11342 12350 11394
rect 12402 11342 12414 11394
rect 14354 11342 14366 11394
rect 14418 11342 14430 11394
rect 10558 11330 10610 11342
rect 17838 11330 17890 11342
rect 18174 11394 18226 11406
rect 19966 11394 20018 11406
rect 18722 11342 18734 11394
rect 18786 11342 18798 11394
rect 19730 11342 19742 11394
rect 19794 11342 19806 11394
rect 18174 11330 18226 11342
rect 19966 11330 20018 11342
rect 21310 11394 21362 11406
rect 22206 11394 22258 11406
rect 21970 11342 21982 11394
rect 22034 11342 22046 11394
rect 21310 11330 21362 11342
rect 22206 11330 22258 11342
rect 22542 11394 22594 11406
rect 24222 11394 24274 11406
rect 23314 11342 23326 11394
rect 23378 11342 23390 11394
rect 23762 11342 23774 11394
rect 23826 11342 23838 11394
rect 22542 11330 22594 11342
rect 24222 11330 24274 11342
rect 24558 11394 24610 11406
rect 26350 11394 26402 11406
rect 25218 11342 25230 11394
rect 25282 11342 25294 11394
rect 24558 11330 24610 11342
rect 26350 11330 26402 11342
rect 26574 11394 26626 11406
rect 26574 11330 26626 11342
rect 26910 11394 26962 11406
rect 26910 11330 26962 11342
rect 27134 11394 27186 11406
rect 27134 11330 27186 11342
rect 29598 11394 29650 11406
rect 29598 11330 29650 11342
rect 29822 11394 29874 11406
rect 29822 11330 29874 11342
rect 31166 11394 31218 11406
rect 31166 11330 31218 11342
rect 31502 11394 31554 11406
rect 31502 11330 31554 11342
rect 31950 11394 32002 11406
rect 31950 11330 32002 11342
rect 32062 11394 32114 11406
rect 32062 11330 32114 11342
rect 32398 11394 32450 11406
rect 48190 11394 48242 11406
rect 33282 11342 33294 11394
rect 33346 11342 33358 11394
rect 34514 11342 34526 11394
rect 34578 11342 34590 11394
rect 35746 11342 35758 11394
rect 35810 11342 35822 11394
rect 36530 11342 36542 11394
rect 36594 11342 36606 11394
rect 38546 11342 38558 11394
rect 38610 11342 38622 11394
rect 40226 11342 40238 11394
rect 40290 11342 40302 11394
rect 40898 11342 40910 11394
rect 40962 11342 40974 11394
rect 45378 11342 45390 11394
rect 45442 11342 45454 11394
rect 45714 11342 45726 11394
rect 45778 11342 45790 11394
rect 47058 11342 47070 11394
rect 47122 11342 47134 11394
rect 32398 11330 32450 11342
rect 48190 11330 48242 11342
rect 49422 11394 49474 11406
rect 49422 11330 49474 11342
rect 49758 11394 49810 11406
rect 49970 11342 49982 11394
rect 50034 11342 50046 11394
rect 50530 11342 50542 11394
rect 50594 11342 50606 11394
rect 54786 11342 54798 11394
rect 54850 11342 54862 11394
rect 55234 11342 55246 11394
rect 55298 11342 55310 11394
rect 49758 11330 49810 11342
rect 7086 11282 7138 11294
rect 2258 11230 2270 11282
rect 2322 11230 2334 11282
rect 4498 11230 4510 11282
rect 4562 11230 4574 11282
rect 5954 11230 5966 11282
rect 6018 11230 6030 11282
rect 7086 11218 7138 11230
rect 7870 11282 7922 11294
rect 7870 11218 7922 11230
rect 8654 11282 8706 11294
rect 8654 11218 8706 11230
rect 9774 11282 9826 11294
rect 17950 11282 18002 11294
rect 13458 11230 13470 11282
rect 13522 11230 13534 11282
rect 9774 11218 9826 11230
rect 17950 11218 18002 11230
rect 22878 11282 22930 11294
rect 22878 11218 22930 11230
rect 25678 11282 25730 11294
rect 29710 11282 29762 11294
rect 26002 11230 26014 11282
rect 26066 11230 26078 11282
rect 25678 11218 25730 11230
rect 29710 11218 29762 11230
rect 30718 11282 30770 11294
rect 30718 11218 30770 11230
rect 31726 11282 31778 11294
rect 31726 11218 31778 11230
rect 32734 11282 32786 11294
rect 32734 11218 32786 11230
rect 33966 11282 34018 11294
rect 45166 11282 45218 11294
rect 37314 11230 37326 11282
rect 37378 11230 37390 11282
rect 33966 11218 34018 11230
rect 45166 11218 45218 11230
rect 47630 11282 47682 11294
rect 47630 11218 47682 11230
rect 49534 11282 49586 11294
rect 51774 11282 51826 11294
rect 50642 11230 50654 11282
rect 50706 11230 50718 11282
rect 49534 11218 49586 11230
rect 51774 11218 51826 11230
rect 54574 11282 54626 11294
rect 56130 11230 56142 11282
rect 56194 11230 56206 11282
rect 57474 11230 57486 11282
rect 57538 11230 57550 11282
rect 54574 11218 54626 11230
rect 2382 11170 2434 11182
rect 2382 11106 2434 11118
rect 2830 11170 2882 11182
rect 2830 11106 2882 11118
rect 3950 11170 4002 11182
rect 8542 11170 8594 11182
rect 6290 11118 6302 11170
rect 6354 11118 6366 11170
rect 3950 11106 4002 11118
rect 8542 11106 8594 11118
rect 8990 11170 9042 11182
rect 8990 11106 9042 11118
rect 10334 11170 10386 11182
rect 10334 11106 10386 11118
rect 13806 11170 13858 11182
rect 13806 11106 13858 11118
rect 20526 11170 20578 11182
rect 20526 11106 20578 11118
rect 22766 11170 22818 11182
rect 22766 11106 22818 11118
rect 27358 11170 27410 11182
rect 27358 11106 27410 11118
rect 28366 11170 28418 11182
rect 28366 11106 28418 11118
rect 30942 11170 30994 11182
rect 30942 11106 30994 11118
rect 32510 11170 32562 11182
rect 32510 11106 32562 11118
rect 34302 11170 34354 11182
rect 34302 11106 34354 11118
rect 41806 11170 41858 11182
rect 41806 11106 41858 11118
rect 42142 11170 42194 11182
rect 42142 11106 42194 11118
rect 42590 11170 42642 11182
rect 42590 11106 42642 11118
rect 43038 11170 43090 11182
rect 43038 11106 43090 11118
rect 45950 11170 46002 11182
rect 51662 11170 51714 11182
rect 48514 11118 48526 11170
rect 48578 11118 48590 11170
rect 56242 11118 56254 11170
rect 56306 11118 56318 11170
rect 45950 11106 46002 11118
rect 51662 11106 51714 11118
rect 1344 11002 58731 11036
rect 1344 10950 15520 11002
rect 15572 10950 15624 11002
rect 15676 10950 15728 11002
rect 15780 10950 29827 11002
rect 29879 10950 29931 11002
rect 29983 10950 30035 11002
rect 30087 10950 44134 11002
rect 44186 10950 44238 11002
rect 44290 10950 44342 11002
rect 44394 10950 58441 11002
rect 58493 10950 58545 11002
rect 58597 10950 58649 11002
rect 58701 10950 58731 11002
rect 1344 10916 58731 10950
rect 2046 10834 2098 10846
rect 2046 10770 2098 10782
rect 5742 10834 5794 10846
rect 5742 10770 5794 10782
rect 16382 10834 16434 10846
rect 16382 10770 16434 10782
rect 25342 10834 25394 10846
rect 25342 10770 25394 10782
rect 25566 10834 25618 10846
rect 32174 10834 32226 10846
rect 35870 10834 35922 10846
rect 26114 10782 26126 10834
rect 26178 10782 26190 10834
rect 26898 10782 26910 10834
rect 26962 10782 26974 10834
rect 33058 10782 33070 10834
rect 33122 10782 33134 10834
rect 25566 10770 25618 10782
rect 32174 10770 32226 10782
rect 35870 10770 35922 10782
rect 36430 10834 36482 10846
rect 36430 10770 36482 10782
rect 36878 10834 36930 10846
rect 36878 10770 36930 10782
rect 42926 10834 42978 10846
rect 42926 10770 42978 10782
rect 43262 10834 43314 10846
rect 43262 10770 43314 10782
rect 45166 10834 45218 10846
rect 53890 10782 53902 10834
rect 53954 10782 53966 10834
rect 45166 10770 45218 10782
rect 1710 10722 1762 10734
rect 7870 10722 7922 10734
rect 22766 10722 22818 10734
rect 35310 10722 35362 10734
rect 3266 10670 3278 10722
rect 3330 10670 3342 10722
rect 12674 10670 12686 10722
rect 12738 10670 12750 10722
rect 13570 10670 13582 10722
rect 13634 10670 13646 10722
rect 14690 10670 14702 10722
rect 14754 10670 14766 10722
rect 20066 10670 20078 10722
rect 20130 10670 20142 10722
rect 27346 10670 27358 10722
rect 27410 10670 27422 10722
rect 31042 10670 31054 10722
rect 31106 10670 31118 10722
rect 1710 10658 1762 10670
rect 7870 10658 7922 10670
rect 22766 10658 22818 10670
rect 35310 10658 35362 10670
rect 36318 10722 36370 10734
rect 36318 10658 36370 10670
rect 37102 10722 37154 10734
rect 37102 10658 37154 10670
rect 37214 10722 37266 10734
rect 42702 10722 42754 10734
rect 39554 10670 39566 10722
rect 39618 10670 39630 10722
rect 37214 10658 37266 10670
rect 42702 10658 42754 10670
rect 46398 10722 46450 10734
rect 46398 10658 46450 10670
rect 48750 10722 48802 10734
rect 55346 10670 55358 10722
rect 55410 10670 55422 10722
rect 48750 10658 48802 10670
rect 8990 10610 9042 10622
rect 10670 10610 10722 10622
rect 19294 10610 19346 10622
rect 25230 10610 25282 10622
rect 27806 10610 27858 10622
rect 2482 10558 2494 10610
rect 2546 10558 2558 10610
rect 6626 10558 6638 10610
rect 6690 10558 6702 10610
rect 7410 10558 7422 10610
rect 7474 10558 7486 10610
rect 8306 10558 8318 10610
rect 8370 10558 8382 10610
rect 9874 10558 9886 10610
rect 9938 10558 9950 10610
rect 10434 10558 10446 10610
rect 10498 10558 10510 10610
rect 12562 10558 12574 10610
rect 12626 10558 12638 10610
rect 14242 10558 14254 10610
rect 14306 10558 14318 10610
rect 14914 10558 14926 10610
rect 14978 10558 14990 10610
rect 19730 10558 19742 10610
rect 19794 10558 19806 10610
rect 21634 10558 21646 10610
rect 21698 10558 21710 10610
rect 22978 10558 22990 10610
rect 23042 10558 23054 10610
rect 23762 10558 23774 10610
rect 23826 10558 23838 10610
rect 24322 10558 24334 10610
rect 24386 10558 24398 10610
rect 26114 10558 26126 10610
rect 26178 10558 26190 10610
rect 27458 10558 27470 10610
rect 27522 10558 27534 10610
rect 8990 10546 9042 10558
rect 10670 10546 10722 10558
rect 19294 10546 19346 10558
rect 25230 10546 25282 10558
rect 27806 10546 27858 10558
rect 28814 10610 28866 10622
rect 31726 10610 31778 10622
rect 29698 10558 29710 10610
rect 29762 10558 29774 10610
rect 30930 10558 30942 10610
rect 30994 10558 31006 10610
rect 28814 10546 28866 10558
rect 31726 10546 31778 10558
rect 33406 10610 33458 10622
rect 33406 10546 33458 10558
rect 34302 10610 34354 10622
rect 34302 10546 34354 10558
rect 34862 10610 34914 10622
rect 34862 10546 34914 10558
rect 35086 10610 35138 10622
rect 35086 10546 35138 10558
rect 35422 10610 35474 10622
rect 35422 10546 35474 10558
rect 35758 10610 35810 10622
rect 38894 10610 38946 10622
rect 40910 10610 40962 10622
rect 36642 10558 36654 10610
rect 36706 10558 36718 10610
rect 39218 10558 39230 10610
rect 39282 10558 39294 10610
rect 40114 10558 40126 10610
rect 40178 10558 40190 10610
rect 35758 10546 35810 10558
rect 38894 10546 38946 10558
rect 40910 10546 40962 10558
rect 41806 10610 41858 10622
rect 43150 10610 43202 10622
rect 44606 10610 44658 10622
rect 42242 10558 42254 10610
rect 42306 10558 42318 10610
rect 44258 10558 44270 10610
rect 44322 10558 44334 10610
rect 41806 10546 41858 10558
rect 43150 10546 43202 10558
rect 44606 10546 44658 10558
rect 44718 10610 44770 10622
rect 44718 10546 44770 10558
rect 45054 10610 45106 10622
rect 45054 10546 45106 10558
rect 45950 10610 46002 10622
rect 45950 10546 46002 10558
rect 46174 10610 46226 10622
rect 47058 10558 47070 10610
rect 47122 10558 47134 10610
rect 49298 10558 49310 10610
rect 49362 10558 49374 10610
rect 51314 10558 51326 10610
rect 51378 10558 51390 10610
rect 54450 10558 54462 10610
rect 54514 10558 54526 10610
rect 57138 10558 57150 10610
rect 57202 10558 57214 10610
rect 46174 10546 46226 10558
rect 5854 10498 5906 10510
rect 5394 10446 5406 10498
rect 5458 10446 5470 10498
rect 5854 10434 5906 10446
rect 6414 10498 6466 10510
rect 6414 10434 6466 10446
rect 10558 10498 10610 10510
rect 15934 10498 15986 10510
rect 10994 10446 11006 10498
rect 11058 10446 11070 10498
rect 15250 10446 15262 10498
rect 15314 10446 15326 10498
rect 10558 10434 10610 10446
rect 15934 10434 15986 10446
rect 16830 10498 16882 10510
rect 16830 10434 16882 10446
rect 17838 10498 17890 10510
rect 17838 10434 17890 10446
rect 18174 10498 18226 10510
rect 18174 10434 18226 10446
rect 19182 10498 19234 10510
rect 22206 10498 22258 10510
rect 33966 10498 34018 10510
rect 41134 10498 41186 10510
rect 46286 10498 46338 10510
rect 19618 10446 19630 10498
rect 19682 10446 19694 10498
rect 23426 10446 23438 10498
rect 23490 10446 23502 10498
rect 28242 10446 28254 10498
rect 28306 10446 28318 10498
rect 29810 10446 29822 10498
rect 29874 10446 29886 10498
rect 30818 10446 30830 10498
rect 30882 10446 30894 10498
rect 39330 10446 39342 10498
rect 39394 10446 39406 10498
rect 41458 10446 41470 10498
rect 41522 10446 41534 10498
rect 43250 10446 43262 10498
rect 43314 10446 43326 10498
rect 19182 10434 19234 10446
rect 22206 10434 22258 10446
rect 33966 10434 34018 10446
rect 41134 10434 41186 10446
rect 46286 10434 46338 10446
rect 46846 10498 46898 10510
rect 51998 10498 52050 10510
rect 57598 10498 57650 10510
rect 49522 10446 49534 10498
rect 49586 10446 49598 10498
rect 51538 10446 51550 10498
rect 51602 10446 51614 10498
rect 55906 10446 55918 10498
rect 55970 10446 55982 10498
rect 56802 10446 56814 10498
rect 56866 10446 56878 10498
rect 46846 10434 46898 10446
rect 51998 10434 52050 10446
rect 57598 10434 57650 10446
rect 18398 10386 18450 10398
rect 6738 10334 6750 10386
rect 6802 10334 6814 10386
rect 10098 10334 10110 10386
rect 10162 10334 10174 10386
rect 18398 10322 18450 10334
rect 18734 10386 18786 10398
rect 18734 10322 18786 10334
rect 20862 10386 20914 10398
rect 20862 10322 20914 10334
rect 28702 10386 28754 10398
rect 35870 10386 35922 10398
rect 31714 10334 31726 10386
rect 31778 10383 31790 10386
rect 32050 10383 32062 10386
rect 31778 10337 32062 10383
rect 31778 10334 31790 10337
rect 32050 10334 32062 10337
rect 32114 10334 32126 10386
rect 33618 10334 33630 10386
rect 33682 10383 33694 10386
rect 33954 10383 33966 10386
rect 33682 10337 33966 10383
rect 33682 10334 33694 10337
rect 33954 10334 33966 10337
rect 34018 10334 34030 10386
rect 28702 10322 28754 10334
rect 35870 10322 35922 10334
rect 45166 10386 45218 10398
rect 45166 10322 45218 10334
rect 46734 10386 46786 10398
rect 46734 10322 46786 10334
rect 1344 10218 58576 10252
rect 1344 10166 8367 10218
rect 8419 10166 8471 10218
rect 8523 10166 8575 10218
rect 8627 10166 22674 10218
rect 22726 10166 22778 10218
rect 22830 10166 22882 10218
rect 22934 10166 36981 10218
rect 37033 10166 37085 10218
rect 37137 10166 37189 10218
rect 37241 10166 51288 10218
rect 51340 10166 51392 10218
rect 51444 10166 51496 10218
rect 51548 10166 58576 10218
rect 1344 10132 58576 10166
rect 11006 10050 11058 10062
rect 40014 10050 40066 10062
rect 29586 9998 29598 10050
rect 29650 9998 29662 10050
rect 35634 9998 35646 10050
rect 35698 9998 35710 10050
rect 11006 9986 11058 9998
rect 40014 9986 40066 9998
rect 48750 10050 48802 10062
rect 50642 9998 50654 10050
rect 50706 9998 50718 10050
rect 48750 9986 48802 9998
rect 5182 9938 5234 9950
rect 2482 9886 2494 9938
rect 2546 9886 2558 9938
rect 4610 9886 4622 9938
rect 4674 9886 4686 9938
rect 5182 9874 5234 9886
rect 5854 9938 5906 9950
rect 5854 9874 5906 9886
rect 12462 9938 12514 9950
rect 12462 9874 12514 9886
rect 12798 9938 12850 9950
rect 32622 9938 32674 9950
rect 17490 9886 17502 9938
rect 17554 9886 17566 9938
rect 19618 9886 19630 9938
rect 19682 9886 19694 9938
rect 25218 9886 25230 9938
rect 25282 9886 25294 9938
rect 26002 9886 26014 9938
rect 26066 9886 26078 9938
rect 27234 9886 27246 9938
rect 27298 9886 27310 9938
rect 27906 9886 27918 9938
rect 27970 9886 27982 9938
rect 29810 9886 29822 9938
rect 29874 9886 29886 9938
rect 12798 9874 12850 9886
rect 32622 9874 32674 9886
rect 34190 9938 34242 9950
rect 36206 9938 36258 9950
rect 39678 9938 39730 9950
rect 34850 9886 34862 9938
rect 34914 9886 34926 9938
rect 39218 9886 39230 9938
rect 39282 9886 39294 9938
rect 34190 9874 34242 9886
rect 36206 9874 36258 9886
rect 39678 9874 39730 9886
rect 40126 9938 40178 9950
rect 54910 9938 54962 9950
rect 45154 9886 45166 9938
rect 45218 9886 45230 9938
rect 47058 9886 47070 9938
rect 47122 9886 47134 9938
rect 56578 9886 56590 9938
rect 56642 9886 56654 9938
rect 40126 9874 40178 9886
rect 54910 9874 54962 9886
rect 11454 9826 11506 9838
rect 16382 9826 16434 9838
rect 30942 9826 30994 9838
rect 1810 9774 1822 9826
rect 1874 9774 1886 9826
rect 6290 9774 6302 9826
rect 6354 9774 6366 9826
rect 7970 9774 7982 9826
rect 8034 9774 8046 9826
rect 9650 9774 9662 9826
rect 9714 9774 9726 9826
rect 10658 9774 10670 9826
rect 10722 9774 10734 9826
rect 14466 9774 14478 9826
rect 14530 9774 14542 9826
rect 15138 9774 15150 9826
rect 15202 9774 15214 9826
rect 16818 9774 16830 9826
rect 16882 9774 16894 9826
rect 20626 9774 20638 9826
rect 20690 9774 20702 9826
rect 21970 9774 21982 9826
rect 22034 9774 22046 9826
rect 23650 9774 23662 9826
rect 23714 9774 23726 9826
rect 25778 9774 25790 9826
rect 25842 9774 25854 9826
rect 26114 9774 26126 9826
rect 26178 9774 26190 9826
rect 27010 9774 27022 9826
rect 27074 9774 27086 9826
rect 28242 9774 28254 9826
rect 28306 9774 28318 9826
rect 29698 9774 29710 9826
rect 29762 9774 29774 9826
rect 30706 9774 30718 9826
rect 30770 9774 30782 9826
rect 11454 9762 11506 9774
rect 16382 9762 16434 9774
rect 30942 9762 30994 9774
rect 32062 9826 32114 9838
rect 32062 9762 32114 9774
rect 33630 9826 33682 9838
rect 33630 9762 33682 9774
rect 34078 9826 34130 9838
rect 34078 9762 34130 9774
rect 34302 9826 34354 9838
rect 42814 9826 42866 9838
rect 35074 9774 35086 9826
rect 35138 9774 35150 9826
rect 38994 9774 39006 9826
rect 39058 9774 39070 9826
rect 40338 9774 40350 9826
rect 40402 9774 40414 9826
rect 41010 9774 41022 9826
rect 41074 9774 41086 9826
rect 34302 9762 34354 9774
rect 42814 9762 42866 9774
rect 44046 9826 44098 9838
rect 45950 9826 46002 9838
rect 48526 9826 48578 9838
rect 44818 9774 44830 9826
rect 44882 9774 44894 9826
rect 45042 9774 45054 9826
rect 45106 9774 45118 9826
rect 46610 9774 46622 9826
rect 46674 9774 46686 9826
rect 47394 9774 47406 9826
rect 47458 9774 47470 9826
rect 44046 9762 44098 9774
rect 45950 9762 46002 9774
rect 48526 9762 48578 9774
rect 48974 9826 49026 9838
rect 48974 9762 49026 9774
rect 49310 9826 49362 9838
rect 50990 9826 51042 9838
rect 49522 9774 49534 9826
rect 49586 9774 49598 9826
rect 50530 9774 50542 9826
rect 50594 9774 50606 9826
rect 49310 9762 49362 9774
rect 50990 9762 51042 9774
rect 52558 9826 52610 9838
rect 52558 9762 52610 9774
rect 53118 9826 53170 9838
rect 53118 9762 53170 9774
rect 55134 9826 55186 9838
rect 55794 9774 55806 9826
rect 55858 9774 55870 9826
rect 57138 9774 57150 9826
rect 57202 9774 57214 9826
rect 55134 9762 55186 9774
rect 12910 9714 12962 9726
rect 15822 9714 15874 9726
rect 21534 9714 21586 9726
rect 31390 9714 31442 9726
rect 33070 9714 33122 9726
rect 6738 9662 6750 9714
rect 6802 9662 6814 9714
rect 9426 9662 9438 9714
rect 9490 9662 9502 9714
rect 11218 9662 11230 9714
rect 11282 9662 11294 9714
rect 13906 9662 13918 9714
rect 13970 9662 13982 9714
rect 20738 9662 20750 9714
rect 20802 9662 20814 9714
rect 22530 9662 22542 9714
rect 22594 9662 22606 9714
rect 23538 9662 23550 9714
rect 23602 9662 23614 9714
rect 26674 9662 26686 9714
rect 26738 9662 26750 9714
rect 27122 9662 27134 9714
rect 27186 9662 27198 9714
rect 31714 9662 31726 9714
rect 31778 9662 31790 9714
rect 12910 9650 12962 9662
rect 15822 9650 15874 9662
rect 21534 9650 21586 9662
rect 31390 9650 31442 9662
rect 33070 9650 33122 9662
rect 33182 9714 33234 9726
rect 33182 9650 33234 9662
rect 40686 9714 40738 9726
rect 40686 9650 40738 9662
rect 41694 9714 41746 9726
rect 41694 9650 41746 9662
rect 42030 9714 42082 9726
rect 42030 9650 42082 9662
rect 42142 9714 42194 9726
rect 43710 9714 43762 9726
rect 43474 9662 43486 9714
rect 43538 9662 43550 9714
rect 42142 9650 42194 9662
rect 43710 9650 43762 9662
rect 45278 9714 45330 9726
rect 45278 9650 45330 9662
rect 45614 9714 45666 9726
rect 45614 9650 45666 9662
rect 45726 9714 45778 9726
rect 53006 9714 53058 9726
rect 46498 9662 46510 9714
rect 46562 9662 46574 9714
rect 46946 9662 46958 9714
rect 47010 9662 47022 9714
rect 57698 9662 57710 9714
rect 57762 9662 57774 9714
rect 45726 9650 45778 9662
rect 53006 9650 53058 9662
rect 8766 9602 8818 9614
rect 8766 9538 8818 9550
rect 10670 9602 10722 9614
rect 10670 9538 10722 9550
rect 12014 9602 12066 9614
rect 21646 9602 21698 9614
rect 20178 9550 20190 9602
rect 20242 9550 20254 9602
rect 12014 9538 12066 9550
rect 21646 9538 21698 9550
rect 32846 9602 32898 9614
rect 32846 9538 32898 9550
rect 38334 9602 38386 9614
rect 38334 9538 38386 9550
rect 40798 9602 40850 9614
rect 40798 9538 40850 9550
rect 41470 9602 41522 9614
rect 41470 9538 41522 9550
rect 41582 9602 41634 9614
rect 41582 9538 41634 9550
rect 42366 9602 42418 9614
rect 42366 9538 42418 9550
rect 42478 9602 42530 9614
rect 42478 9538 42530 9550
rect 42702 9602 42754 9614
rect 42702 9538 42754 9550
rect 43150 9602 43202 9614
rect 43150 9538 43202 9550
rect 43934 9602 43986 9614
rect 43934 9538 43986 9550
rect 48078 9602 48130 9614
rect 48078 9538 48130 9550
rect 52894 9602 52946 9614
rect 55458 9550 55470 9602
rect 55522 9550 55534 9602
rect 52894 9538 52946 9550
rect 1344 9434 58731 9468
rect 1344 9382 15520 9434
rect 15572 9382 15624 9434
rect 15676 9382 15728 9434
rect 15780 9382 29827 9434
rect 29879 9382 29931 9434
rect 29983 9382 30035 9434
rect 30087 9382 44134 9434
rect 44186 9382 44238 9434
rect 44290 9382 44342 9434
rect 44394 9382 58441 9434
rect 58493 9382 58545 9434
rect 58597 9382 58649 9434
rect 58701 9382 58731 9434
rect 1344 9348 58731 9382
rect 2158 9266 2210 9278
rect 1810 9214 1822 9266
rect 1874 9214 1886 9266
rect 2158 9202 2210 9214
rect 3054 9266 3106 9278
rect 3054 9202 3106 9214
rect 3726 9266 3778 9278
rect 3726 9202 3778 9214
rect 4062 9266 4114 9278
rect 4062 9202 4114 9214
rect 4846 9266 4898 9278
rect 22318 9266 22370 9278
rect 6738 9214 6750 9266
rect 6802 9214 6814 9266
rect 20402 9214 20414 9266
rect 20466 9214 20478 9266
rect 4846 9202 4898 9214
rect 22318 9202 22370 9214
rect 29374 9266 29426 9278
rect 29374 9202 29426 9214
rect 31166 9266 31218 9278
rect 31166 9202 31218 9214
rect 31278 9266 31330 9278
rect 31278 9202 31330 9214
rect 39342 9266 39394 9278
rect 39342 9202 39394 9214
rect 39678 9266 39730 9278
rect 39678 9202 39730 9214
rect 40910 9266 40962 9278
rect 40910 9202 40962 9214
rect 43934 9266 43986 9278
rect 43934 9202 43986 9214
rect 44494 9266 44546 9278
rect 44494 9202 44546 9214
rect 44942 9266 44994 9278
rect 44942 9202 44994 9214
rect 45278 9266 45330 9278
rect 45278 9202 45330 9214
rect 46286 9266 46338 9278
rect 46286 9202 46338 9214
rect 47406 9266 47458 9278
rect 47406 9202 47458 9214
rect 53902 9266 53954 9278
rect 57474 9214 57486 9266
rect 57538 9214 57550 9266
rect 53902 9202 53954 9214
rect 2718 9154 2770 9166
rect 9886 9154 9938 9166
rect 16494 9154 16546 9166
rect 5842 9102 5854 9154
rect 5906 9102 5918 9154
rect 7522 9102 7534 9154
rect 7586 9102 7598 9154
rect 10994 9102 11006 9154
rect 11058 9102 11070 9154
rect 15026 9102 15038 9154
rect 15090 9102 15102 9154
rect 2718 9090 2770 9102
rect 9886 9090 9938 9102
rect 16494 9090 16546 9102
rect 16830 9154 16882 9166
rect 27806 9154 27858 9166
rect 23090 9102 23102 9154
rect 23154 9102 23166 9154
rect 24546 9102 24558 9154
rect 24610 9102 24622 9154
rect 16830 9090 16882 9102
rect 27806 9090 27858 9102
rect 30494 9154 30546 9166
rect 46510 9154 46562 9166
rect 32162 9102 32174 9154
rect 32226 9102 32238 9154
rect 37314 9102 37326 9154
rect 37378 9102 37390 9154
rect 40002 9102 40014 9154
rect 40066 9102 40078 9154
rect 41234 9102 41246 9154
rect 41298 9102 41310 9154
rect 41794 9102 41806 9154
rect 41858 9102 41870 9154
rect 30494 9090 30546 9102
rect 46510 9090 46562 9102
rect 50990 9154 51042 9166
rect 50990 9090 51042 9102
rect 52334 9154 52386 9166
rect 52334 9090 52386 9102
rect 53790 9154 53842 9166
rect 53790 9090 53842 9102
rect 54014 9154 54066 9166
rect 54014 9090 54066 9102
rect 54798 9154 54850 9166
rect 54798 9090 54850 9102
rect 54910 9154 54962 9166
rect 56690 9102 56702 9154
rect 56754 9102 56766 9154
rect 54910 9090 54962 9102
rect 28030 9042 28082 9054
rect 29934 9042 29986 9054
rect 5394 8990 5406 9042
rect 5458 8990 5470 9042
rect 7634 8990 7646 9042
rect 7698 8990 7710 9042
rect 9538 8990 9550 9042
rect 9602 8990 9614 9042
rect 10210 8990 10222 9042
rect 10274 8990 10286 9042
rect 13570 8990 13582 9042
rect 13634 8990 13646 9042
rect 13906 8990 13918 9042
rect 13970 8990 13982 9042
rect 17490 8990 17502 9042
rect 17554 8990 17566 9042
rect 18162 8990 18174 9042
rect 18226 8990 18238 9042
rect 22418 8990 22430 9042
rect 22482 8990 22494 9042
rect 22978 8990 22990 9042
rect 23042 8990 23054 9042
rect 24098 8990 24110 9042
rect 24162 8990 24174 9042
rect 25666 8990 25678 9042
rect 25730 8990 25742 9042
rect 25890 8990 25902 9042
rect 25954 8990 25966 9042
rect 26898 8990 26910 9042
rect 26962 8990 26974 9042
rect 27682 8990 27694 9042
rect 27746 8990 27758 9042
rect 28578 8990 28590 9042
rect 28642 8990 28654 9042
rect 28030 8978 28082 8990
rect 29934 8978 29986 8990
rect 31054 9042 31106 9054
rect 31054 8978 31106 8990
rect 31726 9042 31778 9054
rect 31726 8978 31778 8990
rect 32510 9042 32562 9054
rect 32510 8978 32562 8990
rect 33182 9042 33234 9054
rect 33182 8978 33234 8990
rect 33742 9042 33794 9054
rect 44046 9042 44098 9054
rect 34514 8990 34526 9042
rect 34578 8990 34590 9042
rect 36306 8990 36318 9042
rect 36370 8990 36382 9042
rect 36754 8990 36766 9042
rect 36818 8990 36830 9042
rect 37202 8990 37214 9042
rect 37266 8990 37278 9042
rect 38098 8990 38110 9042
rect 38162 8990 38174 9042
rect 42018 8990 42030 9042
rect 42082 8990 42094 9042
rect 42578 8990 42590 9042
rect 42642 8990 42654 9042
rect 43026 8990 43038 9042
rect 43090 8990 43102 9042
rect 33742 8978 33794 8990
rect 44046 8978 44098 8990
rect 45502 9042 45554 9054
rect 45502 8978 45554 8990
rect 45950 9042 46002 9054
rect 51886 9042 51938 9054
rect 55358 9042 55410 9054
rect 47618 8990 47630 9042
rect 47682 8990 47694 9042
rect 48850 8990 48862 9042
rect 48914 8990 48926 9042
rect 49074 8990 49086 9042
rect 49138 8990 49150 9042
rect 49746 8990 49758 9042
rect 49810 8990 49822 9042
rect 51650 8990 51662 9042
rect 51714 8990 51726 9042
rect 53106 8990 53118 9042
rect 53170 8990 53182 9042
rect 56578 8990 56590 9042
rect 56642 8990 56654 9042
rect 57474 8990 57486 9042
rect 57538 8990 57550 9042
rect 45950 8978 46002 8990
rect 51886 8978 51938 8990
rect 55358 8978 55410 8990
rect 15486 8930 15538 8942
rect 9650 8878 9662 8930
rect 9714 8878 9726 8930
rect 13122 8878 13134 8930
rect 13186 8878 13198 8930
rect 15486 8866 15538 8878
rect 15598 8930 15650 8942
rect 15598 8866 15650 8878
rect 16270 8930 16322 8942
rect 16270 8866 16322 8878
rect 20862 8930 20914 8942
rect 27918 8930 27970 8942
rect 23426 8878 23438 8930
rect 23490 8878 23502 8930
rect 24322 8878 24334 8930
rect 24386 8878 24398 8930
rect 20862 8866 20914 8878
rect 27918 8866 27970 8878
rect 29038 8930 29090 8942
rect 35534 8930 35586 8942
rect 30594 8878 30606 8930
rect 30658 8878 30670 8930
rect 34850 8878 34862 8930
rect 34914 8878 34926 8930
rect 29038 8866 29090 8878
rect 35534 8866 35586 8878
rect 35758 8930 35810 8942
rect 35758 8866 35810 8878
rect 38334 8930 38386 8942
rect 38334 8866 38386 8878
rect 38894 8930 38946 8942
rect 38894 8866 38946 8878
rect 45390 8930 45442 8942
rect 46274 8878 46286 8930
rect 46338 8878 46350 8930
rect 47506 8878 47518 8930
rect 47570 8878 47582 8930
rect 52882 8878 52894 8930
rect 52946 8878 52958 8930
rect 45390 8866 45442 8878
rect 8206 8818 8258 8830
rect 8206 8754 8258 8766
rect 8542 8818 8594 8830
rect 8542 8754 8594 8766
rect 21086 8818 21138 8830
rect 21086 8754 21138 8766
rect 21310 8818 21362 8830
rect 21310 8754 21362 8766
rect 21758 8818 21810 8830
rect 21758 8754 21810 8766
rect 26798 8818 26850 8830
rect 26798 8754 26850 8766
rect 27358 8818 27410 8830
rect 27358 8754 27410 8766
rect 30270 8818 30322 8830
rect 30270 8754 30322 8766
rect 35982 8818 36034 8830
rect 35982 8754 36034 8766
rect 38670 8818 38722 8830
rect 38670 8754 38722 8766
rect 43374 8818 43426 8830
rect 43374 8754 43426 8766
rect 43934 8818 43986 8830
rect 43934 8754 43986 8766
rect 49982 8818 50034 8830
rect 49982 8754 50034 8766
rect 54910 8818 54962 8830
rect 54910 8754 54962 8766
rect 55582 8818 55634 8830
rect 55906 8766 55918 8818
rect 55970 8766 55982 8818
rect 55582 8754 55634 8766
rect 1344 8650 58576 8684
rect 1344 8598 8367 8650
rect 8419 8598 8471 8650
rect 8523 8598 8575 8650
rect 8627 8598 22674 8650
rect 22726 8598 22778 8650
rect 22830 8598 22882 8650
rect 22934 8598 36981 8650
rect 37033 8598 37085 8650
rect 37137 8598 37189 8650
rect 37241 8598 51288 8650
rect 51340 8598 51392 8650
rect 51444 8598 51496 8650
rect 51548 8598 58576 8650
rect 1344 8564 58576 8598
rect 33518 8482 33570 8494
rect 22418 8430 22430 8482
rect 22482 8430 22494 8482
rect 33518 8418 33570 8430
rect 35982 8482 36034 8494
rect 54350 8482 54402 8494
rect 41234 8430 41246 8482
rect 41298 8430 41310 8482
rect 55906 8430 55918 8482
rect 55970 8430 55982 8482
rect 57138 8430 57150 8482
rect 57202 8430 57214 8482
rect 35982 8418 36034 8430
rect 54350 8418 54402 8430
rect 5182 8370 5234 8382
rect 30606 8370 30658 8382
rect 46510 8370 46562 8382
rect 4610 8318 4622 8370
rect 4674 8318 4686 8370
rect 7746 8318 7758 8370
rect 7810 8318 7822 8370
rect 9762 8318 9774 8370
rect 9826 8318 9838 8370
rect 11890 8318 11902 8370
rect 11954 8318 11966 8370
rect 15026 8318 15038 8370
rect 15090 8318 15102 8370
rect 18498 8318 18510 8370
rect 18562 8318 18574 8370
rect 20066 8318 20078 8370
rect 20130 8318 20142 8370
rect 25554 8318 25566 8370
rect 25618 8318 25630 8370
rect 29586 8318 29598 8370
rect 29650 8318 29662 8370
rect 34738 8318 34750 8370
rect 34802 8318 34814 8370
rect 39890 8318 39902 8370
rect 39954 8318 39966 8370
rect 45378 8318 45390 8370
rect 45442 8318 45454 8370
rect 5182 8306 5234 8318
rect 30606 8306 30658 8318
rect 46510 8306 46562 8318
rect 47294 8370 47346 8382
rect 47294 8306 47346 8318
rect 47406 8370 47458 8382
rect 47406 8306 47458 8318
rect 49310 8370 49362 8382
rect 53230 8370 53282 8382
rect 55134 8370 55186 8382
rect 50194 8318 50206 8370
rect 50258 8318 50270 8370
rect 54674 8318 54686 8370
rect 54738 8318 54750 8370
rect 49310 8306 49362 8318
rect 53230 8306 53282 8318
rect 55134 8306 55186 8318
rect 56254 8370 56306 8382
rect 57362 8318 57374 8370
rect 57426 8318 57438 8370
rect 56254 8306 56306 8318
rect 12462 8258 12514 8270
rect 1810 8206 1822 8258
rect 1874 8206 1886 8258
rect 6178 8206 6190 8258
rect 6242 8206 6254 8258
rect 8978 8206 8990 8258
rect 9042 8206 9054 8258
rect 12462 8194 12514 8206
rect 13022 8258 13074 8270
rect 16494 8258 16546 8270
rect 17726 8258 17778 8270
rect 25902 8258 25954 8270
rect 13570 8206 13582 8258
rect 13634 8206 13646 8258
rect 17154 8206 17166 8258
rect 17218 8206 17230 8258
rect 18610 8206 18622 8258
rect 18674 8206 18686 8258
rect 20626 8206 20638 8258
rect 20690 8206 20702 8258
rect 22194 8206 22206 8258
rect 22258 8206 22270 8258
rect 22754 8206 22766 8258
rect 22818 8206 22830 8258
rect 23090 8206 23102 8258
rect 23154 8206 23166 8258
rect 23986 8206 23998 8258
rect 24050 8206 24062 8258
rect 24322 8206 24334 8258
rect 24386 8206 24398 8258
rect 13022 8194 13074 8206
rect 16494 8194 16546 8206
rect 17726 8194 17778 8206
rect 25902 8194 25954 8206
rect 26014 8258 26066 8270
rect 26014 8194 26066 8206
rect 26238 8258 26290 8270
rect 26238 8194 26290 8206
rect 26350 8258 26402 8270
rect 30046 8258 30098 8270
rect 36094 8258 36146 8270
rect 45726 8258 45778 8270
rect 27570 8206 27582 8258
rect 27634 8206 27646 8258
rect 27906 8206 27918 8258
rect 27970 8206 27982 8258
rect 31938 8206 31950 8258
rect 32002 8206 32014 8258
rect 32722 8206 32734 8258
rect 32786 8206 32798 8258
rect 33170 8206 33182 8258
rect 33234 8206 33246 8258
rect 37762 8206 37774 8258
rect 37826 8206 37838 8258
rect 38658 8206 38670 8258
rect 38722 8206 38734 8258
rect 42578 8206 42590 8258
rect 42642 8206 42654 8258
rect 26350 8194 26402 8206
rect 30046 8194 30098 8206
rect 36094 8194 36146 8206
rect 45726 8194 45778 8206
rect 46062 8258 46114 8270
rect 46062 8194 46114 8206
rect 46398 8258 46450 8270
rect 46398 8194 46450 8206
rect 47070 8258 47122 8270
rect 49534 8258 49586 8270
rect 54910 8258 54962 8270
rect 48178 8206 48190 8258
rect 48242 8206 48254 8258
rect 49970 8206 49982 8258
rect 50034 8206 50046 8258
rect 47070 8194 47122 8206
rect 49534 8194 49586 8206
rect 54910 8194 54962 8206
rect 55246 8258 55298 8270
rect 55246 8194 55298 8206
rect 55470 8258 55522 8270
rect 55470 8194 55522 8206
rect 56478 8258 56530 8270
rect 57138 8206 57150 8258
rect 57202 8206 57214 8258
rect 58034 8206 58046 8258
rect 58098 8206 58110 8258
rect 56478 8194 56530 8206
rect 12686 8146 12738 8158
rect 14254 8146 14306 8158
rect 2482 8094 2494 8146
rect 2546 8094 2558 8146
rect 7186 8094 7198 8146
rect 7250 8094 7262 8146
rect 13794 8094 13806 8146
rect 13858 8094 13870 8146
rect 12686 8082 12738 8094
rect 14254 8082 14306 8094
rect 14366 8146 14418 8158
rect 14366 8082 14418 8094
rect 14702 8146 14754 8158
rect 14702 8082 14754 8094
rect 15262 8146 15314 8158
rect 15262 8082 15314 8094
rect 15598 8146 15650 8158
rect 15598 8082 15650 8094
rect 15934 8146 15986 8158
rect 15934 8082 15986 8094
rect 17838 8146 17890 8158
rect 17838 8082 17890 8094
rect 19182 8146 19234 8158
rect 32174 8146 32226 8158
rect 27010 8094 27022 8146
rect 27074 8094 27086 8146
rect 28466 8094 28478 8146
rect 28530 8094 28542 8146
rect 31266 8094 31278 8146
rect 31330 8094 31342 8146
rect 19182 8082 19234 8094
rect 32174 8082 32226 8094
rect 33742 8146 33794 8158
rect 35982 8146 36034 8158
rect 40238 8146 40290 8158
rect 43934 8146 43986 8158
rect 35186 8094 35198 8146
rect 35250 8094 35262 8146
rect 37426 8094 37438 8146
rect 37490 8094 37502 8146
rect 42130 8094 42142 8146
rect 42194 8094 42206 8146
rect 43698 8094 43710 8146
rect 43762 8094 43774 8146
rect 33742 8082 33794 8094
rect 35982 8082 36034 8094
rect 40238 8082 40290 8094
rect 43934 8082 43986 8094
rect 44830 8146 44882 8158
rect 44830 8082 44882 8094
rect 47518 8146 47570 8158
rect 54574 8146 54626 8158
rect 48290 8094 48302 8146
rect 48354 8094 48366 8146
rect 48738 8094 48750 8146
rect 48802 8094 48814 8146
rect 47518 8082 47570 8094
rect 54574 8082 54626 8094
rect 8766 8034 8818 8046
rect 5730 7982 5742 8034
rect 5794 7982 5806 8034
rect 8766 7970 8818 7982
rect 12798 8034 12850 8046
rect 12798 7970 12850 7982
rect 14030 8034 14082 8046
rect 14030 7970 14082 7982
rect 14926 8034 14978 8046
rect 14926 7970 14978 7982
rect 15486 8034 15538 8046
rect 15486 7970 15538 7982
rect 21422 8034 21474 8046
rect 29150 8034 29202 8046
rect 21746 7982 21758 8034
rect 21810 7982 21822 8034
rect 28354 7982 28366 8034
rect 28418 7982 28430 8034
rect 21422 7970 21474 7982
rect 29150 7970 29202 7982
rect 30942 8034 30994 8046
rect 30942 7970 30994 7982
rect 35534 8034 35586 8046
rect 35534 7970 35586 7982
rect 44942 8034 44994 8046
rect 44942 7970 44994 7982
rect 46622 8034 46674 8046
rect 46622 7970 46674 7982
rect 53342 8034 53394 8046
rect 53342 7970 53394 7982
rect 53454 8034 53506 8046
rect 53454 7970 53506 7982
rect 54126 8034 54178 8046
rect 54126 7970 54178 7982
rect 1344 7866 58731 7900
rect 1344 7814 15520 7866
rect 15572 7814 15624 7866
rect 15676 7814 15728 7866
rect 15780 7814 29827 7866
rect 29879 7814 29931 7866
rect 29983 7814 30035 7866
rect 30087 7814 44134 7866
rect 44186 7814 44238 7866
rect 44290 7814 44342 7866
rect 44394 7814 58441 7866
rect 58493 7814 58545 7866
rect 58597 7814 58649 7866
rect 58701 7814 58731 7866
rect 1344 7780 58731 7814
rect 2270 7698 2322 7710
rect 2270 7634 2322 7646
rect 2494 7698 2546 7710
rect 2494 7634 2546 7646
rect 3838 7698 3890 7710
rect 3838 7634 3890 7646
rect 4510 7698 4562 7710
rect 4510 7634 4562 7646
rect 4958 7698 5010 7710
rect 4958 7634 5010 7646
rect 6638 7698 6690 7710
rect 17502 7698 17554 7710
rect 15026 7646 15038 7698
rect 15090 7646 15102 7698
rect 6638 7634 6690 7646
rect 17502 7634 17554 7646
rect 19294 7698 19346 7710
rect 19294 7634 19346 7646
rect 25230 7698 25282 7710
rect 25230 7634 25282 7646
rect 30830 7698 30882 7710
rect 30830 7634 30882 7646
rect 34526 7698 34578 7710
rect 34526 7634 34578 7646
rect 35422 7698 35474 7710
rect 35422 7634 35474 7646
rect 36094 7698 36146 7710
rect 36094 7634 36146 7646
rect 36318 7698 36370 7710
rect 36318 7634 36370 7646
rect 37326 7698 37378 7710
rect 37326 7634 37378 7646
rect 37774 7698 37826 7710
rect 37774 7634 37826 7646
rect 38670 7698 38722 7710
rect 44830 7698 44882 7710
rect 40002 7646 40014 7698
rect 40066 7646 40078 7698
rect 41122 7646 41134 7698
rect 41186 7646 41198 7698
rect 38670 7634 38722 7646
rect 44830 7634 44882 7646
rect 47630 7698 47682 7710
rect 47630 7634 47682 7646
rect 47854 7698 47906 7710
rect 55010 7646 55022 7698
rect 55074 7646 55086 7698
rect 47854 7634 47906 7646
rect 2830 7586 2882 7598
rect 2830 7522 2882 7534
rect 3166 7586 3218 7598
rect 14030 7586 14082 7598
rect 30942 7586 30994 7598
rect 34190 7586 34242 7598
rect 10322 7534 10334 7586
rect 10386 7534 10398 7586
rect 18946 7534 18958 7586
rect 19010 7534 19022 7586
rect 27794 7534 27806 7586
rect 27858 7534 27870 7586
rect 28802 7534 28814 7586
rect 28866 7534 28878 7586
rect 31266 7534 31278 7586
rect 31330 7534 31342 7586
rect 3166 7522 3218 7534
rect 14030 7522 14082 7534
rect 30942 7522 30994 7534
rect 34190 7522 34242 7534
rect 36430 7586 36482 7598
rect 36430 7522 36482 7534
rect 36878 7586 36930 7598
rect 36878 7522 36930 7534
rect 38782 7586 38834 7598
rect 46958 7586 47010 7598
rect 39330 7534 39342 7586
rect 39394 7534 39406 7586
rect 41570 7534 41582 7586
rect 41634 7534 41646 7586
rect 43250 7534 43262 7586
rect 43314 7534 43326 7586
rect 38782 7522 38834 7534
rect 46958 7522 47010 7534
rect 50318 7586 50370 7598
rect 54114 7534 54126 7586
rect 54178 7534 54190 7586
rect 50318 7522 50370 7534
rect 3502 7474 3554 7486
rect 3502 7410 3554 7422
rect 5406 7474 5458 7486
rect 5406 7410 5458 7422
rect 5630 7474 5682 7486
rect 5630 7410 5682 7422
rect 5966 7474 6018 7486
rect 5966 7410 6018 7422
rect 6190 7474 6242 7486
rect 6190 7410 6242 7422
rect 6862 7474 6914 7486
rect 6862 7410 6914 7422
rect 7198 7474 7250 7486
rect 29822 7474 29874 7486
rect 8194 7422 8206 7474
rect 8258 7422 8270 7474
rect 9650 7422 9662 7474
rect 9714 7422 9726 7474
rect 13570 7422 13582 7474
rect 13634 7422 13646 7474
rect 16370 7422 16382 7474
rect 16434 7422 16446 7474
rect 18050 7422 18062 7474
rect 18114 7422 18126 7474
rect 18834 7422 18846 7474
rect 18898 7422 18910 7474
rect 20402 7422 20414 7474
rect 20466 7422 20478 7474
rect 22306 7422 22318 7474
rect 22370 7422 22382 7474
rect 22978 7422 22990 7474
rect 23042 7422 23054 7474
rect 23538 7422 23550 7474
rect 23602 7422 23614 7474
rect 26786 7422 26798 7474
rect 26850 7422 26862 7474
rect 27010 7422 27022 7474
rect 27074 7422 27086 7474
rect 28354 7422 28366 7474
rect 28418 7422 28430 7474
rect 28690 7422 28702 7474
rect 28754 7422 28766 7474
rect 7198 7410 7250 7422
rect 29822 7410 29874 7422
rect 30382 7474 30434 7486
rect 30382 7410 30434 7422
rect 33518 7474 33570 7486
rect 35310 7474 35362 7486
rect 33730 7422 33742 7474
rect 33794 7422 33806 7474
rect 33518 7410 33570 7422
rect 35310 7410 35362 7422
rect 35534 7474 35586 7486
rect 35534 7410 35586 7422
rect 35982 7474 36034 7486
rect 43822 7474 43874 7486
rect 39106 7422 39118 7474
rect 39170 7422 39182 7474
rect 40114 7422 40126 7474
rect 40178 7422 40190 7474
rect 40898 7422 40910 7474
rect 40962 7422 40974 7474
rect 41458 7422 41470 7474
rect 41522 7422 41534 7474
rect 42354 7422 42366 7474
rect 42418 7422 42430 7474
rect 43474 7422 43486 7474
rect 43538 7422 43550 7474
rect 35982 7410 36034 7422
rect 43822 7410 43874 7422
rect 44606 7474 44658 7486
rect 44606 7410 44658 7422
rect 44942 7474 44994 7486
rect 47518 7474 47570 7486
rect 46386 7422 46398 7474
rect 46450 7422 46462 7474
rect 44942 7410 44994 7422
rect 47518 7410 47570 7422
rect 48078 7474 48130 7486
rect 48078 7410 48130 7422
rect 48190 7474 48242 7486
rect 50542 7474 50594 7486
rect 56926 7474 56978 7486
rect 49522 7422 49534 7474
rect 49586 7422 49598 7474
rect 51538 7422 51550 7474
rect 51602 7422 51614 7474
rect 52994 7422 53006 7474
rect 53058 7422 53070 7474
rect 54338 7422 54350 7474
rect 54402 7422 54414 7474
rect 54898 7422 54910 7474
rect 54962 7422 54974 7474
rect 57250 7422 57262 7474
rect 57314 7422 57326 7474
rect 48190 7410 48242 7422
rect 50542 7410 50594 7422
rect 56926 7410 56978 7422
rect 3950 7362 4002 7374
rect 3950 7298 4002 7310
rect 5518 7362 5570 7374
rect 5518 7298 5570 7310
rect 6750 7362 6802 7374
rect 6750 7298 6802 7310
rect 7310 7362 7362 7374
rect 7310 7298 7362 7310
rect 7758 7362 7810 7374
rect 7758 7298 7810 7310
rect 9102 7362 9154 7374
rect 14478 7362 14530 7374
rect 12450 7310 12462 7362
rect 12514 7310 12526 7362
rect 13234 7310 13246 7362
rect 13298 7310 13310 7362
rect 9102 7298 9154 7310
rect 14478 7298 14530 7310
rect 15934 7362 15986 7374
rect 19854 7362 19906 7374
rect 25790 7362 25842 7374
rect 32286 7362 32338 7374
rect 16706 7310 16718 7362
rect 16770 7310 16782 7362
rect 18386 7310 18398 7362
rect 18450 7310 18462 7362
rect 20850 7310 20862 7362
rect 20914 7310 20926 7362
rect 29138 7310 29150 7362
rect 29202 7310 29214 7362
rect 15934 7298 15986 7310
rect 19854 7298 19906 7310
rect 25790 7298 25842 7310
rect 32286 7298 32338 7310
rect 33854 7362 33906 7374
rect 33854 7298 33906 7310
rect 34974 7362 35026 7374
rect 44382 7362 44434 7374
rect 56814 7362 56866 7374
rect 42802 7310 42814 7362
rect 42866 7310 42878 7362
rect 46162 7310 46174 7362
rect 46226 7310 46238 7362
rect 49186 7310 49198 7362
rect 49250 7310 49262 7362
rect 51426 7310 51438 7362
rect 51490 7310 51502 7362
rect 34974 7298 35026 7310
rect 44382 7298 44434 7310
rect 56814 7298 56866 7310
rect 14702 7250 14754 7262
rect 15710 7250 15762 7262
rect 30830 7250 30882 7262
rect 15362 7198 15374 7250
rect 15426 7198 15438 7250
rect 23202 7198 23214 7250
rect 23266 7198 23278 7250
rect 14702 7186 14754 7198
rect 15710 7186 15762 7198
rect 30830 7186 30882 7198
rect 38670 7250 38722 7262
rect 50878 7250 50930 7262
rect 49522 7198 49534 7250
rect 49586 7198 49598 7250
rect 53106 7198 53118 7250
rect 53170 7198 53182 7250
rect 38670 7186 38722 7198
rect 50878 7186 50930 7198
rect 1344 7082 58576 7116
rect 1344 7030 8367 7082
rect 8419 7030 8471 7082
rect 8523 7030 8575 7082
rect 8627 7030 22674 7082
rect 22726 7030 22778 7082
rect 22830 7030 22882 7082
rect 22934 7030 36981 7082
rect 37033 7030 37085 7082
rect 37137 7030 37189 7082
rect 37241 7030 51288 7082
rect 51340 7030 51392 7082
rect 51444 7030 51496 7082
rect 51548 7030 58576 7082
rect 1344 6996 58576 7030
rect 19966 6914 20018 6926
rect 19966 6850 20018 6862
rect 20190 6914 20242 6926
rect 20190 6850 20242 6862
rect 20638 6914 20690 6926
rect 20638 6850 20690 6862
rect 28254 6914 28306 6926
rect 36318 6914 36370 6926
rect 58046 6914 58098 6926
rect 35410 6862 35422 6914
rect 35474 6862 35486 6914
rect 39778 6862 39790 6914
rect 39842 6862 39854 6914
rect 49298 6862 49310 6914
rect 49362 6862 49374 6914
rect 50866 6862 50878 6914
rect 50930 6911 50942 6914
rect 51874 6911 51886 6914
rect 50930 6865 51886 6911
rect 50930 6862 50942 6865
rect 51874 6862 51886 6865
rect 51938 6862 51950 6914
rect 28254 6850 28306 6862
rect 36318 6850 36370 6862
rect 58046 6850 58098 6862
rect 23102 6802 23154 6814
rect 35086 6802 35138 6814
rect 2594 6750 2606 6802
rect 2658 6750 2670 6802
rect 4722 6750 4734 6802
rect 4786 6750 4798 6802
rect 6402 6750 6414 6802
rect 6466 6750 6478 6802
rect 14354 6750 14366 6802
rect 14418 6750 14430 6802
rect 28578 6750 28590 6802
rect 28642 6750 28654 6802
rect 23102 6738 23154 6750
rect 35086 6738 35138 6750
rect 35982 6802 36034 6814
rect 50094 6802 50146 6814
rect 55806 6802 55858 6814
rect 43026 6750 43038 6802
rect 43090 6750 43102 6802
rect 45938 6750 45950 6802
rect 46002 6750 46014 6802
rect 49522 6750 49534 6802
rect 49586 6750 49598 6802
rect 50418 6750 50430 6802
rect 50482 6750 50494 6802
rect 57250 6750 57262 6802
rect 57314 6750 57326 6802
rect 35982 6738 36034 6750
rect 50094 6738 50146 6750
rect 55806 6738 55858 6750
rect 7534 6690 7586 6702
rect 12126 6690 12178 6702
rect 1922 6638 1934 6690
rect 1986 6638 1998 6690
rect 5730 6638 5742 6690
rect 5794 6638 5806 6690
rect 6290 6638 6302 6690
rect 6354 6638 6366 6690
rect 7858 6638 7870 6690
rect 7922 6638 7934 6690
rect 8530 6638 8542 6690
rect 8594 6638 8606 6690
rect 7534 6626 7586 6638
rect 12126 6626 12178 6638
rect 12238 6690 12290 6702
rect 12238 6626 12290 6638
rect 12574 6690 12626 6702
rect 12574 6626 12626 6638
rect 13470 6690 13522 6702
rect 15486 6690 15538 6702
rect 20526 6690 20578 6702
rect 14018 6638 14030 6690
rect 14082 6638 14094 6690
rect 16258 6638 16270 6690
rect 16322 6638 16334 6690
rect 16818 6638 16830 6690
rect 16882 6638 16894 6690
rect 18610 6638 18622 6690
rect 18674 6638 18686 6690
rect 19058 6638 19070 6690
rect 19122 6638 19134 6690
rect 13470 6626 13522 6638
rect 15486 6626 15538 6638
rect 20526 6626 20578 6638
rect 22766 6690 22818 6702
rect 28030 6690 28082 6702
rect 26114 6638 26126 6690
rect 26178 6638 26190 6690
rect 26674 6638 26686 6690
rect 26738 6638 26750 6690
rect 22766 6626 22818 6638
rect 28030 6626 28082 6638
rect 31054 6690 31106 6702
rect 31054 6626 31106 6638
rect 31278 6690 31330 6702
rect 31278 6626 31330 6638
rect 32622 6690 32674 6702
rect 33966 6690 34018 6702
rect 33394 6638 33406 6690
rect 33458 6638 33470 6690
rect 32622 6626 32674 6638
rect 33966 6626 34018 6638
rect 34302 6690 34354 6702
rect 34302 6626 34354 6638
rect 34862 6690 34914 6702
rect 34862 6626 34914 6638
rect 35758 6690 35810 6702
rect 38894 6690 38946 6702
rect 44046 6690 44098 6702
rect 38546 6638 38558 6690
rect 38610 6638 38622 6690
rect 39890 6638 39902 6690
rect 39954 6638 39966 6690
rect 42354 6638 42366 6690
rect 42418 6638 42430 6690
rect 43586 6638 43598 6690
rect 43650 6638 43662 6690
rect 35758 6626 35810 6638
rect 38894 6626 38946 6638
rect 44046 6626 44098 6638
rect 44158 6690 44210 6702
rect 47742 6690 47794 6702
rect 51774 6690 51826 6702
rect 53566 6690 53618 6702
rect 45826 6638 45838 6690
rect 45890 6638 45902 6690
rect 46946 6638 46958 6690
rect 47010 6638 47022 6690
rect 48850 6638 48862 6690
rect 48914 6638 48926 6690
rect 52994 6638 53006 6690
rect 53058 6638 53070 6690
rect 44158 6626 44210 6638
rect 47742 6626 47794 6638
rect 51774 6626 51826 6638
rect 53566 6626 53618 6638
rect 54014 6690 54066 6702
rect 54014 6626 54066 6638
rect 54350 6690 54402 6702
rect 58158 6690 58210 6702
rect 57138 6638 57150 6690
rect 57202 6638 57214 6690
rect 54350 6626 54402 6638
rect 58158 6626 58210 6638
rect 20750 6578 20802 6590
rect 6514 6526 6526 6578
rect 6578 6526 6590 6578
rect 17490 6526 17502 6578
rect 17554 6526 17566 6578
rect 17826 6526 17838 6578
rect 17890 6526 17902 6578
rect 20750 6514 20802 6526
rect 21870 6578 21922 6590
rect 28478 6578 28530 6590
rect 30830 6578 30882 6590
rect 25218 6526 25230 6578
rect 25282 6526 25294 6578
rect 27346 6526 27358 6578
rect 27410 6526 27422 6578
rect 29138 6526 29150 6578
rect 29202 6526 29214 6578
rect 21870 6514 21922 6526
rect 28478 6514 28530 6526
rect 30830 6514 30882 6526
rect 31166 6578 31218 6590
rect 31166 6514 31218 6526
rect 31614 6578 31666 6590
rect 31614 6514 31666 6526
rect 31950 6578 32002 6590
rect 31950 6514 32002 6526
rect 32286 6578 32338 6590
rect 32286 6514 32338 6526
rect 32398 6578 32450 6590
rect 37550 6578 37602 6590
rect 47854 6578 47906 6590
rect 32834 6526 32846 6578
rect 32898 6526 32910 6578
rect 33282 6526 33294 6578
rect 33346 6526 33358 6578
rect 41682 6526 41694 6578
rect 41746 6526 41758 6578
rect 43698 6526 43710 6578
rect 43762 6526 43774 6578
rect 45714 6526 45726 6578
rect 45778 6526 45790 6578
rect 32398 6514 32450 6526
rect 37550 6514 37602 6526
rect 47854 6514 47906 6526
rect 50318 6578 50370 6590
rect 50318 6514 50370 6526
rect 50878 6578 50930 6590
rect 50878 6514 50930 6526
rect 51326 6578 51378 6590
rect 51326 6514 51378 6526
rect 53678 6578 53730 6590
rect 53678 6514 53730 6526
rect 57598 6578 57650 6590
rect 57598 6514 57650 6526
rect 11342 6466 11394 6478
rect 10770 6414 10782 6466
rect 10834 6414 10846 6466
rect 11342 6402 11394 6414
rect 11902 6466 11954 6478
rect 15150 6466 15202 6478
rect 29710 6466 29762 6478
rect 12898 6414 12910 6466
rect 12962 6414 12974 6466
rect 23314 6414 23326 6466
rect 23378 6414 23390 6466
rect 24322 6414 24334 6466
rect 24386 6414 24398 6466
rect 11902 6402 11954 6414
rect 15150 6402 15202 6414
rect 29710 6402 29762 6414
rect 34078 6466 34130 6478
rect 34078 6402 34130 6414
rect 37662 6466 37714 6478
rect 42142 6466 42194 6478
rect 40786 6414 40798 6466
rect 40850 6414 40862 6466
rect 37662 6402 37714 6414
rect 42142 6402 42194 6414
rect 48078 6466 48130 6478
rect 48078 6402 48130 6414
rect 54126 6466 54178 6478
rect 54126 6402 54178 6414
rect 55694 6466 55746 6478
rect 55694 6402 55746 6414
rect 55918 6466 55970 6478
rect 55918 6402 55970 6414
rect 56142 6466 56194 6478
rect 56142 6402 56194 6414
rect 58046 6466 58098 6478
rect 58046 6402 58098 6414
rect 1344 6298 58731 6332
rect 1344 6246 15520 6298
rect 15572 6246 15624 6298
rect 15676 6246 15728 6298
rect 15780 6246 29827 6298
rect 29879 6246 29931 6298
rect 29983 6246 30035 6298
rect 30087 6246 44134 6298
rect 44186 6246 44238 6298
rect 44290 6246 44342 6298
rect 44394 6246 58441 6298
rect 58493 6246 58545 6298
rect 58597 6246 58649 6298
rect 58701 6246 58731 6298
rect 1344 6212 58731 6246
rect 1934 6130 1986 6142
rect 1934 6066 1986 6078
rect 2494 6130 2546 6142
rect 8990 6130 9042 6142
rect 4722 6078 4734 6130
rect 4786 6078 4798 6130
rect 5282 6078 5294 6130
rect 5346 6078 5358 6130
rect 8194 6078 8206 6130
rect 8258 6078 8270 6130
rect 2494 6066 2546 6078
rect 8990 6066 9042 6078
rect 9774 6130 9826 6142
rect 9774 6066 9826 6078
rect 10222 6130 10274 6142
rect 10222 6066 10274 6078
rect 13918 6130 13970 6142
rect 14814 6130 14866 6142
rect 24670 6130 24722 6142
rect 14466 6078 14478 6130
rect 14530 6078 14542 6130
rect 22754 6078 22766 6130
rect 22818 6078 22830 6130
rect 13918 6066 13970 6078
rect 14814 6066 14866 6078
rect 24670 6066 24722 6078
rect 27246 6130 27298 6142
rect 33182 6130 33234 6142
rect 32386 6078 32398 6130
rect 32450 6078 32462 6130
rect 27246 6066 27298 6078
rect 33182 6066 33234 6078
rect 34750 6130 34802 6142
rect 34750 6066 34802 6078
rect 38110 6130 38162 6142
rect 38110 6066 38162 6078
rect 38222 6130 38274 6142
rect 38222 6066 38274 6078
rect 39006 6130 39058 6142
rect 54126 6130 54178 6142
rect 53554 6078 53566 6130
rect 53618 6078 53630 6130
rect 39006 6066 39058 6078
rect 54126 6066 54178 6078
rect 57822 6130 57874 6142
rect 57822 6066 57874 6078
rect 8654 6018 8706 6030
rect 3266 5966 3278 6018
rect 3330 5966 3342 6018
rect 4610 5966 4622 6018
rect 4674 5966 4686 6018
rect 6626 5966 6638 6018
rect 6690 5966 6702 6018
rect 8654 5954 8706 5966
rect 10446 6018 10498 6030
rect 10446 5954 10498 5966
rect 10782 6018 10834 6030
rect 10782 5954 10834 5966
rect 11118 6018 11170 6030
rect 11118 5954 11170 5966
rect 11230 6018 11282 6030
rect 11230 5954 11282 5966
rect 11902 6018 11954 6030
rect 11902 5954 11954 5966
rect 12238 6018 12290 6030
rect 12238 5954 12290 5966
rect 12350 6018 12402 6030
rect 12350 5954 12402 5966
rect 13022 6018 13074 6030
rect 21646 6018 21698 6030
rect 19842 5966 19854 6018
rect 19906 5966 19918 6018
rect 13022 5954 13074 5966
rect 21646 5954 21698 5966
rect 23662 6018 23714 6030
rect 33966 6018 34018 6030
rect 37326 6018 37378 6030
rect 25218 5966 25230 6018
rect 25282 5966 25294 6018
rect 27794 5966 27806 6018
rect 27858 5966 27870 6018
rect 28802 5966 28814 6018
rect 28866 5966 28878 6018
rect 31826 5966 31838 6018
rect 31890 5966 31902 6018
rect 34178 5966 34190 6018
rect 34242 5966 34254 6018
rect 23662 5954 23714 5966
rect 33966 5954 34018 5966
rect 37326 5954 37378 5966
rect 38670 6018 38722 6030
rect 50990 6018 51042 6030
rect 54014 6018 54066 6030
rect 41234 5966 41246 6018
rect 41298 5966 41310 6018
rect 43586 5966 43598 6018
rect 43650 5966 43662 6018
rect 51874 5966 51886 6018
rect 51938 5966 51950 6018
rect 38670 5954 38722 5966
rect 50990 5954 51042 5966
rect 54014 5954 54066 5966
rect 54686 6018 54738 6030
rect 54686 5954 54738 5966
rect 54798 6018 54850 6030
rect 54798 5954 54850 5966
rect 55806 6018 55858 6030
rect 55806 5954 55858 5966
rect 58046 6018 58098 6030
rect 58046 5954 58098 5966
rect 6302 5906 6354 5918
rect 12574 5906 12626 5918
rect 3602 5854 3614 5906
rect 3666 5854 3678 5906
rect 5506 5854 5518 5906
rect 5570 5854 5582 5906
rect 5954 5854 5966 5906
rect 6018 5854 6030 5906
rect 7746 5854 7758 5906
rect 7810 5854 7822 5906
rect 6302 5842 6354 5854
rect 12574 5842 12626 5854
rect 12798 5906 12850 5918
rect 12798 5842 12850 5854
rect 13358 5906 13410 5918
rect 13358 5842 13410 5854
rect 13806 5906 13858 5918
rect 13806 5842 13858 5854
rect 14030 5906 14082 5918
rect 22094 5906 22146 5918
rect 15810 5854 15822 5906
rect 15874 5854 15886 5906
rect 16146 5854 16158 5906
rect 16210 5854 16222 5906
rect 17826 5854 17838 5906
rect 17890 5854 17902 5906
rect 18946 5854 18958 5906
rect 19010 5854 19022 5906
rect 14030 5842 14082 5854
rect 22094 5842 22146 5854
rect 22542 5906 22594 5918
rect 27470 5906 27522 5918
rect 32958 5906 33010 5918
rect 25330 5854 25342 5906
rect 25394 5854 25406 5906
rect 26002 5854 26014 5906
rect 26066 5854 26078 5906
rect 26562 5854 26574 5906
rect 26626 5854 26638 5906
rect 28914 5854 28926 5906
rect 28978 5854 28990 5906
rect 29698 5854 29710 5906
rect 29762 5854 29774 5906
rect 31378 5854 31390 5906
rect 31442 5854 31454 5906
rect 32274 5854 32286 5906
rect 32338 5854 32350 5906
rect 22542 5842 22594 5854
rect 27470 5842 27522 5854
rect 32958 5842 33010 5854
rect 33294 5906 33346 5918
rect 33294 5842 33346 5854
rect 33854 5906 33906 5918
rect 40238 5906 40290 5918
rect 46286 5906 46338 5918
rect 47182 5906 47234 5918
rect 34290 5854 34302 5906
rect 34354 5854 34366 5906
rect 35522 5854 35534 5906
rect 35586 5854 35598 5906
rect 36530 5854 36542 5906
rect 36594 5854 36606 5906
rect 39778 5854 39790 5906
rect 39842 5854 39854 5906
rect 42466 5854 42478 5906
rect 42530 5854 42542 5906
rect 44258 5854 44270 5906
rect 44322 5854 44334 5906
rect 44706 5854 44718 5906
rect 44770 5854 44782 5906
rect 46498 5854 46510 5906
rect 46562 5854 46574 5906
rect 33854 5842 33906 5854
rect 40238 5842 40290 5854
rect 46286 5842 46338 5854
rect 47182 5842 47234 5854
rect 47630 5906 47682 5918
rect 47630 5842 47682 5854
rect 48862 5906 48914 5918
rect 54462 5906 54514 5918
rect 49298 5854 49310 5906
rect 49362 5854 49374 5906
rect 50418 5854 50430 5906
rect 50482 5854 50494 5906
rect 53218 5854 53230 5906
rect 53282 5854 53294 5906
rect 48862 5842 48914 5854
rect 54462 5842 54514 5854
rect 56030 5906 56082 5918
rect 56030 5842 56082 5854
rect 56590 5906 56642 5918
rect 57486 5906 57538 5918
rect 57026 5854 57038 5906
rect 57090 5854 57102 5906
rect 56590 5842 56642 5854
rect 57486 5842 57538 5854
rect 58158 5906 58210 5918
rect 58158 5842 58210 5854
rect 47854 5794 47906 5806
rect 13122 5742 13134 5794
rect 13186 5742 13198 5794
rect 16706 5742 16718 5794
rect 16770 5742 16782 5794
rect 18274 5742 18286 5794
rect 18338 5742 18350 5794
rect 31042 5742 31054 5794
rect 31106 5742 31118 5794
rect 35074 5742 35086 5794
rect 35138 5742 35150 5794
rect 41010 5742 41022 5794
rect 41074 5742 41086 5794
rect 45826 5742 45838 5794
rect 45890 5742 45902 5794
rect 47854 5730 47906 5742
rect 49758 5794 49810 5806
rect 49758 5730 49810 5742
rect 50094 5794 50146 5806
rect 50094 5730 50146 5742
rect 50206 5794 50258 5806
rect 50206 5730 50258 5742
rect 50878 5794 50930 5806
rect 50878 5730 50930 5742
rect 51662 5794 51714 5806
rect 55682 5742 55694 5794
rect 55746 5742 55758 5794
rect 51662 5730 51714 5742
rect 5966 5682 6018 5694
rect 5966 5618 6018 5630
rect 11230 5682 11282 5694
rect 38334 5682 38386 5694
rect 50766 5682 50818 5694
rect 26338 5630 26350 5682
rect 26402 5630 26414 5682
rect 48178 5630 48190 5682
rect 48242 5630 48254 5682
rect 11230 5618 11282 5630
rect 38334 5618 38386 5630
rect 50766 5618 50818 5630
rect 54126 5682 54178 5694
rect 54126 5618 54178 5630
rect 1344 5514 58576 5548
rect 1344 5462 8367 5514
rect 8419 5462 8471 5514
rect 8523 5462 8575 5514
rect 8627 5462 22674 5514
rect 22726 5462 22778 5514
rect 22830 5462 22882 5514
rect 22934 5462 36981 5514
rect 37033 5462 37085 5514
rect 37137 5462 37189 5514
rect 37241 5462 51288 5514
rect 51340 5462 51392 5514
rect 51444 5462 51496 5514
rect 51548 5462 58576 5514
rect 1344 5428 58576 5462
rect 5070 5346 5122 5358
rect 5070 5282 5122 5294
rect 9102 5346 9154 5358
rect 9102 5282 9154 5294
rect 12910 5346 12962 5358
rect 26798 5346 26850 5358
rect 26226 5294 26238 5346
rect 26290 5294 26302 5346
rect 12910 5282 12962 5294
rect 26798 5282 26850 5294
rect 29262 5346 29314 5358
rect 29262 5282 29314 5294
rect 29598 5346 29650 5358
rect 29598 5282 29650 5294
rect 30606 5346 30658 5358
rect 30606 5282 30658 5294
rect 32622 5346 32674 5358
rect 32622 5282 32674 5294
rect 41134 5346 41186 5358
rect 41134 5282 41186 5294
rect 47966 5346 48018 5358
rect 47966 5282 48018 5294
rect 48974 5346 49026 5358
rect 48974 5282 49026 5294
rect 49422 5346 49474 5358
rect 49422 5282 49474 5294
rect 49758 5346 49810 5358
rect 49758 5282 49810 5294
rect 51102 5346 51154 5358
rect 55234 5294 55246 5346
rect 55298 5294 55310 5346
rect 51102 5282 51154 5294
rect 3502 5234 3554 5246
rect 3502 5170 3554 5182
rect 4958 5234 5010 5246
rect 4958 5170 5010 5182
rect 5854 5234 5906 5246
rect 8878 5234 8930 5246
rect 8194 5182 8206 5234
rect 8258 5182 8270 5234
rect 5854 5170 5906 5182
rect 8878 5170 8930 5182
rect 9214 5234 9266 5246
rect 12014 5234 12066 5246
rect 9874 5182 9886 5234
rect 9938 5182 9950 5234
rect 9214 5170 9266 5182
rect 12014 5170 12066 5182
rect 12462 5234 12514 5246
rect 12462 5170 12514 5182
rect 15486 5234 15538 5246
rect 20302 5234 20354 5246
rect 25678 5234 25730 5246
rect 35086 5234 35138 5246
rect 17042 5182 17054 5234
rect 17106 5182 17118 5234
rect 23314 5182 23326 5234
rect 23378 5182 23390 5234
rect 25330 5182 25342 5234
rect 25394 5182 25406 5234
rect 30146 5182 30158 5234
rect 30210 5182 30222 5234
rect 31714 5182 31726 5234
rect 31778 5182 31790 5234
rect 33506 5182 33518 5234
rect 33570 5182 33582 5234
rect 34514 5182 34526 5234
rect 34578 5182 34590 5234
rect 15486 5170 15538 5182
rect 20302 5170 20354 5182
rect 25678 5170 25730 5182
rect 35086 5170 35138 5182
rect 35534 5234 35586 5246
rect 35534 5170 35586 5182
rect 35758 5234 35810 5246
rect 43486 5234 43538 5246
rect 37090 5182 37102 5234
rect 37154 5182 37166 5234
rect 43698 5182 43710 5234
rect 43762 5182 43774 5234
rect 53442 5182 53454 5234
rect 53506 5182 53518 5234
rect 35758 5170 35810 5182
rect 43486 5170 43538 5182
rect 9550 5122 9602 5134
rect 6626 5070 6638 5122
rect 6690 5070 6702 5122
rect 9550 5058 9602 5070
rect 10446 5122 10498 5134
rect 10446 5058 10498 5070
rect 10670 5122 10722 5134
rect 10670 5058 10722 5070
rect 10782 5122 10834 5134
rect 10782 5058 10834 5070
rect 11006 5122 11058 5134
rect 17390 5122 17442 5134
rect 25902 5122 25954 5134
rect 29374 5122 29426 5134
rect 32286 5122 32338 5134
rect 16706 5070 16718 5122
rect 16770 5070 16782 5122
rect 18274 5070 18286 5122
rect 18338 5070 18350 5122
rect 19170 5070 19182 5122
rect 19234 5070 19246 5122
rect 19506 5070 19518 5122
rect 19570 5070 19582 5122
rect 22306 5070 22318 5122
rect 22370 5070 22382 5122
rect 22642 5070 22654 5122
rect 22706 5070 22718 5122
rect 23762 5070 23774 5122
rect 23826 5070 23838 5122
rect 24210 5070 24222 5122
rect 24274 5070 24286 5122
rect 27570 5070 27582 5122
rect 27634 5070 27646 5122
rect 28354 5070 28366 5122
rect 28418 5070 28430 5122
rect 31266 5070 31278 5122
rect 31330 5070 31342 5122
rect 31490 5070 31502 5122
rect 31554 5070 31566 5122
rect 11006 5058 11058 5070
rect 17390 5058 17442 5070
rect 25902 5058 25954 5070
rect 29374 5058 29426 5070
rect 32286 5058 32338 5070
rect 32510 5122 32562 5134
rect 32510 5058 32562 5070
rect 33070 5122 33122 5134
rect 34414 5122 34466 5134
rect 40686 5122 40738 5134
rect 44830 5122 44882 5134
rect 33954 5070 33966 5122
rect 34018 5070 34030 5122
rect 38770 5070 38782 5122
rect 38834 5070 38846 5122
rect 39890 5070 39902 5122
rect 39954 5070 39966 5122
rect 41906 5070 41918 5122
rect 41970 5070 41982 5122
rect 33070 5058 33122 5070
rect 34414 5058 34466 5070
rect 40686 5058 40738 5070
rect 44830 5058 44882 5070
rect 46622 5122 46674 5134
rect 48750 5122 48802 5134
rect 51438 5122 51490 5134
rect 48514 5070 48526 5122
rect 48578 5070 48590 5122
rect 49746 5070 49758 5122
rect 49810 5070 49822 5122
rect 46622 5058 46674 5070
rect 48750 5058 48802 5070
rect 51438 5058 51490 5070
rect 51662 5122 51714 5134
rect 51662 5058 51714 5070
rect 51774 5122 51826 5134
rect 51774 5058 51826 5070
rect 51998 5122 52050 5134
rect 54014 5122 54066 5134
rect 53106 5070 53118 5122
rect 53170 5070 53182 5122
rect 51998 5058 52050 5070
rect 54014 5058 54066 5070
rect 54350 5122 54402 5134
rect 56590 5122 56642 5134
rect 55906 5070 55918 5122
rect 55970 5070 55982 5122
rect 56914 5070 56926 5122
rect 56978 5070 56990 5122
rect 54350 5058 54402 5070
rect 56590 5058 56642 5070
rect 4846 5010 4898 5022
rect 9774 5010 9826 5022
rect 7858 4958 7870 5010
rect 7922 4958 7934 5010
rect 4846 4946 4898 4958
rect 9774 4946 9826 4958
rect 10222 5010 10274 5022
rect 10222 4946 10274 4958
rect 11342 5010 11394 5022
rect 11342 4946 11394 4958
rect 12798 5010 12850 5022
rect 28590 5010 28642 5022
rect 13682 4958 13694 5010
rect 13746 4958 13758 5010
rect 15138 4958 15150 5010
rect 15202 4958 15214 5010
rect 16482 4958 16494 5010
rect 16546 4958 16558 5010
rect 12798 4946 12850 4958
rect 28590 4946 28642 4958
rect 30494 5010 30546 5022
rect 39230 5010 39282 5022
rect 40350 5010 40402 5022
rect 37538 4958 37550 5010
rect 37602 4958 37614 5010
rect 39666 4958 39678 5010
rect 39730 4958 39742 5010
rect 30494 4946 30546 4958
rect 39230 4946 39282 4958
rect 40350 4946 40402 4958
rect 41022 5010 41074 5022
rect 41022 4946 41074 4958
rect 41134 5010 41186 5022
rect 41134 4946 41186 4958
rect 41694 5010 41746 5022
rect 49086 5010 49138 5022
rect 42354 4958 42366 5010
rect 42418 4958 42430 5010
rect 47170 4958 47182 5010
rect 47234 4958 47246 5010
rect 41694 4946 41746 4958
rect 49086 4946 49138 4958
rect 51102 5010 51154 5022
rect 51102 4946 51154 4958
rect 51214 5010 51266 5022
rect 51214 4946 51266 4958
rect 52670 5010 52722 5022
rect 52670 4946 52722 4958
rect 54238 5010 54290 5022
rect 54238 4946 54290 4958
rect 3950 4898 4002 4910
rect 3950 4834 4002 4846
rect 4398 4898 4450 4910
rect 11230 4898 11282 4910
rect 32622 4898 32674 4910
rect 6402 4846 6414 4898
rect 6466 4846 6478 4898
rect 13570 4846 13582 4898
rect 13634 4846 13646 4898
rect 4398 4834 4450 4846
rect 11230 4834 11282 4846
rect 32622 4834 32674 4846
rect 34190 4898 34242 4910
rect 34190 4834 34242 4846
rect 34526 4898 34578 4910
rect 42702 4898 42754 4910
rect 36082 4846 36094 4898
rect 36146 4846 36158 4898
rect 34526 4834 34578 4846
rect 42702 4834 42754 4846
rect 43710 4898 43762 4910
rect 43710 4834 43762 4846
rect 45166 4898 45218 4910
rect 45166 4834 45218 4846
rect 1344 4730 58731 4764
rect 1344 4678 15520 4730
rect 15572 4678 15624 4730
rect 15676 4678 15728 4730
rect 15780 4678 29827 4730
rect 29879 4678 29931 4730
rect 29983 4678 30035 4730
rect 30087 4678 44134 4730
rect 44186 4678 44238 4730
rect 44290 4678 44342 4730
rect 44394 4678 58441 4730
rect 58493 4678 58545 4730
rect 58597 4678 58649 4730
rect 58701 4678 58731 4730
rect 1344 4644 58731 4678
rect 8990 4562 9042 4574
rect 8990 4498 9042 4510
rect 10110 4562 10162 4574
rect 10110 4498 10162 4510
rect 11342 4562 11394 4574
rect 11342 4498 11394 4510
rect 15934 4562 15986 4574
rect 15934 4498 15986 4510
rect 17726 4562 17778 4574
rect 17726 4498 17778 4510
rect 24334 4562 24386 4574
rect 24334 4498 24386 4510
rect 25454 4562 25506 4574
rect 34078 4562 34130 4574
rect 33618 4510 33630 4562
rect 33682 4510 33694 4562
rect 25454 4498 25506 4510
rect 34078 4498 34130 4510
rect 35086 4562 35138 4574
rect 35086 4498 35138 4510
rect 40238 4562 40290 4574
rect 40238 4498 40290 4510
rect 46734 4562 46786 4574
rect 46734 4498 46786 4510
rect 8094 4450 8146 4462
rect 8094 4386 8146 4398
rect 8430 4450 8482 4462
rect 8430 4386 8482 4398
rect 9886 4450 9938 4462
rect 9886 4386 9938 4398
rect 10894 4450 10946 4462
rect 10894 4386 10946 4398
rect 12126 4450 12178 4462
rect 12126 4386 12178 4398
rect 12910 4450 12962 4462
rect 14702 4450 14754 4462
rect 14018 4398 14030 4450
rect 14082 4398 14094 4450
rect 12910 4386 12962 4398
rect 14702 4386 14754 4398
rect 15038 4450 15090 4462
rect 24670 4450 24722 4462
rect 33854 4450 33906 4462
rect 40126 4450 40178 4462
rect 18498 4398 18510 4450
rect 18562 4398 18574 4450
rect 20402 4398 20414 4450
rect 20466 4398 20478 4450
rect 20962 4398 20974 4450
rect 21026 4398 21038 4450
rect 23986 4398 23998 4450
rect 24050 4398 24062 4450
rect 27122 4398 27134 4450
rect 27186 4398 27198 4450
rect 28802 4398 28814 4450
rect 28866 4398 28878 4450
rect 29474 4398 29486 4450
rect 29538 4398 29550 4450
rect 30594 4398 30606 4450
rect 30658 4398 30670 4450
rect 38882 4398 38894 4450
rect 38946 4398 38958 4450
rect 15038 4386 15090 4398
rect 24670 4386 24722 4398
rect 33854 4386 33906 4398
rect 40126 4386 40178 4398
rect 43262 4450 43314 4462
rect 51998 4450 52050 4462
rect 44594 4398 44606 4450
rect 44658 4398 44670 4450
rect 43262 4386 43314 4398
rect 51998 4386 52050 4398
rect 52222 4450 52274 4462
rect 52222 4386 52274 4398
rect 7646 4338 7698 4350
rect 4386 4286 4398 4338
rect 4450 4286 4462 4338
rect 7646 4274 7698 4286
rect 10558 4338 10610 4350
rect 10558 4274 10610 4286
rect 11454 4338 11506 4350
rect 11454 4274 11506 4286
rect 11902 4338 11954 4350
rect 15374 4338 15426 4350
rect 29822 4338 29874 4350
rect 33294 4338 33346 4350
rect 12674 4286 12686 4338
rect 12738 4286 12750 4338
rect 13234 4286 13246 4338
rect 13298 4286 13310 4338
rect 13794 4286 13806 4338
rect 13858 4286 13870 4338
rect 16706 4286 16718 4338
rect 16770 4286 16782 4338
rect 17490 4286 17502 4338
rect 17554 4286 17566 4338
rect 18050 4286 18062 4338
rect 18114 4286 18126 4338
rect 19394 4286 19406 4338
rect 19458 4286 19470 4338
rect 20850 4286 20862 4338
rect 20914 4286 20926 4338
rect 21970 4286 21982 4338
rect 22034 4286 22046 4338
rect 22754 4286 22766 4338
rect 22818 4286 22830 4338
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 26226 4286 26238 4338
rect 26290 4286 26302 4338
rect 26562 4286 26574 4338
rect 26626 4286 26638 4338
rect 27794 4286 27806 4338
rect 27858 4286 27870 4338
rect 28914 4286 28926 4338
rect 28978 4286 28990 4338
rect 30930 4286 30942 4338
rect 30994 4286 31006 4338
rect 31938 4286 31950 4338
rect 32002 4286 32014 4338
rect 11902 4274 11954 4286
rect 15374 4274 15426 4286
rect 29822 4274 29874 4286
rect 33294 4274 33346 4286
rect 34190 4338 34242 4350
rect 40462 4338 40514 4350
rect 47406 4338 47458 4350
rect 38210 4286 38222 4338
rect 38274 4286 38286 4338
rect 39330 4286 39342 4338
rect 39394 4286 39406 4338
rect 41122 4286 41134 4338
rect 41186 4286 41198 4338
rect 42466 4286 42478 4338
rect 42530 4286 42542 4338
rect 45378 4286 45390 4338
rect 45442 4286 45454 4338
rect 34190 4274 34242 4286
rect 40462 4274 40514 4286
rect 47406 4274 47458 4286
rect 8878 4226 8930 4238
rect 16270 4226 16322 4238
rect 25566 4226 25618 4238
rect 28478 4226 28530 4238
rect 5058 4174 5070 4226
rect 5122 4174 5134 4226
rect 7186 4174 7198 4226
rect 7250 4174 7262 4226
rect 10210 4174 10222 4226
rect 10274 4174 10286 4226
rect 13682 4174 13694 4226
rect 13746 4174 13758 4226
rect 20962 4174 20974 4226
rect 21026 4174 21038 4226
rect 22866 4174 22878 4226
rect 22930 4174 22942 4226
rect 26674 4174 26686 4226
rect 26738 4174 26750 4226
rect 27570 4174 27582 4226
rect 27634 4174 27646 4226
rect 8878 4162 8930 4174
rect 16270 4162 16322 4174
rect 25566 4162 25618 4174
rect 28478 4162 28530 4174
rect 29934 4226 29986 4238
rect 29934 4162 29986 4174
rect 32510 4226 32562 4238
rect 32510 4162 32562 4174
rect 34638 4226 34690 4238
rect 34638 4162 34690 4174
rect 37886 4226 37938 4238
rect 47070 4226 47122 4238
rect 39106 4174 39118 4226
rect 39170 4174 39182 4226
rect 41458 4174 41470 4226
rect 41522 4174 41534 4226
rect 43922 4174 43934 4226
rect 43986 4174 43998 4226
rect 47842 4174 47854 4226
rect 47906 4174 47918 4226
rect 51874 4174 51886 4226
rect 51938 4174 51950 4226
rect 37886 4162 37938 4174
rect 47070 4162 47122 4174
rect 7758 4114 7810 4126
rect 7758 4050 7810 4062
rect 11566 4114 11618 4126
rect 11566 4050 11618 4062
rect 12238 4114 12290 4126
rect 12238 4050 12290 4062
rect 1344 3946 58576 3980
rect 1344 3894 8367 3946
rect 8419 3894 8471 3946
rect 8523 3894 8575 3946
rect 8627 3894 22674 3946
rect 22726 3894 22778 3946
rect 22830 3894 22882 3946
rect 22934 3894 36981 3946
rect 37033 3894 37085 3946
rect 37137 3894 37189 3946
rect 37241 3894 51288 3946
rect 51340 3894 51392 3946
rect 51444 3894 51496 3946
rect 51548 3894 58576 3946
rect 1344 3860 58576 3894
rect 16046 3778 16098 3790
rect 28590 3778 28642 3790
rect 29710 3778 29762 3790
rect 40798 3778 40850 3790
rect 16370 3726 16382 3778
rect 16434 3726 16446 3778
rect 28914 3726 28926 3778
rect 28978 3726 28990 3778
rect 29362 3726 29374 3778
rect 29426 3726 29438 3778
rect 38098 3726 38110 3778
rect 38162 3726 38174 3778
rect 16046 3714 16098 3726
rect 28590 3714 28642 3726
rect 29710 3714 29762 3726
rect 40798 3714 40850 3726
rect 6302 3666 6354 3678
rect 6302 3602 6354 3614
rect 6750 3666 6802 3678
rect 6750 3602 6802 3614
rect 7198 3666 7250 3678
rect 7198 3602 7250 3614
rect 7646 3666 7698 3678
rect 15822 3666 15874 3678
rect 21758 3666 21810 3678
rect 29934 3666 29986 3678
rect 9314 3614 9326 3666
rect 9378 3614 9390 3666
rect 11442 3614 11454 3666
rect 11506 3614 11518 3666
rect 13458 3614 13470 3666
rect 13522 3614 13534 3666
rect 16930 3614 16942 3666
rect 16994 3614 17006 3666
rect 19058 3614 19070 3666
rect 19122 3614 19134 3666
rect 20962 3614 20974 3666
rect 21026 3614 21038 3666
rect 23986 3614 23998 3666
rect 24050 3614 24062 3666
rect 27794 3614 27806 3666
rect 27858 3614 27870 3666
rect 7646 3602 7698 3614
rect 15822 3602 15874 3614
rect 21758 3602 21810 3614
rect 29934 3602 29986 3614
rect 33406 3666 33458 3678
rect 33406 3602 33458 3614
rect 34638 3666 34690 3678
rect 47406 3666 47458 3678
rect 38546 3614 38558 3666
rect 38610 3614 38622 3666
rect 41122 3614 41134 3666
rect 41186 3614 41198 3666
rect 41906 3614 41918 3666
rect 41970 3614 41982 3666
rect 34638 3602 34690 3614
rect 47406 3602 47458 3614
rect 56590 3666 56642 3678
rect 57362 3614 57374 3666
rect 57426 3614 57438 3666
rect 56590 3602 56642 3614
rect 28366 3554 28418 3566
rect 3154 3502 3166 3554
rect 3218 3502 3230 3554
rect 4722 3502 4734 3554
rect 4786 3502 4798 3554
rect 8082 3502 8094 3554
rect 8146 3502 8158 3554
rect 12114 3502 12126 3554
rect 12178 3502 12190 3554
rect 13682 3502 13694 3554
rect 13746 3502 13758 3554
rect 14690 3502 14702 3554
rect 14754 3502 14766 3554
rect 19842 3502 19854 3554
rect 19906 3502 19918 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 22418 3502 22430 3554
rect 22482 3502 22494 3554
rect 22978 3502 22990 3554
rect 23042 3502 23054 3554
rect 24994 3502 25006 3554
rect 25058 3502 25070 3554
rect 28366 3490 28418 3502
rect 30606 3554 30658 3566
rect 30606 3490 30658 3502
rect 35086 3554 35138 3566
rect 35086 3490 35138 3502
rect 37662 3554 37714 3566
rect 37662 3490 37714 3502
rect 38334 3554 38386 3566
rect 43486 3554 43538 3566
rect 41458 3502 41470 3554
rect 41522 3502 41534 3554
rect 42578 3502 42590 3554
rect 42642 3502 42654 3554
rect 38334 3490 38386 3502
rect 43486 3490 43538 3502
rect 43822 3554 43874 3566
rect 52782 3554 52834 3566
rect 45042 3502 45054 3554
rect 45106 3502 45118 3554
rect 45826 3502 45838 3554
rect 45890 3502 45902 3554
rect 47506 3502 47518 3554
rect 47570 3502 47582 3554
rect 47954 3502 47966 3554
rect 48018 3502 48030 3554
rect 43822 3490 43874 3502
rect 52782 3490 52834 3502
rect 56926 3554 56978 3566
rect 56926 3490 56978 3502
rect 2718 3442 2770 3454
rect 2718 3378 2770 3390
rect 2942 3442 2994 3454
rect 2942 3378 2994 3390
rect 4958 3442 5010 3454
rect 4958 3378 5010 3390
rect 5854 3442 5906 3454
rect 5854 3378 5906 3390
rect 7870 3442 7922 3454
rect 7870 3378 7922 3390
rect 8878 3442 8930 3454
rect 30942 3442 30994 3454
rect 15250 3390 15262 3442
rect 15314 3390 15326 3442
rect 25666 3390 25678 3442
rect 25730 3390 25742 3442
rect 8878 3378 8930 3390
rect 30942 3378 30994 3390
rect 31278 3442 31330 3454
rect 32846 3442 32898 3454
rect 32498 3390 32510 3442
rect 32562 3390 32574 3442
rect 31278 3378 31330 3390
rect 32846 3378 32898 3390
rect 34190 3442 34242 3454
rect 34190 3378 34242 3390
rect 37326 3442 37378 3454
rect 37326 3378 37378 3390
rect 41022 3442 41074 3454
rect 43710 3442 43762 3454
rect 51998 3442 52050 3454
rect 42130 3390 42142 3442
rect 42194 3390 42206 3442
rect 45938 3390 45950 3442
rect 46002 3390 46014 3442
rect 41022 3378 41074 3390
rect 43710 3378 43762 3390
rect 51998 3378 52050 3390
rect 52222 3442 52274 3454
rect 52222 3378 52274 3390
rect 30270 3330 30322 3342
rect 30270 3266 30322 3278
rect 33742 3330 33794 3342
rect 45042 3278 45054 3330
rect 45106 3278 45118 3330
rect 33742 3266 33794 3278
rect 1344 3162 58731 3196
rect 1344 3110 15520 3162
rect 15572 3110 15624 3162
rect 15676 3110 15728 3162
rect 15780 3110 29827 3162
rect 29879 3110 29931 3162
rect 29983 3110 30035 3162
rect 30087 3110 44134 3162
rect 44186 3110 44238 3162
rect 44290 3110 44342 3162
rect 44394 3110 58441 3162
rect 58493 3110 58545 3162
rect 58597 3110 58649 3162
rect 58701 3110 58731 3162
rect 1344 3076 58731 3110
<< via1 >>
rect 8367 36822 8419 36874
rect 8471 36822 8523 36874
rect 8575 36822 8627 36874
rect 22674 36822 22726 36874
rect 22778 36822 22830 36874
rect 22882 36822 22934 36874
rect 36981 36822 37033 36874
rect 37085 36822 37137 36874
rect 37189 36822 37241 36874
rect 51288 36822 51340 36874
rect 51392 36822 51444 36874
rect 51496 36822 51548 36874
rect 4622 36542 4674 36594
rect 8766 36542 8818 36594
rect 12574 36542 12626 36594
rect 14814 36542 14866 36594
rect 17390 36542 17442 36594
rect 19294 36542 19346 36594
rect 21534 36542 21586 36594
rect 23214 36542 23266 36594
rect 25678 36542 25730 36594
rect 27358 36542 27410 36594
rect 31278 36542 31330 36594
rect 35422 36542 35474 36594
rect 36542 36542 36594 36594
rect 41918 36542 41970 36594
rect 43038 36542 43090 36594
rect 43934 36542 43986 36594
rect 55022 36542 55074 36594
rect 56926 36542 56978 36594
rect 1822 36430 1874 36482
rect 5854 36430 5906 36482
rect 9774 36430 9826 36482
rect 14366 36430 14418 36482
rect 25006 36430 25058 36482
rect 28478 36430 28530 36482
rect 32622 36430 32674 36482
rect 37214 36430 37266 36482
rect 37998 36430 38050 36482
rect 38558 36430 38610 36482
rect 40798 36430 40850 36482
rect 41358 36430 41410 36482
rect 42254 36430 42306 36482
rect 46734 36430 46786 36482
rect 48862 36430 48914 36482
rect 49422 36430 49474 36482
rect 52782 36430 52834 36482
rect 53118 36430 53170 36482
rect 53790 36430 53842 36482
rect 55470 36430 55522 36482
rect 2494 36318 2546 36370
rect 6638 36318 6690 36370
rect 10446 36318 10498 36370
rect 15822 36318 15874 36370
rect 29150 36318 29202 36370
rect 33294 36318 33346 36370
rect 39230 36318 39282 36370
rect 39902 36318 39954 36370
rect 46062 36318 46114 36370
rect 47406 36318 47458 36370
rect 48302 36318 48354 36370
rect 49198 36318 49250 36370
rect 50542 36318 50594 36370
rect 51662 36318 51714 36370
rect 56478 36318 56530 36370
rect 13246 36206 13298 36258
rect 13694 36206 13746 36258
rect 16158 36206 16210 36258
rect 16942 36206 16994 36258
rect 18510 36206 18562 36258
rect 18846 36206 18898 36258
rect 20302 36206 20354 36258
rect 21086 36206 21138 36258
rect 22542 36206 22594 36258
rect 22766 36206 22818 36258
rect 24110 36206 24162 36258
rect 24670 36206 24722 36258
rect 26686 36206 26738 36258
rect 27806 36206 27858 36258
rect 42590 36206 42642 36258
rect 47742 36206 47794 36258
rect 50206 36206 50258 36258
rect 53566 36206 53618 36258
rect 54462 36206 54514 36258
rect 56030 36206 56082 36258
rect 15520 36038 15572 36090
rect 15624 36038 15676 36090
rect 15728 36038 15780 36090
rect 29827 36038 29879 36090
rect 29931 36038 29983 36090
rect 30035 36038 30087 36090
rect 44134 36038 44186 36090
rect 44238 36038 44290 36090
rect 44342 36038 44394 36090
rect 58441 36038 58493 36090
rect 58545 36038 58597 36090
rect 58649 36038 58701 36090
rect 9886 35870 9938 35922
rect 10670 35870 10722 35922
rect 21646 35870 21698 35922
rect 35534 35870 35586 35922
rect 51438 35870 51490 35922
rect 54686 35870 54738 35922
rect 54798 35870 54850 35922
rect 56030 35870 56082 35922
rect 2942 35758 2994 35810
rect 4958 35758 5010 35810
rect 16270 35758 16322 35810
rect 22766 35758 22818 35810
rect 37774 35758 37826 35810
rect 39790 35758 39842 35810
rect 40910 35758 40962 35810
rect 42702 35758 42754 35810
rect 44718 35758 44770 35810
rect 47630 35758 47682 35810
rect 48750 35758 48802 35810
rect 49086 35758 49138 35810
rect 50654 35758 50706 35810
rect 51774 35758 51826 35810
rect 55582 35758 55634 35810
rect 56702 35758 56754 35810
rect 1710 35646 1762 35698
rect 3838 35646 3890 35698
rect 4174 35646 4226 35698
rect 7646 35646 7698 35698
rect 11678 35646 11730 35698
rect 13134 35646 13186 35698
rect 16494 35646 16546 35698
rect 18286 35646 18338 35698
rect 21422 35646 21474 35698
rect 22542 35646 22594 35698
rect 22654 35646 22706 35698
rect 24222 35646 24274 35698
rect 26014 35646 26066 35698
rect 29598 35646 29650 35698
rect 33070 35646 33122 35698
rect 35870 35646 35922 35698
rect 36430 35646 36482 35698
rect 39902 35646 39954 35698
rect 41134 35646 41186 35698
rect 41694 35646 41746 35698
rect 43934 35646 43986 35698
rect 44830 35646 44882 35698
rect 46398 35646 46450 35698
rect 46846 35646 46898 35698
rect 47966 35646 48018 35698
rect 52782 35646 52834 35698
rect 53566 35646 53618 35698
rect 54574 35646 54626 35698
rect 55246 35646 55298 35698
rect 56478 35646 56530 35698
rect 56814 35646 56866 35698
rect 2158 35534 2210 35586
rect 7086 35534 7138 35586
rect 8094 35534 8146 35586
rect 8878 35534 8930 35586
rect 11118 35534 11170 35586
rect 12126 35534 12178 35586
rect 13806 35534 13858 35586
rect 15934 35534 15986 35586
rect 17838 35534 17890 35586
rect 18958 35534 19010 35586
rect 21086 35534 21138 35586
rect 24446 35534 24498 35586
rect 25678 35534 25730 35586
rect 26798 35534 26850 35586
rect 28926 35534 28978 35586
rect 30382 35534 30434 35586
rect 32510 35534 32562 35586
rect 33742 35534 33794 35586
rect 34526 35534 34578 35586
rect 37438 35534 37490 35586
rect 40126 35534 40178 35586
rect 42254 35534 42306 35586
rect 43822 35534 43874 35586
rect 45614 35534 45666 35586
rect 50878 35534 50930 35586
rect 52110 35534 52162 35586
rect 21758 35422 21810 35474
rect 22094 35422 22146 35474
rect 24558 35422 24610 35474
rect 40238 35422 40290 35474
rect 8367 35254 8419 35306
rect 8471 35254 8523 35306
rect 8575 35254 8627 35306
rect 22674 35254 22726 35306
rect 22778 35254 22830 35306
rect 22882 35254 22934 35306
rect 36981 35254 37033 35306
rect 37085 35254 37137 35306
rect 37189 35254 37241 35306
rect 51288 35254 51340 35306
rect 51392 35254 51444 35306
rect 51496 35254 51548 35306
rect 30494 35086 30546 35138
rect 35086 35086 35138 35138
rect 52894 35086 52946 35138
rect 53230 35086 53282 35138
rect 5070 34974 5122 35026
rect 5630 34974 5682 35026
rect 11790 34974 11842 35026
rect 14926 34974 14978 35026
rect 16046 34974 16098 35026
rect 18174 34974 18226 35026
rect 25566 34974 25618 35026
rect 30158 34974 30210 35026
rect 32174 34974 32226 35026
rect 36990 34974 37042 35026
rect 44046 34974 44098 35026
rect 45838 34974 45890 35026
rect 49086 34974 49138 35026
rect 51214 34974 51266 35026
rect 52670 34974 52722 35026
rect 56702 34974 56754 35026
rect 58158 34974 58210 35026
rect 1822 34862 1874 34914
rect 2270 34862 2322 34914
rect 2606 34862 2658 34914
rect 3166 34862 3218 34914
rect 3502 34862 3554 34914
rect 4062 34862 4114 34914
rect 8542 34862 8594 34914
rect 8990 34862 9042 34914
rect 12350 34862 12402 34914
rect 15262 34862 15314 34914
rect 20302 34862 20354 34914
rect 20526 34862 20578 34914
rect 21646 34862 21698 34914
rect 22430 34862 22482 34914
rect 22766 34862 22818 34914
rect 23998 34862 24050 34914
rect 25902 34862 25954 34914
rect 26462 34862 26514 34914
rect 28142 34862 28194 34914
rect 31278 34862 31330 34914
rect 32958 34862 33010 34914
rect 33742 34862 33794 34914
rect 33966 34862 34018 34914
rect 35758 34862 35810 34914
rect 40014 34862 40066 34914
rect 40462 34862 40514 34914
rect 42590 34862 42642 34914
rect 42926 34862 42978 34914
rect 46062 34862 46114 34914
rect 47630 34862 47682 34914
rect 47854 34862 47906 34914
rect 49422 34862 49474 34914
rect 50318 34862 50370 34914
rect 50542 34862 50594 34914
rect 54574 34862 54626 34914
rect 55470 34862 55522 34914
rect 57150 34862 57202 34914
rect 7758 34750 7810 34802
rect 9662 34750 9714 34802
rect 12126 34750 12178 34802
rect 13022 34750 13074 34802
rect 13806 34750 13858 34802
rect 14142 34750 14194 34802
rect 18734 34750 18786 34802
rect 19070 34750 19122 34802
rect 19630 34750 19682 34802
rect 21310 34750 21362 34802
rect 21422 34750 21474 34802
rect 21870 34750 21922 34802
rect 23438 34750 23490 34802
rect 25230 34750 25282 34802
rect 26350 34750 26402 34802
rect 27246 34750 27298 34802
rect 27582 34750 27634 34802
rect 28366 34750 28418 34802
rect 29374 34750 29426 34802
rect 29710 34750 29762 34802
rect 32734 34750 32786 34802
rect 33294 34750 33346 34802
rect 37102 34750 37154 34802
rect 37326 34750 37378 34802
rect 37886 34750 37938 34802
rect 39566 34750 39618 34802
rect 41022 34750 41074 34802
rect 44942 34750 44994 34802
rect 46846 34750 46898 34802
rect 49870 34750 49922 34802
rect 51550 34750 51602 34802
rect 54238 34750 54290 34802
rect 56142 34750 56194 34802
rect 57598 34750 57650 34802
rect 4622 34638 4674 34690
rect 26126 34638 26178 34690
rect 32846 34638 32898 34690
rect 33854 34638 33906 34690
rect 34190 34638 34242 34690
rect 34862 34638 34914 34690
rect 36430 34638 36482 34690
rect 37550 34638 37602 34690
rect 37774 34638 37826 34690
rect 38446 34638 38498 34690
rect 51662 34638 51714 34690
rect 51886 34638 51938 34690
rect 15520 34470 15572 34522
rect 15624 34470 15676 34522
rect 15728 34470 15780 34522
rect 29827 34470 29879 34522
rect 29931 34470 29983 34522
rect 30035 34470 30087 34522
rect 44134 34470 44186 34522
rect 44238 34470 44290 34522
rect 44342 34470 44394 34522
rect 58441 34470 58493 34522
rect 58545 34470 58597 34522
rect 58649 34470 58701 34522
rect 2718 34302 2770 34354
rect 4062 34302 4114 34354
rect 5406 34302 5458 34354
rect 6638 34302 6690 34354
rect 6974 34302 7026 34354
rect 7870 34302 7922 34354
rect 8766 34302 8818 34354
rect 9886 34302 9938 34354
rect 11902 34302 11954 34354
rect 17838 34302 17890 34354
rect 20414 34302 20466 34354
rect 21758 34302 21810 34354
rect 24222 34302 24274 34354
rect 28814 34302 28866 34354
rect 29374 34302 29426 34354
rect 30942 34302 30994 34354
rect 33182 34302 33234 34354
rect 36542 34302 36594 34354
rect 36766 34302 36818 34354
rect 42702 34302 42754 34354
rect 48190 34302 48242 34354
rect 50542 34302 50594 34354
rect 55134 34302 55186 34354
rect 3054 34190 3106 34242
rect 3502 34190 3554 34242
rect 4622 34190 4674 34242
rect 16606 34190 16658 34242
rect 21534 34190 21586 34242
rect 22094 34190 22146 34242
rect 28254 34190 28306 34242
rect 33518 34190 33570 34242
rect 35310 34190 35362 34242
rect 37998 34190 38050 34242
rect 40014 34190 40066 34242
rect 43710 34190 43762 34242
rect 45166 34190 45218 34242
rect 48862 34190 48914 34242
rect 49086 34190 49138 34242
rect 49422 34190 49474 34242
rect 50430 34190 50482 34242
rect 54686 34190 54738 34242
rect 56590 34190 56642 34242
rect 1710 34078 1762 34130
rect 3390 34078 3442 34130
rect 3726 34078 3778 34130
rect 4174 34078 4226 34130
rect 4398 34078 4450 34130
rect 4734 34078 4786 34130
rect 7310 34078 7362 34130
rect 8206 34078 8258 34130
rect 10222 34078 10274 34130
rect 12798 34078 12850 34130
rect 16270 34078 16322 34130
rect 18958 34078 19010 34130
rect 19518 34078 19570 34130
rect 19854 34078 19906 34130
rect 20302 34078 20354 34130
rect 20526 34078 20578 34130
rect 20974 34078 21026 34130
rect 21758 34078 21810 34130
rect 23102 34078 23154 34130
rect 23998 34078 24050 34130
rect 24558 34078 24610 34130
rect 25678 34078 25730 34130
rect 27582 34078 27634 34130
rect 31502 34078 31554 34130
rect 32174 34078 32226 34130
rect 34750 34078 34802 34130
rect 35982 34078 36034 34130
rect 36878 34078 36930 34130
rect 38222 34078 38274 34130
rect 39118 34078 39170 34130
rect 39566 34078 39618 34130
rect 40126 34078 40178 34130
rect 41022 34078 41074 34130
rect 41582 34078 41634 34130
rect 44158 34078 44210 34130
rect 46286 34078 46338 34130
rect 47070 34078 47122 34130
rect 47518 34078 47570 34130
rect 47742 34078 47794 34130
rect 48750 34078 48802 34130
rect 49534 34078 49586 34130
rect 50094 34078 50146 34130
rect 50654 34078 50706 34130
rect 51550 34078 51602 34130
rect 52894 34078 52946 34130
rect 53342 34078 53394 34130
rect 54238 34078 54290 34130
rect 54574 34078 54626 34130
rect 56702 34078 56754 34130
rect 57262 34078 57314 34130
rect 2158 33966 2210 34018
rect 5854 33966 5906 34018
rect 10670 33966 10722 34018
rect 11118 33966 11170 34018
rect 12350 33966 12402 34018
rect 13470 33966 13522 34018
rect 15598 33966 15650 34018
rect 18286 33966 18338 34018
rect 18734 33966 18786 34018
rect 22430 33966 22482 34018
rect 23326 33966 23378 34018
rect 24110 33966 24162 34018
rect 24558 33966 24610 34018
rect 24782 33966 24834 34018
rect 26014 33966 26066 34018
rect 26910 33966 26962 34018
rect 27918 33966 27970 34018
rect 29934 33966 29986 34018
rect 30494 33966 30546 34018
rect 32398 33966 32450 34018
rect 33966 33966 34018 34018
rect 34078 33966 34130 34018
rect 36206 33966 36258 34018
rect 40910 33966 40962 34018
rect 51102 33966 51154 34018
rect 58158 33966 58210 34018
rect 4062 33854 4114 33906
rect 25342 33854 25394 33906
rect 29710 33854 29762 33906
rect 40014 33854 40066 33906
rect 49422 33854 49474 33906
rect 8367 33686 8419 33738
rect 8471 33686 8523 33738
rect 8575 33686 8627 33738
rect 22674 33686 22726 33738
rect 22778 33686 22830 33738
rect 22882 33686 22934 33738
rect 36981 33686 37033 33738
rect 37085 33686 37137 33738
rect 37189 33686 37241 33738
rect 51288 33686 51340 33738
rect 51392 33686 51444 33738
rect 51496 33686 51548 33738
rect 35422 33518 35474 33570
rect 50766 33518 50818 33570
rect 51214 33518 51266 33570
rect 54462 33518 54514 33570
rect 4622 33406 4674 33458
rect 6190 33406 6242 33458
rect 8206 33406 8258 33458
rect 11566 33406 11618 33458
rect 12014 33406 12066 33458
rect 12574 33406 12626 33458
rect 12910 33406 12962 33458
rect 14366 33406 14418 33458
rect 14926 33406 14978 33458
rect 15710 33406 15762 33458
rect 16830 33406 16882 33458
rect 18958 33406 19010 33458
rect 20302 33406 20354 33458
rect 21982 33406 22034 33458
rect 26126 33406 26178 33458
rect 27918 33406 27970 33458
rect 28254 33406 28306 33458
rect 28590 33406 28642 33458
rect 29598 33406 29650 33458
rect 30158 33406 30210 33458
rect 33966 33406 34018 33458
rect 38558 33406 38610 33458
rect 39006 33406 39058 33458
rect 41246 33406 41298 33458
rect 43822 33406 43874 33458
rect 45390 33406 45442 33458
rect 46734 33406 46786 33458
rect 48862 33406 48914 33458
rect 53118 33406 53170 33458
rect 55806 33406 55858 33458
rect 57598 33406 57650 33458
rect 1822 33294 1874 33346
rect 11118 33294 11170 33346
rect 15262 33294 15314 33346
rect 16158 33294 16210 33346
rect 19854 33294 19906 33346
rect 20190 33294 20242 33346
rect 21198 33294 21250 33346
rect 21534 33294 21586 33346
rect 23214 33294 23266 33346
rect 24110 33294 24162 33346
rect 24894 33294 24946 33346
rect 25230 33294 25282 33346
rect 27246 33294 27298 33346
rect 27694 33294 27746 33346
rect 29486 33294 29538 33346
rect 30494 33294 30546 33346
rect 32622 33294 32674 33346
rect 33406 33294 33458 33346
rect 34302 33294 34354 33346
rect 34974 33294 35026 33346
rect 35534 33294 35586 33346
rect 37102 33294 37154 33346
rect 37662 33294 37714 33346
rect 39118 33294 39170 33346
rect 39454 33294 39506 33346
rect 40574 33294 40626 33346
rect 42702 33294 42754 33346
rect 43934 33294 43986 33346
rect 44382 33294 44434 33346
rect 45166 33294 45218 33346
rect 46286 33294 46338 33346
rect 48190 33294 48242 33346
rect 49198 33294 49250 33346
rect 49534 33294 49586 33346
rect 49758 33294 49810 33346
rect 50094 33294 50146 33346
rect 50766 33294 50818 33346
rect 53230 33294 53282 33346
rect 53566 33294 53618 33346
rect 53790 33294 53842 33346
rect 56030 33294 56082 33346
rect 57934 33294 57986 33346
rect 2494 33182 2546 33234
rect 10334 33182 10386 33234
rect 13582 33182 13634 33234
rect 13918 33182 13970 33234
rect 22766 33182 22818 33234
rect 32174 33182 32226 33234
rect 34526 33182 34578 33234
rect 35422 33182 35474 33234
rect 40350 33182 40402 33234
rect 41694 33182 41746 33234
rect 43374 33182 43426 33234
rect 43710 33182 43762 33234
rect 45838 33182 45890 33234
rect 46174 33182 46226 33234
rect 47294 33182 47346 33234
rect 49982 33182 50034 33234
rect 50430 33182 50482 33234
rect 51214 33182 51266 33234
rect 51326 33182 51378 33234
rect 54126 33182 54178 33234
rect 54574 33182 54626 33234
rect 5182 33070 5234 33122
rect 5854 33070 5906 33122
rect 6638 33070 6690 33122
rect 7086 33070 7138 33122
rect 7534 33070 7586 33122
rect 20862 33070 20914 33122
rect 21422 33070 21474 33122
rect 24334 33070 24386 33122
rect 25118 33070 25170 33122
rect 25678 33070 25730 33122
rect 26574 33070 26626 33122
rect 28478 33070 28530 33122
rect 30942 33070 30994 33122
rect 34638 33070 34690 33122
rect 36430 33070 36482 33122
rect 40798 33070 40850 33122
rect 40910 33070 40962 33122
rect 49310 33070 49362 33122
rect 51774 33070 51826 33122
rect 53006 33070 53058 33122
rect 54014 33070 54066 33122
rect 15520 32902 15572 32954
rect 15624 32902 15676 32954
rect 15728 32902 15780 32954
rect 29827 32902 29879 32954
rect 29931 32902 29983 32954
rect 30035 32902 30087 32954
rect 44134 32902 44186 32954
rect 44238 32902 44290 32954
rect 44342 32902 44394 32954
rect 58441 32902 58493 32954
rect 58545 32902 58597 32954
rect 58649 32902 58701 32954
rect 2494 32734 2546 32786
rect 7198 32734 7250 32786
rect 8878 32734 8930 32786
rect 9662 32734 9714 32786
rect 11790 32734 11842 32786
rect 15262 32734 15314 32786
rect 17726 32734 17778 32786
rect 20190 32734 20242 32786
rect 23214 32734 23266 32786
rect 23886 32734 23938 32786
rect 24446 32734 24498 32786
rect 27694 32734 27746 32786
rect 29822 32734 29874 32786
rect 33294 32734 33346 32786
rect 38782 32734 38834 32786
rect 42814 32734 42866 32786
rect 43934 32734 43986 32786
rect 53230 32734 53282 32786
rect 56142 32734 56194 32786
rect 58158 32734 58210 32786
rect 1822 32622 1874 32674
rect 1934 32622 1986 32674
rect 2382 32622 2434 32674
rect 2718 32622 2770 32674
rect 6638 32622 6690 32674
rect 6750 32622 6802 32674
rect 7982 32622 8034 32674
rect 8318 32622 8370 32674
rect 10782 32622 10834 32674
rect 16158 32622 16210 32674
rect 18958 32622 19010 32674
rect 21758 32622 21810 32674
rect 23102 32622 23154 32674
rect 26238 32622 26290 32674
rect 30382 32622 30434 32674
rect 30606 32622 30658 32674
rect 34414 32622 34466 32674
rect 36318 32622 36370 32674
rect 36542 32622 36594 32674
rect 36990 32622 37042 32674
rect 38670 32622 38722 32674
rect 39342 32622 39394 32674
rect 41918 32622 41970 32674
rect 43822 32622 43874 32674
rect 47854 32622 47906 32674
rect 48750 32622 48802 32674
rect 50542 32622 50594 32674
rect 51998 32622 52050 32674
rect 54910 32622 54962 32674
rect 55806 32622 55858 32674
rect 55918 32622 55970 32674
rect 56590 32622 56642 32674
rect 2158 32510 2210 32562
rect 2942 32510 2994 32562
rect 3278 32510 3330 32562
rect 6414 32510 6466 32562
rect 8542 32510 8594 32562
rect 9438 32510 9490 32562
rect 9774 32510 9826 32562
rect 10110 32510 10162 32562
rect 10670 32510 10722 32562
rect 13246 32510 13298 32562
rect 14590 32510 14642 32562
rect 15150 32510 15202 32562
rect 15374 32510 15426 32562
rect 15822 32510 15874 32562
rect 18062 32510 18114 32562
rect 26126 32510 26178 32562
rect 28590 32510 28642 32562
rect 28926 32510 28978 32562
rect 29374 32510 29426 32562
rect 30270 32510 30322 32562
rect 30830 32510 30882 32562
rect 31838 32510 31890 32562
rect 32286 32510 32338 32562
rect 33070 32510 33122 32562
rect 33182 32510 33234 32562
rect 34302 32510 34354 32562
rect 36654 32510 36706 32562
rect 37438 32510 37490 32562
rect 38446 32510 38498 32562
rect 39118 32510 39170 32562
rect 39454 32510 39506 32562
rect 40350 32510 40402 32562
rect 41470 32510 41522 32562
rect 42030 32510 42082 32562
rect 43374 32510 43426 32562
rect 44046 32510 44098 32562
rect 44830 32510 44882 32562
rect 46286 32510 46338 32562
rect 46622 32510 46674 32562
rect 48078 32510 48130 32562
rect 49422 32510 49474 32562
rect 52894 32510 52946 32562
rect 54238 32510 54290 32562
rect 57486 32510 57538 32562
rect 4062 32398 4114 32450
rect 6190 32398 6242 32450
rect 11454 32398 11506 32450
rect 14702 32398 14754 32450
rect 16046 32398 16098 32450
rect 16830 32398 16882 32450
rect 19518 32398 19570 32450
rect 20750 32398 20802 32450
rect 21422 32398 21474 32450
rect 28030 32398 28082 32450
rect 28254 32398 28306 32450
rect 31390 32398 31442 32450
rect 37774 32398 37826 32450
rect 40238 32398 40290 32450
rect 40910 32398 40962 32450
rect 43262 32398 43314 32450
rect 44494 32398 44546 32450
rect 45390 32398 45442 32450
rect 46734 32398 46786 32450
rect 47182 32398 47234 32450
rect 50878 32398 50930 32450
rect 51438 32398 51490 32450
rect 54014 32398 54066 32450
rect 55470 32398 55522 32450
rect 57150 32398 57202 32450
rect 13022 32286 13074 32338
rect 16382 32286 16434 32338
rect 26238 32286 26290 32338
rect 29150 32286 29202 32338
rect 34414 32286 34466 32338
rect 38782 32286 38834 32338
rect 41246 32286 41298 32338
rect 41918 32286 41970 32338
rect 8367 32118 8419 32170
rect 8471 32118 8523 32170
rect 8575 32118 8627 32170
rect 22674 32118 22726 32170
rect 22778 32118 22830 32170
rect 22882 32118 22934 32170
rect 36981 32118 37033 32170
rect 37085 32118 37137 32170
rect 37189 32118 37241 32170
rect 51288 32118 51340 32170
rect 51392 32118 51444 32170
rect 51496 32118 51548 32170
rect 32398 31950 32450 32002
rect 33406 31950 33458 32002
rect 37438 31950 37490 32002
rect 46958 31950 47010 32002
rect 53342 31950 53394 32002
rect 55806 31950 55858 32002
rect 7198 31838 7250 31890
rect 7534 31838 7586 31890
rect 18510 31838 18562 31890
rect 20190 31838 20242 31890
rect 21534 31838 21586 31890
rect 27134 31838 27186 31890
rect 31838 31838 31890 31890
rect 33854 31838 33906 31890
rect 36430 31838 36482 31890
rect 37774 31838 37826 31890
rect 43710 31838 43762 31890
rect 45726 31838 45778 31890
rect 51326 31838 51378 31890
rect 53678 31838 53730 31890
rect 1822 31726 1874 31778
rect 2270 31726 2322 31778
rect 3838 31726 3890 31778
rect 3950 31726 4002 31778
rect 5966 31726 6018 31778
rect 8430 31726 8482 31778
rect 9550 31726 9602 31778
rect 10670 31726 10722 31778
rect 14254 31726 14306 31778
rect 14814 31726 14866 31778
rect 15150 31726 15202 31778
rect 15822 31726 15874 31778
rect 16158 31726 16210 31778
rect 16494 31726 16546 31778
rect 17054 31726 17106 31778
rect 18286 31726 18338 31778
rect 19406 31726 19458 31778
rect 19742 31726 19794 31778
rect 20302 31726 20354 31778
rect 25902 31726 25954 31778
rect 26238 31726 26290 31778
rect 26574 31726 26626 31778
rect 27358 31726 27410 31778
rect 27694 31726 27746 31778
rect 30158 31726 30210 31778
rect 33294 31726 33346 31778
rect 34526 31726 34578 31778
rect 34750 31726 34802 31778
rect 35534 31726 35586 31778
rect 35982 31726 36034 31778
rect 37886 31726 37938 31778
rect 39678 31726 39730 31778
rect 40126 31726 40178 31778
rect 40574 31726 40626 31778
rect 41022 31726 41074 31778
rect 41358 31726 41410 31778
rect 42478 31726 42530 31778
rect 42702 31726 42754 31778
rect 44718 31726 44770 31778
rect 45054 31726 45106 31778
rect 45614 31726 45666 31778
rect 46174 31726 46226 31778
rect 48190 31726 48242 31778
rect 49086 31726 49138 31778
rect 51998 31726 52050 31778
rect 53566 31726 53618 31778
rect 54686 31726 54738 31778
rect 54910 31726 54962 31778
rect 55134 31726 55186 31778
rect 56030 31726 56082 31778
rect 56926 31726 56978 31778
rect 57262 31726 57314 31778
rect 3278 31614 3330 31666
rect 4286 31614 4338 31666
rect 4622 31614 4674 31666
rect 4958 31614 5010 31666
rect 5630 31614 5682 31666
rect 5742 31614 5794 31666
rect 6638 31614 6690 31666
rect 6974 31614 7026 31666
rect 8318 31614 8370 31666
rect 9214 31614 9266 31666
rect 9326 31614 9378 31666
rect 15598 31614 15650 31666
rect 16382 31614 16434 31666
rect 17390 31614 17442 31666
rect 18734 31614 18786 31666
rect 21646 31614 21698 31666
rect 23326 31614 23378 31666
rect 25566 31614 25618 31666
rect 29150 31614 29202 31666
rect 31502 31614 31554 31666
rect 32734 31614 32786 31666
rect 33406 31614 33458 31666
rect 38894 31614 38946 31666
rect 41134 31614 41186 31666
rect 42926 31614 42978 31666
rect 44942 31614 44994 31666
rect 47070 31614 47122 31666
rect 48078 31614 48130 31666
rect 50094 31614 50146 31666
rect 2718 31502 2770 31554
rect 2942 31502 2994 31554
rect 3166 31502 3218 31554
rect 4062 31502 4114 31554
rect 8094 31502 8146 31554
rect 8878 31502 8930 31554
rect 9886 31502 9938 31554
rect 10334 31502 10386 31554
rect 10782 31502 10834 31554
rect 11006 31502 11058 31554
rect 17278 31502 17330 31554
rect 17950 31502 18002 31554
rect 23214 31502 23266 31554
rect 24110 31502 24162 31554
rect 24334 31502 24386 31554
rect 24446 31502 24498 31554
rect 24558 31502 24610 31554
rect 25678 31502 25730 31554
rect 27582 31502 27634 31554
rect 28590 31502 28642 31554
rect 32510 31502 32562 31554
rect 39230 31502 39282 31554
rect 43598 31502 43650 31554
rect 43822 31502 43874 31554
rect 44046 31502 44098 31554
rect 50878 31502 50930 31554
rect 51774 31502 51826 31554
rect 15520 31334 15572 31386
rect 15624 31334 15676 31386
rect 15728 31334 15780 31386
rect 29827 31334 29879 31386
rect 29931 31334 29983 31386
rect 30035 31334 30087 31386
rect 44134 31334 44186 31386
rect 44238 31334 44290 31386
rect 44342 31334 44394 31386
rect 58441 31334 58493 31386
rect 58545 31334 58597 31386
rect 58649 31334 58701 31386
rect 15822 31166 15874 31218
rect 16382 31166 16434 31218
rect 18958 31166 19010 31218
rect 19294 31166 19346 31218
rect 19406 31166 19458 31218
rect 20302 31166 20354 31218
rect 21422 31166 21474 31218
rect 23886 31166 23938 31218
rect 33182 31166 33234 31218
rect 40014 31166 40066 31218
rect 40910 31166 40962 31218
rect 45390 31166 45442 31218
rect 15710 31054 15762 31106
rect 19742 31054 19794 31106
rect 22318 31054 22370 31106
rect 23998 31054 24050 31106
rect 26014 31054 26066 31106
rect 28254 31054 28306 31106
rect 33294 31054 33346 31106
rect 34750 31054 34802 31106
rect 35198 31054 35250 31106
rect 36318 31054 36370 31106
rect 38670 31054 38722 31106
rect 45502 31054 45554 31106
rect 45950 31054 46002 31106
rect 55246 31054 55298 31106
rect 56590 31054 56642 31106
rect 58046 31054 58098 31106
rect 1710 30942 1762 30994
rect 2830 30942 2882 30994
rect 6190 30942 6242 30994
rect 10110 30942 10162 30994
rect 14814 30942 14866 30994
rect 15038 30942 15090 30994
rect 15486 30942 15538 30994
rect 19518 30942 19570 30994
rect 20414 30942 20466 30994
rect 22878 30942 22930 30994
rect 26686 30942 26738 30994
rect 26910 30942 26962 30994
rect 29150 30942 29202 30994
rect 29822 30942 29874 30994
rect 31614 30942 31666 30994
rect 34078 30942 34130 30994
rect 37550 30942 37602 30994
rect 40350 30942 40402 30994
rect 42590 30942 42642 30994
rect 43934 30942 43986 30994
rect 45166 30942 45218 30994
rect 46398 30942 46450 30994
rect 46734 30942 46786 30994
rect 47966 30942 48018 30994
rect 49086 30942 49138 30994
rect 49422 30942 49474 30994
rect 51662 30942 51714 30994
rect 53006 30942 53058 30994
rect 53790 30942 53842 30994
rect 55470 30942 55522 30994
rect 57038 30942 57090 30994
rect 2270 30830 2322 30882
rect 3614 30830 3666 30882
rect 5742 30830 5794 30882
rect 6862 30830 6914 30882
rect 8990 30830 9042 30882
rect 9662 30830 9714 30882
rect 10782 30830 10834 30882
rect 12910 30830 12962 30882
rect 14926 30830 14978 30882
rect 17614 30830 17666 30882
rect 18398 30830 18450 30882
rect 20862 30830 20914 30882
rect 28366 30830 28418 30882
rect 28926 30830 28978 30882
rect 29374 30830 29426 30882
rect 30606 30830 30658 30882
rect 31838 30830 31890 30882
rect 32286 30830 32338 30882
rect 33070 30830 33122 30882
rect 34414 30830 34466 30882
rect 36094 30830 36146 30882
rect 41470 30830 41522 30882
rect 42478 30830 42530 30882
rect 48862 30830 48914 30882
rect 49310 30830 49362 30882
rect 51774 30830 51826 30882
rect 54238 30830 54290 30882
rect 56142 30830 56194 30882
rect 57374 30830 57426 30882
rect 15822 30718 15874 30770
rect 18622 30718 18674 30770
rect 28478 30718 28530 30770
rect 41246 30718 41298 30770
rect 44494 30718 44546 30770
rect 50766 30718 50818 30770
rect 8367 30550 8419 30602
rect 8471 30550 8523 30602
rect 8575 30550 8627 30602
rect 22674 30550 22726 30602
rect 22778 30550 22830 30602
rect 22882 30550 22934 30602
rect 36981 30550 37033 30602
rect 37085 30550 37137 30602
rect 37189 30550 37241 30602
rect 51288 30550 51340 30602
rect 51392 30550 51444 30602
rect 51496 30550 51548 30602
rect 6974 30382 7026 30434
rect 7310 30382 7362 30434
rect 19630 30382 19682 30434
rect 19966 30382 20018 30434
rect 23998 30382 24050 30434
rect 31726 30382 31778 30434
rect 55358 30382 55410 30434
rect 10670 30270 10722 30322
rect 16606 30270 16658 30322
rect 18510 30270 18562 30322
rect 21534 30270 21586 30322
rect 24558 30270 24610 30322
rect 27694 30270 27746 30322
rect 34078 30270 34130 30322
rect 38558 30270 38610 30322
rect 40686 30270 40738 30322
rect 43038 30270 43090 30322
rect 45838 30270 45890 30322
rect 48974 30270 49026 30322
rect 54462 30270 54514 30322
rect 57150 30270 57202 30322
rect 2942 30158 2994 30210
rect 3614 30158 3666 30210
rect 4398 30158 4450 30210
rect 5630 30158 5682 30210
rect 5966 30158 6018 30210
rect 7534 30158 7586 30210
rect 7870 30158 7922 30210
rect 9998 30158 10050 30210
rect 10558 30158 10610 30210
rect 11342 30158 11394 30210
rect 15038 30158 15090 30210
rect 18846 30158 18898 30210
rect 26014 30158 26066 30210
rect 27918 30158 27970 30210
rect 28590 30158 28642 30210
rect 29150 30158 29202 30210
rect 29486 30158 29538 30210
rect 30046 30158 30098 30210
rect 31390 30158 31442 30210
rect 32398 30158 32450 30210
rect 33182 30158 33234 30210
rect 33630 30158 33682 30210
rect 37662 30158 37714 30210
rect 40014 30158 40066 30210
rect 43486 30158 43538 30210
rect 44270 30158 44322 30210
rect 47182 30158 47234 30210
rect 50430 30158 50482 30210
rect 52670 30158 52722 30210
rect 53230 30158 53282 30210
rect 55694 30158 55746 30210
rect 56702 30158 56754 30210
rect 57934 30158 57986 30210
rect 1710 30046 1762 30098
rect 2046 30046 2098 30098
rect 4734 30046 4786 30098
rect 4958 30046 5010 30098
rect 6414 30046 6466 30098
rect 6638 30046 6690 30098
rect 6750 30046 6802 30098
rect 8094 30046 8146 30098
rect 10222 30046 10274 30098
rect 10782 30046 10834 30098
rect 11118 30046 11170 30098
rect 14926 30046 14978 30098
rect 16382 30046 16434 30098
rect 19294 30046 19346 30098
rect 20190 30046 20242 30098
rect 21646 30046 21698 30098
rect 23326 30046 23378 30098
rect 23886 30046 23938 30098
rect 24782 30046 24834 30098
rect 29374 30046 29426 30098
rect 31614 30046 31666 30098
rect 36990 30046 37042 30098
rect 37214 30046 37266 30098
rect 38782 30046 38834 30098
rect 42814 30046 42866 30098
rect 46286 30046 46338 30098
rect 48526 30046 48578 30098
rect 49422 30046 49474 30098
rect 53342 30046 53394 30098
rect 54126 30046 54178 30098
rect 57598 30046 57650 30098
rect 2382 29934 2434 29986
rect 3726 29934 3778 29986
rect 3950 29934 4002 29986
rect 4510 29934 4562 29986
rect 5742 29934 5794 29986
rect 7198 29934 7250 29986
rect 7646 29934 7698 29986
rect 8542 29934 8594 29986
rect 13694 29934 13746 29986
rect 17054 29934 17106 29986
rect 23214 29934 23266 29986
rect 23998 29934 24050 29986
rect 26574 29934 26626 29986
rect 37326 29934 37378 29986
rect 45166 29934 45218 29986
rect 51774 29934 51826 29986
rect 52782 29934 52834 29986
rect 54350 29934 54402 29986
rect 57710 29934 57762 29986
rect 15520 29766 15572 29818
rect 15624 29766 15676 29818
rect 15728 29766 15780 29818
rect 29827 29766 29879 29818
rect 29931 29766 29983 29818
rect 30035 29766 30087 29818
rect 44134 29766 44186 29818
rect 44238 29766 44290 29818
rect 44342 29766 44394 29818
rect 58441 29766 58493 29818
rect 58545 29766 58597 29818
rect 58649 29766 58701 29818
rect 13806 29598 13858 29650
rect 19966 29598 20018 29650
rect 20526 29598 20578 29650
rect 20750 29598 20802 29650
rect 21534 29598 21586 29650
rect 25678 29598 25730 29650
rect 29262 29598 29314 29650
rect 31950 29598 32002 29650
rect 32062 29598 32114 29650
rect 32398 29598 32450 29650
rect 35534 29598 35586 29650
rect 42926 29598 42978 29650
rect 47966 29598 48018 29650
rect 48078 29598 48130 29650
rect 48974 29598 49026 29650
rect 15374 29486 15426 29538
rect 18174 29486 18226 29538
rect 20190 29486 20242 29538
rect 20862 29486 20914 29538
rect 21310 29486 21362 29538
rect 23662 29486 23714 29538
rect 28030 29486 28082 29538
rect 29934 29486 29986 29538
rect 34526 29486 34578 29538
rect 34638 29486 34690 29538
rect 35422 29486 35474 29538
rect 36990 29486 37042 29538
rect 42814 29486 42866 29538
rect 45726 29486 45778 29538
rect 50206 29486 50258 29538
rect 51550 29486 51602 29538
rect 53790 29486 53842 29538
rect 54350 29486 54402 29538
rect 55806 29486 55858 29538
rect 55918 29486 55970 29538
rect 56926 29486 56978 29538
rect 1822 29374 1874 29426
rect 5294 29374 5346 29426
rect 10222 29374 10274 29426
rect 13582 29374 13634 29426
rect 14702 29374 14754 29426
rect 19294 29374 19346 29426
rect 19742 29374 19794 29426
rect 20302 29374 20354 29426
rect 21198 29374 21250 29426
rect 23774 29374 23826 29426
rect 24334 29374 24386 29426
rect 29038 29374 29090 29426
rect 30606 29374 30658 29426
rect 31614 29374 31666 29426
rect 32174 29374 32226 29426
rect 33630 29374 33682 29426
rect 36542 29374 36594 29426
rect 37774 29374 37826 29426
rect 38222 29374 38274 29426
rect 39902 29374 39954 29426
rect 44158 29374 44210 29426
rect 45278 29374 45330 29426
rect 50094 29374 50146 29426
rect 53006 29374 53058 29426
rect 54574 29374 54626 29426
rect 54798 29374 54850 29426
rect 56142 29374 56194 29426
rect 56590 29374 56642 29426
rect 57710 29374 57762 29426
rect 2606 29262 2658 29314
rect 4734 29262 4786 29314
rect 6078 29262 6130 29314
rect 8206 29262 8258 29314
rect 10894 29262 10946 29314
rect 13022 29262 13074 29314
rect 14926 29262 14978 29314
rect 17726 29262 17778 29314
rect 21870 29262 21922 29314
rect 25790 29262 25842 29314
rect 27470 29262 27522 29314
rect 30270 29262 30322 29314
rect 31390 29262 31442 29314
rect 33294 29262 33346 29314
rect 34078 29262 34130 29314
rect 36094 29262 36146 29314
rect 37326 29262 37378 29314
rect 39566 29262 39618 29314
rect 40350 29262 40402 29314
rect 43934 29262 43986 29314
rect 44942 29262 44994 29314
rect 46174 29262 46226 29314
rect 51214 29262 51266 29314
rect 57150 29262 57202 29314
rect 58158 29262 58210 29314
rect 31278 29150 31330 29202
rect 34526 29150 34578 29202
rect 35646 29150 35698 29202
rect 43598 29150 43650 29202
rect 48190 29150 48242 29202
rect 8367 28982 8419 29034
rect 8471 28982 8523 29034
rect 8575 28982 8627 29034
rect 22674 28982 22726 29034
rect 22778 28982 22830 29034
rect 22882 28982 22934 29034
rect 36981 28982 37033 29034
rect 37085 28982 37137 29034
rect 37189 28982 37241 29034
rect 51288 28982 51340 29034
rect 51392 28982 51444 29034
rect 51496 28982 51548 29034
rect 8318 28814 8370 28866
rect 8654 28814 8706 28866
rect 9886 28814 9938 28866
rect 12798 28814 12850 28866
rect 14926 28814 14978 28866
rect 21982 28814 22034 28866
rect 25118 28814 25170 28866
rect 27918 28814 27970 28866
rect 33854 28814 33906 28866
rect 37438 28814 37490 28866
rect 38222 28814 38274 28866
rect 43710 28814 43762 28866
rect 44046 28814 44098 28866
rect 44942 28814 44994 28866
rect 49198 28814 49250 28866
rect 55694 28814 55746 28866
rect 3054 28702 3106 28754
rect 5070 28702 5122 28754
rect 5742 28702 5794 28754
rect 10446 28702 10498 28754
rect 15150 28702 15202 28754
rect 19742 28702 19794 28754
rect 20638 28702 20690 28754
rect 23438 28702 23490 28754
rect 24446 28702 24498 28754
rect 24894 28702 24946 28754
rect 25902 28702 25954 28754
rect 27134 28702 27186 28754
rect 28478 28702 28530 28754
rect 30046 28702 30098 28754
rect 30494 28702 30546 28754
rect 31166 28702 31218 28754
rect 33294 28702 33346 28754
rect 37662 28702 37714 28754
rect 42702 28702 42754 28754
rect 43374 28702 43426 28754
rect 46398 28702 46450 28754
rect 49758 28702 49810 28754
rect 50318 28702 50370 28754
rect 52782 28702 52834 28754
rect 57934 28702 57986 28754
rect 1934 28590 1986 28642
rect 2158 28590 2210 28642
rect 2830 28590 2882 28642
rect 3278 28590 3330 28642
rect 3726 28590 3778 28642
rect 4734 28590 4786 28642
rect 5518 28590 5570 28642
rect 5966 28590 6018 28642
rect 6078 28590 6130 28642
rect 6750 28590 6802 28642
rect 9438 28590 9490 28642
rect 10222 28590 10274 28642
rect 10670 28590 10722 28642
rect 11118 28590 11170 28642
rect 11454 28590 11506 28642
rect 11678 28590 11730 28642
rect 12014 28590 12066 28642
rect 14254 28590 14306 28642
rect 15374 28590 15426 28642
rect 18846 28590 18898 28642
rect 19070 28590 19122 28642
rect 21198 28590 21250 28642
rect 22990 28590 23042 28642
rect 23326 28590 23378 28642
rect 23998 28590 24050 28642
rect 30606 28590 30658 28642
rect 32846 28590 32898 28642
rect 33182 28590 33234 28642
rect 33406 28590 33458 28642
rect 33742 28590 33794 28642
rect 35982 28590 36034 28642
rect 36878 28590 36930 28642
rect 38782 28590 38834 28642
rect 39566 28590 39618 28642
rect 40798 28590 40850 28642
rect 41582 28590 41634 28642
rect 44270 28590 44322 28642
rect 45278 28590 45330 28642
rect 48190 28590 48242 28642
rect 49982 28590 50034 28642
rect 51438 28590 51490 28642
rect 51886 28590 51938 28642
rect 53230 28590 53282 28642
rect 54574 28590 54626 28642
rect 55022 28590 55074 28642
rect 56366 28590 56418 28642
rect 2494 28478 2546 28530
rect 3502 28478 3554 28530
rect 3950 28478 4002 28530
rect 4062 28478 4114 28530
rect 4398 28478 4450 28530
rect 6974 28478 7026 28530
rect 7086 28478 7138 28530
rect 7646 28478 7698 28530
rect 7982 28478 8034 28530
rect 9998 28478 10050 28530
rect 10894 28478 10946 28530
rect 12238 28478 12290 28530
rect 12350 28478 12402 28530
rect 12686 28478 12738 28530
rect 12798 28478 12850 28530
rect 14478 28478 14530 28530
rect 20190 28478 20242 28530
rect 21534 28478 21586 28530
rect 21982 28478 22034 28530
rect 22094 28478 22146 28530
rect 24334 28478 24386 28530
rect 27134 28478 27186 28530
rect 31502 28478 31554 28530
rect 36318 28478 36370 28530
rect 37102 28478 37154 28530
rect 37214 28478 37266 28530
rect 39678 28478 39730 28530
rect 40686 28478 40738 28530
rect 45054 28478 45106 28530
rect 45502 28478 45554 28530
rect 45614 28478 45666 28530
rect 46622 28478 46674 28530
rect 52110 28478 52162 28530
rect 57374 28478 57426 28530
rect 4510 28366 4562 28418
rect 9886 28366 9938 28418
rect 11454 28366 11506 28418
rect 13918 28366 13970 28418
rect 21422 28366 21474 28418
rect 24558 28366 24610 28418
rect 25454 28366 25506 28418
rect 25790 28366 25842 28418
rect 31278 28366 31330 28418
rect 34526 28366 34578 28418
rect 35758 28366 35810 28418
rect 36206 28366 36258 28418
rect 38222 28366 38274 28418
rect 38670 28366 38722 28418
rect 44942 28366 44994 28418
rect 15520 28198 15572 28250
rect 15624 28198 15676 28250
rect 15728 28198 15780 28250
rect 29827 28198 29879 28250
rect 29931 28198 29983 28250
rect 30035 28198 30087 28250
rect 44134 28198 44186 28250
rect 44238 28198 44290 28250
rect 44342 28198 44394 28250
rect 58441 28198 58493 28250
rect 58545 28198 58597 28250
rect 58649 28198 58701 28250
rect 1710 28030 1762 28082
rect 2718 28030 2770 28082
rect 3054 28030 3106 28082
rect 4734 28030 4786 28082
rect 7422 28030 7474 28082
rect 9550 28030 9602 28082
rect 10334 28030 10386 28082
rect 10782 28030 10834 28082
rect 11006 28030 11058 28082
rect 16494 28030 16546 28082
rect 18062 28030 18114 28082
rect 18510 28030 18562 28082
rect 20526 28030 20578 28082
rect 22318 28030 22370 28082
rect 22542 28030 22594 28082
rect 35422 28030 35474 28082
rect 39902 28030 39954 28082
rect 41022 28030 41074 28082
rect 49310 28030 49362 28082
rect 49534 28030 49586 28082
rect 49758 28030 49810 28082
rect 52222 28030 52274 28082
rect 54238 28030 54290 28082
rect 57262 28030 57314 28082
rect 2046 27918 2098 27970
rect 4286 27918 4338 27970
rect 7982 27918 8034 27970
rect 12126 27918 12178 27970
rect 15262 27918 15314 27970
rect 16606 27918 16658 27970
rect 18622 27918 18674 27970
rect 25454 27918 25506 27970
rect 30270 27918 30322 27970
rect 32174 27918 32226 27970
rect 37326 27918 37378 27970
rect 39566 27918 39618 27970
rect 40910 27918 40962 27970
rect 42478 27918 42530 27970
rect 47294 27918 47346 27970
rect 48190 27918 48242 27970
rect 51886 27918 51938 27970
rect 52446 27918 52498 27970
rect 2382 27806 2434 27858
rect 3278 27806 3330 27858
rect 4062 27806 4114 27858
rect 7086 27806 7138 27858
rect 8430 27806 8482 27858
rect 9886 27806 9938 27858
rect 10670 27806 10722 27858
rect 11454 27806 11506 27858
rect 18286 27806 18338 27858
rect 19406 27806 19458 27858
rect 20302 27806 20354 27858
rect 20862 27806 20914 27858
rect 22206 27806 22258 27858
rect 24222 27806 24274 27858
rect 25902 27806 25954 27858
rect 27694 27806 27746 27858
rect 28030 27806 28082 27858
rect 28814 27806 28866 27858
rect 30942 27806 30994 27858
rect 34190 27806 34242 27858
rect 34638 27806 34690 27858
rect 34974 27806 35026 27858
rect 35310 27806 35362 27858
rect 35646 27806 35698 27858
rect 37438 27806 37490 27858
rect 38222 27806 38274 27858
rect 41246 27806 41298 27858
rect 42702 27806 42754 27858
rect 43374 27806 43426 27858
rect 43710 27806 43762 27858
rect 44270 27806 44322 27858
rect 45502 27806 45554 27858
rect 45950 27806 46002 27858
rect 46846 27806 46898 27858
rect 47630 27806 47682 27858
rect 47854 27806 47906 27858
rect 48078 27806 48130 27858
rect 49198 27862 49250 27914
rect 52558 27918 52610 27970
rect 54126 27918 54178 27970
rect 55022 27918 55074 27970
rect 57822 27918 57874 27970
rect 50206 27806 50258 27858
rect 50318 27806 50370 27858
rect 50542 27806 50594 27858
rect 50878 27806 50930 27858
rect 51438 27806 51490 27858
rect 53006 27806 53058 27858
rect 54350 27806 54402 27858
rect 54686 27806 54738 27858
rect 55134 27806 55186 27858
rect 55470 27806 55522 27858
rect 57038 27806 57090 27858
rect 5182 27694 5234 27746
rect 8990 27694 9042 27746
rect 14254 27694 14306 27746
rect 14814 27694 14866 27746
rect 18958 27694 19010 27746
rect 19854 27694 19906 27746
rect 20414 27694 20466 27746
rect 21758 27694 21810 27746
rect 22878 27694 22930 27746
rect 24334 27694 24386 27746
rect 24670 27694 24722 27746
rect 25230 27694 25282 27746
rect 25566 27694 25618 27746
rect 28142 27694 28194 27746
rect 28478 27694 28530 27746
rect 28590 27694 28642 27746
rect 32286 27694 32338 27746
rect 33742 27694 33794 27746
rect 40014 27694 40066 27746
rect 42366 27694 42418 27746
rect 45054 27694 45106 27746
rect 46958 27694 47010 27746
rect 48862 27694 48914 27746
rect 51550 27694 51602 27746
rect 52894 27694 52946 27746
rect 53902 27694 53954 27746
rect 57150 27694 57202 27746
rect 57710 27694 57762 27746
rect 4734 27582 4786 27634
rect 5182 27582 5234 27634
rect 25902 27582 25954 27634
rect 26238 27582 26290 27634
rect 58046 27582 58098 27634
rect 8367 27414 8419 27466
rect 8471 27414 8523 27466
rect 8575 27414 8627 27466
rect 22674 27414 22726 27466
rect 22778 27414 22830 27466
rect 22882 27414 22934 27466
rect 36981 27414 37033 27466
rect 37085 27414 37137 27466
rect 37189 27414 37241 27466
rect 51288 27414 51340 27466
rect 51392 27414 51444 27466
rect 51496 27414 51548 27466
rect 16494 27246 16546 27298
rect 20078 27246 20130 27298
rect 34414 27246 34466 27298
rect 43822 27246 43874 27298
rect 46622 27246 46674 27298
rect 46958 27246 47010 27298
rect 47294 27246 47346 27298
rect 47742 27246 47794 27298
rect 49086 27246 49138 27298
rect 50654 27246 50706 27298
rect 52782 27246 52834 27298
rect 57150 27246 57202 27298
rect 4622 27134 4674 27186
rect 8542 27134 8594 27186
rect 15598 27134 15650 27186
rect 17278 27134 17330 27186
rect 26014 27134 26066 27186
rect 30942 27134 30994 27186
rect 31726 27134 31778 27186
rect 33854 27134 33906 27186
rect 35646 27134 35698 27186
rect 36318 27134 36370 27186
rect 37998 27134 38050 27186
rect 40014 27134 40066 27186
rect 42926 27134 42978 27186
rect 44942 27134 44994 27186
rect 52110 27134 52162 27186
rect 1710 27022 1762 27074
rect 5630 27022 5682 27074
rect 10894 27022 10946 27074
rect 11230 27022 11282 27074
rect 11790 27022 11842 27074
rect 15486 27022 15538 27074
rect 15710 27022 15762 27074
rect 16158 27022 16210 27074
rect 17838 27022 17890 27074
rect 18062 27022 18114 27074
rect 18398 27022 18450 27074
rect 18622 27022 18674 27074
rect 18846 27022 18898 27074
rect 19742 27022 19794 27074
rect 21982 27022 22034 27074
rect 22206 27022 22258 27074
rect 22542 27022 22594 27074
rect 22990 27022 23042 27074
rect 23662 27022 23714 27074
rect 24222 27022 24274 27074
rect 27470 27022 27522 27074
rect 31278 27022 31330 27074
rect 34078 27022 34130 27074
rect 34638 27022 34690 27074
rect 36094 27022 36146 27074
rect 37102 27022 37154 27074
rect 37326 27022 37378 27074
rect 39678 27022 39730 27074
rect 42030 27022 42082 27074
rect 42254 27022 42306 27074
rect 43262 27022 43314 27074
rect 43486 27022 43538 27074
rect 45390 27022 45442 27074
rect 46062 27022 46114 27074
rect 46286 27022 46338 27074
rect 47854 27022 47906 27074
rect 48526 27022 48578 27074
rect 51550 27022 51602 27074
rect 51886 27022 51938 27074
rect 55134 27022 55186 27074
rect 56030 27022 56082 27074
rect 57262 27022 57314 27074
rect 57486 27022 57538 27074
rect 2494 26910 2546 26962
rect 6414 26910 6466 26962
rect 9998 26910 10050 26962
rect 10334 26910 10386 26962
rect 11566 26910 11618 26962
rect 12014 26910 12066 26962
rect 12126 26910 12178 26962
rect 12686 26910 12738 26962
rect 16382 26910 16434 26962
rect 18174 26910 18226 26962
rect 19518 26910 19570 26962
rect 22654 26910 22706 26962
rect 22878 26910 22930 26962
rect 24334 26910 24386 26962
rect 26238 26910 26290 26962
rect 27918 26910 27970 26962
rect 29262 26910 29314 26962
rect 30494 26910 30546 26962
rect 32062 26910 32114 26962
rect 33294 26910 33346 26962
rect 34302 26910 34354 26962
rect 34862 26910 34914 26962
rect 34974 26910 35026 26962
rect 39790 26910 39842 26962
rect 40126 26910 40178 26962
rect 47182 26910 47234 26962
rect 47742 26910 47794 26962
rect 48190 26910 48242 26962
rect 49198 26910 49250 26962
rect 50542 26910 50594 26962
rect 10670 26798 10722 26850
rect 11230 26798 11282 26850
rect 16494 26798 16546 26850
rect 19182 26798 19234 26850
rect 21534 26798 21586 26850
rect 22318 26798 22370 26850
rect 24782 26798 24834 26850
rect 30046 26798 30098 26850
rect 32174 26798 32226 26850
rect 32398 26798 32450 26850
rect 32846 26798 32898 26850
rect 38894 26798 38946 26850
rect 48302 26798 48354 26850
rect 49086 26798 49138 26850
rect 49870 26798 49922 26850
rect 50654 26854 50706 26906
rect 52894 26910 52946 26962
rect 53342 26910 53394 26962
rect 53454 26910 53506 26962
rect 54126 26910 54178 26962
rect 54798 26910 54850 26962
rect 56702 26910 56754 26962
rect 52782 26798 52834 26850
rect 53678 26798 53730 26850
rect 15520 26630 15572 26682
rect 15624 26630 15676 26682
rect 15728 26630 15780 26682
rect 29827 26630 29879 26682
rect 29931 26630 29983 26682
rect 30035 26630 30087 26682
rect 44134 26630 44186 26682
rect 44238 26630 44290 26682
rect 44342 26630 44394 26682
rect 58441 26630 58493 26682
rect 58545 26630 58597 26682
rect 58649 26630 58701 26682
rect 2494 26462 2546 26514
rect 3054 26462 3106 26514
rect 6414 26462 6466 26514
rect 7198 26462 7250 26514
rect 8878 26462 8930 26514
rect 10446 26462 10498 26514
rect 24334 26462 24386 26514
rect 25230 26462 25282 26514
rect 30718 26462 30770 26514
rect 33406 26462 33458 26514
rect 33518 26462 33570 26514
rect 34526 26462 34578 26514
rect 35758 26462 35810 26514
rect 36206 26462 36258 26514
rect 36318 26462 36370 26514
rect 36766 26462 36818 26514
rect 39678 26462 39730 26514
rect 40798 26462 40850 26514
rect 45390 26462 45442 26514
rect 47518 26462 47570 26514
rect 2046 26350 2098 26402
rect 3502 26350 3554 26402
rect 4062 26350 4114 26402
rect 4622 26350 4674 26402
rect 8318 26350 8370 26402
rect 8990 26350 9042 26402
rect 10222 26350 10274 26402
rect 11454 26350 11506 26402
rect 20526 26350 20578 26402
rect 20638 26350 20690 26402
rect 23550 26350 23602 26402
rect 24558 26350 24610 26402
rect 28478 26350 28530 26402
rect 30942 26350 30994 26402
rect 33182 26350 33234 26402
rect 33742 26350 33794 26402
rect 34302 26350 34354 26402
rect 34862 26350 34914 26402
rect 35310 26350 35362 26402
rect 38334 26350 38386 26402
rect 40126 26350 40178 26402
rect 41022 26350 41074 26402
rect 44494 26350 44546 26402
rect 46622 26350 46674 26402
rect 49086 26350 49138 26402
rect 51662 26350 51714 26402
rect 52558 26350 52610 26402
rect 54798 26350 54850 26402
rect 55918 26350 55970 26402
rect 1822 26238 1874 26290
rect 2830 26238 2882 26290
rect 3278 26238 3330 26290
rect 3838 26238 3890 26290
rect 4174 26238 4226 26290
rect 4510 26238 4562 26290
rect 6078 26238 6130 26290
rect 6526 26238 6578 26290
rect 6750 26238 6802 26290
rect 7534 26238 7586 26290
rect 7982 26238 8034 26290
rect 8654 26238 8706 26290
rect 10110 26238 10162 26290
rect 10782 26238 10834 26290
rect 15038 26238 15090 26290
rect 16382 26238 16434 26290
rect 17950 26238 18002 26290
rect 18958 26238 19010 26290
rect 20302 26238 20354 26290
rect 21310 26238 21362 26290
rect 21534 26238 21586 26290
rect 21982 26238 22034 26290
rect 22654 26238 22706 26290
rect 22878 26238 22930 26290
rect 23774 26238 23826 26290
rect 24670 26238 24722 26290
rect 25566 26238 25618 26290
rect 29374 26238 29426 26290
rect 31054 26238 31106 26290
rect 31614 26238 31666 26290
rect 32398 26238 32450 26290
rect 33070 26238 33122 26290
rect 33854 26238 33906 26290
rect 34190 26238 34242 26290
rect 37102 26238 37154 26290
rect 38222 26238 38274 26290
rect 38558 26238 38610 26290
rect 40350 26238 40402 26290
rect 41134 26238 41186 26290
rect 44606 26238 44658 26290
rect 46062 26238 46114 26290
rect 46510 26238 46562 26290
rect 50430 26238 50482 26290
rect 53230 26238 53282 26290
rect 53454 26238 53506 26290
rect 55134 26238 55186 26290
rect 57150 26238 57202 26290
rect 9774 26126 9826 26178
rect 13582 26126 13634 26178
rect 16494 26126 16546 26178
rect 17726 26126 17778 26178
rect 21422 26126 21474 26178
rect 22318 26126 22370 26178
rect 27582 26126 27634 26178
rect 28478 26126 28530 26178
rect 37998 26126 38050 26178
rect 39118 26126 39170 26178
rect 40014 26126 40066 26178
rect 46958 26126 47010 26178
rect 47966 26126 48018 26178
rect 48974 26126 49026 26178
rect 52110 26126 52162 26178
rect 54910 26126 54962 26178
rect 55694 26126 55746 26178
rect 55806 26126 55858 26178
rect 56702 26126 56754 26178
rect 57598 26126 57650 26178
rect 58046 26126 58098 26178
rect 4622 26014 4674 26066
rect 14814 26014 14866 26066
rect 19182 26014 19234 26066
rect 23214 26014 23266 26066
rect 24110 26014 24162 26066
rect 36430 26014 36482 26066
rect 39342 26014 39394 26066
rect 44494 26014 44546 26066
rect 47182 26014 47234 26066
rect 8367 25846 8419 25898
rect 8471 25846 8523 25898
rect 8575 25846 8627 25898
rect 22674 25846 22726 25898
rect 22778 25846 22830 25898
rect 22882 25846 22934 25898
rect 36981 25846 37033 25898
rect 37085 25846 37137 25898
rect 37189 25846 37241 25898
rect 51288 25846 51340 25898
rect 51392 25846 51444 25898
rect 51496 25846 51548 25898
rect 8542 25678 8594 25730
rect 32062 25678 32114 25730
rect 33966 25678 34018 25730
rect 36990 25678 37042 25730
rect 46958 25678 47010 25730
rect 54014 25678 54066 25730
rect 4846 25566 4898 25618
rect 8206 25566 8258 25618
rect 12462 25566 12514 25618
rect 13694 25566 13746 25618
rect 16046 25566 16098 25618
rect 17166 25566 17218 25618
rect 18734 25566 18786 25618
rect 19630 25566 19682 25618
rect 23886 25566 23938 25618
rect 29598 25566 29650 25618
rect 31614 25566 31666 25618
rect 31950 25566 32002 25618
rect 34974 25566 35026 25618
rect 39454 25566 39506 25618
rect 41694 25566 41746 25618
rect 42478 25566 42530 25618
rect 45166 25566 45218 25618
rect 46174 25566 46226 25618
rect 47070 25566 47122 25618
rect 47742 25566 47794 25618
rect 49534 25566 49586 25618
rect 51662 25566 51714 25618
rect 53230 25566 53282 25618
rect 56030 25566 56082 25618
rect 56478 25566 56530 25618
rect 2046 25454 2098 25506
rect 11454 25454 11506 25506
rect 12014 25454 12066 25506
rect 14366 25454 14418 25506
rect 15598 25454 15650 25506
rect 15822 25454 15874 25506
rect 16382 25454 16434 25506
rect 19406 25454 19458 25506
rect 21758 25454 21810 25506
rect 26462 25454 26514 25506
rect 27918 25454 27970 25506
rect 29150 25454 29202 25506
rect 30046 25454 30098 25506
rect 30718 25454 30770 25506
rect 31166 25454 31218 25506
rect 33518 25454 33570 25506
rect 34190 25454 34242 25506
rect 34862 25454 34914 25506
rect 35646 25454 35698 25506
rect 38222 25454 38274 25506
rect 38558 25454 38610 25506
rect 39678 25454 39730 25506
rect 41134 25454 41186 25506
rect 42590 25454 42642 25506
rect 43150 25454 43202 25506
rect 43934 25454 43986 25506
rect 44718 25454 44770 25506
rect 45390 25454 45442 25506
rect 48638 25454 48690 25506
rect 49086 25454 49138 25506
rect 51214 25454 51266 25506
rect 51550 25454 51602 25506
rect 53678 25454 53730 25506
rect 55134 25454 55186 25506
rect 55918 25454 55970 25506
rect 57262 25454 57314 25506
rect 57710 25454 57762 25506
rect 2718 25342 2770 25394
rect 7646 25342 7698 25394
rect 7982 25342 8034 25394
rect 10334 25342 10386 25394
rect 10670 25342 10722 25394
rect 10894 25342 10946 25394
rect 11230 25342 11282 25394
rect 11678 25342 11730 25394
rect 11902 25342 11954 25394
rect 21646 25342 21698 25394
rect 27806 25342 27858 25394
rect 28030 25342 28082 25394
rect 29822 25342 29874 25394
rect 32958 25342 33010 25394
rect 33182 25342 33234 25394
rect 35870 25342 35922 25394
rect 37326 25342 37378 25394
rect 37774 25342 37826 25394
rect 37886 25342 37938 25394
rect 38334 25342 38386 25394
rect 38782 25342 38834 25394
rect 44270 25342 44322 25394
rect 46510 25342 46562 25394
rect 50094 25342 50146 25394
rect 54238 25342 54290 25394
rect 56142 25342 56194 25394
rect 9998 25230 10050 25282
rect 10446 25230 10498 25282
rect 11118 25230 11170 25282
rect 14030 25230 14082 25282
rect 16718 25230 16770 25282
rect 20190 25230 20242 25282
rect 21422 25230 21474 25282
rect 28702 25230 28754 25282
rect 32734 25230 32786 25282
rect 36430 25230 36482 25282
rect 37102 25230 37154 25282
rect 37550 25230 37602 25282
rect 38894 25230 38946 25282
rect 39118 25230 39170 25282
rect 44158 25230 44210 25282
rect 47182 25230 47234 25282
rect 48190 25230 48242 25282
rect 50206 25230 50258 25282
rect 50430 25230 50482 25282
rect 52110 25230 52162 25282
rect 53118 25230 53170 25282
rect 53342 25230 53394 25282
rect 54126 25230 54178 25282
rect 15520 25062 15572 25114
rect 15624 25062 15676 25114
rect 15728 25062 15780 25114
rect 29827 25062 29879 25114
rect 29931 25062 29983 25114
rect 30035 25062 30087 25114
rect 44134 25062 44186 25114
rect 44238 25062 44290 25114
rect 44342 25062 44394 25114
rect 58441 25062 58493 25114
rect 58545 25062 58597 25114
rect 58649 25062 58701 25114
rect 2158 24894 2210 24946
rect 3166 24894 3218 24946
rect 4846 24894 4898 24946
rect 22878 24894 22930 24946
rect 23662 24894 23714 24946
rect 23886 24894 23938 24946
rect 24110 24894 24162 24946
rect 27134 24894 27186 24946
rect 32286 24894 32338 24946
rect 42254 24894 42306 24946
rect 42590 24894 42642 24946
rect 3390 24782 3442 24834
rect 4062 24782 4114 24834
rect 4622 24782 4674 24834
rect 11118 24782 11170 24834
rect 17502 24782 17554 24834
rect 21422 24782 21474 24834
rect 22990 24782 23042 24834
rect 25230 24782 25282 24834
rect 29150 24782 29202 24834
rect 30494 24782 30546 24834
rect 34078 24782 34130 24834
rect 36766 24782 36818 24834
rect 36878 24782 36930 24834
rect 38110 24782 38162 24834
rect 38670 24782 38722 24834
rect 39230 24782 39282 24834
rect 41918 24782 41970 24834
rect 42814 24782 42866 24834
rect 44046 24782 44098 24834
rect 45502 24782 45554 24834
rect 45838 24782 45890 24834
rect 50542 24782 50594 24834
rect 51438 24782 51490 24834
rect 53454 24782 53506 24834
rect 55358 24782 55410 24834
rect 56590 24782 56642 24834
rect 2494 24670 2546 24722
rect 3054 24670 3106 24722
rect 3502 24670 3554 24722
rect 3950 24670 4002 24722
rect 4510 24670 4562 24722
rect 5742 24670 5794 24722
rect 10334 24670 10386 24722
rect 15486 24670 15538 24722
rect 15934 24670 15986 24722
rect 18286 24670 18338 24722
rect 19630 24670 19682 24722
rect 21646 24670 21698 24722
rect 23774 24670 23826 24722
rect 25342 24670 25394 24722
rect 25678 24670 25730 24722
rect 27582 24670 27634 24722
rect 29262 24670 29314 24722
rect 29822 24670 29874 24722
rect 31726 24670 31778 24722
rect 32174 24670 32226 24722
rect 32398 24670 32450 24722
rect 33182 24670 33234 24722
rect 33406 24670 33458 24722
rect 34862 24670 34914 24722
rect 35982 24670 36034 24722
rect 37102 24670 37154 24722
rect 38446 24670 38498 24722
rect 39118 24670 39170 24722
rect 40014 24670 40066 24722
rect 42142 24670 42194 24722
rect 42366 24670 42418 24722
rect 42926 24670 42978 24722
rect 43934 24670 43986 24722
rect 44270 24670 44322 24722
rect 44606 24670 44658 24722
rect 45054 24670 45106 24722
rect 47854 24670 47906 24722
rect 48638 24670 48690 24722
rect 49422 24670 49474 24722
rect 50430 24670 50482 24722
rect 50766 24670 50818 24722
rect 51326 24670 51378 24722
rect 51550 24670 51602 24722
rect 52222 24670 52274 24722
rect 54014 24670 54066 24722
rect 54686 24670 54738 24722
rect 56030 24670 56082 24722
rect 56814 24670 56866 24722
rect 57038 24670 57090 24722
rect 6526 24558 6578 24610
rect 8654 24558 8706 24610
rect 13358 24558 13410 24610
rect 15038 24558 15090 24610
rect 19742 24558 19794 24610
rect 27918 24558 27970 24610
rect 30942 24558 30994 24610
rect 31502 24558 31554 24610
rect 34414 24558 34466 24610
rect 36206 24558 36258 24610
rect 36318 24558 36370 24610
rect 37998 24558 38050 24610
rect 38782 24558 38834 24610
rect 39566 24558 39618 24610
rect 46398 24558 46450 24610
rect 47406 24558 47458 24610
rect 47630 24558 47682 24610
rect 48190 24558 48242 24610
rect 48862 24558 48914 24610
rect 49310 24558 49362 24610
rect 55806 24558 55858 24610
rect 58158 24558 58210 24610
rect 4062 24446 4114 24498
rect 28030 24446 28082 24498
rect 46062 24446 46114 24498
rect 55694 24446 55746 24498
rect 8367 24278 8419 24330
rect 8471 24278 8523 24330
rect 8575 24278 8627 24330
rect 22674 24278 22726 24330
rect 22778 24278 22830 24330
rect 22882 24278 22934 24330
rect 36981 24278 37033 24330
rect 37085 24278 37137 24330
rect 37189 24278 37241 24330
rect 51288 24278 51340 24330
rect 51392 24278 51444 24330
rect 51496 24278 51548 24330
rect 7534 24110 7586 24162
rect 18510 24110 18562 24162
rect 32510 24110 32562 24162
rect 42030 24110 42082 24162
rect 47854 24110 47906 24162
rect 51998 24110 52050 24162
rect 55246 24110 55298 24162
rect 55582 24110 55634 24162
rect 6638 23998 6690 24050
rect 9438 23998 9490 24050
rect 10222 23998 10274 24050
rect 16382 23998 16434 24050
rect 17726 23998 17778 24050
rect 17950 23998 18002 24050
rect 18286 23998 18338 24050
rect 19630 23998 19682 24050
rect 21422 23998 21474 24050
rect 27022 23998 27074 24050
rect 30158 23998 30210 24050
rect 33630 23998 33682 24050
rect 35534 23998 35586 24050
rect 37550 23998 37602 24050
rect 38446 23998 38498 24050
rect 40574 23998 40626 24050
rect 45278 23998 45330 24050
rect 46510 23998 46562 24050
rect 48526 23998 48578 24050
rect 51326 23998 51378 24050
rect 53342 23998 53394 24050
rect 2046 23886 2098 23938
rect 2382 23886 2434 23938
rect 3054 23886 3106 23938
rect 4062 23886 4114 23938
rect 6414 23886 6466 23938
rect 6862 23886 6914 23938
rect 7646 23886 7698 23938
rect 8206 23886 8258 23938
rect 10894 23886 10946 23938
rect 13470 23886 13522 23938
rect 19518 23886 19570 23938
rect 24334 23886 24386 23938
rect 24670 23886 24722 23938
rect 26126 23886 26178 23938
rect 26798 23886 26850 23938
rect 27806 23886 27858 23938
rect 28478 23886 28530 23938
rect 28590 23886 28642 23938
rect 29262 23886 29314 23938
rect 29486 23886 29538 23938
rect 30718 23886 30770 23938
rect 32062 23886 32114 23938
rect 32398 23886 32450 23938
rect 32958 23886 33010 23938
rect 34078 23886 34130 23938
rect 35870 23886 35922 23938
rect 37102 23886 37154 23938
rect 39902 23886 39954 23938
rect 41246 23886 41298 23938
rect 41694 23886 41746 23938
rect 42702 23886 42754 23938
rect 46062 23886 46114 23938
rect 48190 23886 48242 23938
rect 49086 23886 49138 23938
rect 49422 23886 49474 23938
rect 49758 23886 49810 23938
rect 50430 23886 50482 23938
rect 51662 23886 51714 23938
rect 52558 23886 52610 23938
rect 56814 23886 56866 23938
rect 57598 23886 57650 23938
rect 2606 23774 2658 23826
rect 3278 23774 3330 23826
rect 3390 23774 3442 23826
rect 4398 23774 4450 23826
rect 7086 23774 7138 23826
rect 7870 23774 7922 23826
rect 8094 23774 8146 23826
rect 10558 23774 10610 23826
rect 11342 23774 11394 23826
rect 11454 23774 11506 23826
rect 11902 23774 11954 23826
rect 12014 23774 12066 23826
rect 12574 23774 12626 23826
rect 14254 23774 14306 23826
rect 18846 23774 18898 23826
rect 19182 23774 19234 23826
rect 19742 23774 19794 23826
rect 21758 23774 21810 23826
rect 23326 23774 23378 23826
rect 25342 23774 25394 23826
rect 30494 23774 30546 23826
rect 33070 23774 33122 23826
rect 35198 23774 35250 23826
rect 39006 23774 39058 23826
rect 40910 23774 40962 23826
rect 41470 23774 41522 23826
rect 45726 23774 45778 23826
rect 45838 23774 45890 23826
rect 52894 23774 52946 23826
rect 56254 23774 56306 23826
rect 58158 23774 58210 23826
rect 2158 23662 2210 23714
rect 2718 23662 2770 23714
rect 2942 23662 2994 23714
rect 3726 23662 3778 23714
rect 3950 23662 4002 23714
rect 4510 23662 4562 23714
rect 4734 23662 4786 23714
rect 7534 23662 7586 23714
rect 11118 23662 11170 23714
rect 12238 23662 12290 23714
rect 17390 23662 17442 23714
rect 23214 23662 23266 23714
rect 24558 23662 24610 23714
rect 25230 23662 25282 23714
rect 25790 23662 25842 23714
rect 27582 23662 27634 23714
rect 27694 23662 27746 23714
rect 28030 23662 28082 23714
rect 34638 23662 34690 23714
rect 41022 23662 41074 23714
rect 42926 23662 42978 23714
rect 43598 23662 43650 23714
rect 44942 23662 44994 23714
rect 45166 23662 45218 23714
rect 45390 23662 45442 23714
rect 46846 23662 46898 23714
rect 47182 23662 47234 23714
rect 49310 23662 49362 23714
rect 49870 23662 49922 23714
rect 50094 23662 50146 23714
rect 50542 23662 50594 23714
rect 50766 23662 50818 23714
rect 52782 23662 52834 23714
rect 55358 23662 55410 23714
rect 15520 23494 15572 23546
rect 15624 23494 15676 23546
rect 15728 23494 15780 23546
rect 29827 23494 29879 23546
rect 29931 23494 29983 23546
rect 30035 23494 30087 23546
rect 44134 23494 44186 23546
rect 44238 23494 44290 23546
rect 44342 23494 44394 23546
rect 58441 23494 58493 23546
rect 58545 23494 58597 23546
rect 58649 23494 58701 23546
rect 8430 23326 8482 23378
rect 14030 23326 14082 23378
rect 15150 23326 15202 23378
rect 15710 23326 15762 23378
rect 16382 23326 16434 23378
rect 20638 23326 20690 23378
rect 28926 23326 28978 23378
rect 31390 23326 31442 23378
rect 32174 23326 32226 23378
rect 32398 23326 32450 23378
rect 33294 23326 33346 23378
rect 33966 23326 34018 23378
rect 35534 23326 35586 23378
rect 35870 23326 35922 23378
rect 37550 23326 37602 23378
rect 42814 23326 42866 23378
rect 43486 23326 43538 23378
rect 44718 23326 44770 23378
rect 47630 23326 47682 23378
rect 47966 23326 48018 23378
rect 50206 23326 50258 23378
rect 50990 23326 51042 23378
rect 23550 23214 23602 23266
rect 25902 23214 25954 23266
rect 26014 23214 26066 23266
rect 27358 23214 27410 23266
rect 27694 23214 27746 23266
rect 28030 23214 28082 23266
rect 28254 23214 28306 23266
rect 30494 23214 30546 23266
rect 31166 23214 31218 23266
rect 31614 23214 31666 23266
rect 31726 23214 31778 23266
rect 33518 23214 33570 23266
rect 34862 23214 34914 23266
rect 35310 23214 35362 23266
rect 35758 23214 35810 23266
rect 36766 23214 36818 23266
rect 37774 23214 37826 23266
rect 37886 23214 37938 23266
rect 39678 23214 39730 23266
rect 41470 23214 41522 23266
rect 45278 23214 45330 23266
rect 47406 23214 47458 23266
rect 50654 23214 50706 23266
rect 51550 23214 51602 23266
rect 55022 23214 55074 23266
rect 1822 23102 1874 23154
rect 5182 23102 5234 23154
rect 8766 23102 8818 23154
rect 9774 23102 9826 23154
rect 13694 23102 13746 23154
rect 14142 23102 14194 23154
rect 14254 23102 14306 23154
rect 14926 23102 14978 23154
rect 15262 23102 15314 23154
rect 15598 23102 15650 23154
rect 15934 23102 15986 23154
rect 17390 23102 17442 23154
rect 20862 23102 20914 23154
rect 24110 23102 24162 23154
rect 26686 23102 26738 23154
rect 29486 23102 29538 23154
rect 30830 23102 30882 23154
rect 32510 23102 32562 23154
rect 32958 23102 33010 23154
rect 34302 23102 34354 23154
rect 35198 23102 35250 23154
rect 36094 23102 36146 23154
rect 36430 23102 36482 23154
rect 39230 23102 39282 23154
rect 43262 23102 43314 23154
rect 43822 23102 43874 23154
rect 45166 23102 45218 23154
rect 45390 23102 45442 23154
rect 47294 23102 47346 23154
rect 48078 23102 48130 23154
rect 49086 23102 49138 23154
rect 51326 23102 51378 23154
rect 54350 23102 54402 23154
rect 54910 23102 54962 23154
rect 56926 23102 56978 23154
rect 2494 22990 2546 23042
rect 4622 22990 4674 23042
rect 5966 22990 6018 23042
rect 8094 22990 8146 23042
rect 10558 22990 10610 23042
rect 12686 22990 12738 23042
rect 13358 22990 13410 23042
rect 18174 22990 18226 23042
rect 20302 22990 20354 23042
rect 21982 22990 22034 23042
rect 24446 22990 24498 23042
rect 25566 22990 25618 23042
rect 26910 22990 26962 23042
rect 27806 22990 27858 23042
rect 30270 22990 30322 23042
rect 37214 22990 37266 23042
rect 38334 22990 38386 23042
rect 38782 22990 38834 23042
rect 41582 22990 41634 23042
rect 46062 22990 46114 23042
rect 46958 22990 47010 23042
rect 48190 22990 48242 23042
rect 48862 22990 48914 23042
rect 49758 22990 49810 23042
rect 52446 22990 52498 23042
rect 54798 22990 54850 23042
rect 56702 22990 56754 23042
rect 57598 22990 57650 23042
rect 25902 22878 25954 22930
rect 29262 22878 29314 22930
rect 33182 22878 33234 22930
rect 41694 22878 41746 22930
rect 44046 22878 44098 22930
rect 44382 22878 44434 22930
rect 51886 22878 51938 22930
rect 52222 22878 52274 22930
rect 8367 22710 8419 22762
rect 8471 22710 8523 22762
rect 8575 22710 8627 22762
rect 22674 22710 22726 22762
rect 22778 22710 22830 22762
rect 22882 22710 22934 22762
rect 36981 22710 37033 22762
rect 37085 22710 37137 22762
rect 37189 22710 37241 22762
rect 51288 22710 51340 22762
rect 51392 22710 51444 22762
rect 51496 22710 51548 22762
rect 7758 22542 7810 22594
rect 8094 22542 8146 22594
rect 27246 22542 27298 22594
rect 37774 22542 37826 22594
rect 38222 22542 38274 22594
rect 48526 22542 48578 22594
rect 55022 22542 55074 22594
rect 56142 22542 56194 22594
rect 3054 22430 3106 22482
rect 6078 22430 6130 22482
rect 11006 22430 11058 22482
rect 24110 22430 24162 22482
rect 25006 22430 25058 22482
rect 34750 22430 34802 22482
rect 35646 22430 35698 22482
rect 38782 22430 38834 22482
rect 39902 22430 39954 22482
rect 43262 22430 43314 22482
rect 54462 22430 54514 22482
rect 55918 22430 55970 22482
rect 2942 22318 2994 22370
rect 3278 22318 3330 22370
rect 3502 22318 3554 22370
rect 4510 22318 4562 22370
rect 6302 22318 6354 22370
rect 10894 22318 10946 22370
rect 11118 22318 11170 22370
rect 11678 22318 11730 22370
rect 13022 22318 13074 22370
rect 14030 22318 14082 22370
rect 14702 22318 14754 22370
rect 15038 22318 15090 22370
rect 15262 22318 15314 22370
rect 15710 22318 15762 22370
rect 16270 22318 16322 22370
rect 21534 22318 21586 22370
rect 22430 22318 22482 22370
rect 22878 22318 22930 22370
rect 25790 22318 25842 22370
rect 26126 22318 26178 22370
rect 26350 22318 26402 22370
rect 27358 22318 27410 22370
rect 27582 22318 27634 22370
rect 28366 22318 28418 22370
rect 28590 22318 28642 22370
rect 30158 22318 30210 22370
rect 30830 22318 30882 22370
rect 31166 22318 31218 22370
rect 32846 22318 32898 22370
rect 33406 22318 33458 22370
rect 33966 22318 34018 22370
rect 36206 22318 36258 22370
rect 37326 22318 37378 22370
rect 38334 22318 38386 22370
rect 41694 22318 41746 22370
rect 42590 22318 42642 22370
rect 44382 22318 44434 22370
rect 45166 22318 45218 22370
rect 45502 22318 45554 22370
rect 46510 22318 46562 22370
rect 49870 22318 49922 22370
rect 50430 22318 50482 22370
rect 50654 22318 50706 22370
rect 50990 22318 51042 22370
rect 51550 22318 51602 22370
rect 51886 22318 51938 22370
rect 52894 22318 52946 22370
rect 53230 22318 53282 22370
rect 54238 22318 54290 22370
rect 55806 22318 55858 22370
rect 57038 22318 57090 22370
rect 57262 22318 57314 22370
rect 2606 22206 2658 22258
rect 4174 22206 4226 22258
rect 5966 22206 6018 22258
rect 6526 22206 6578 22258
rect 7086 22206 7138 22258
rect 7422 22206 7474 22258
rect 8990 22206 9042 22258
rect 9326 22206 9378 22258
rect 10558 22206 10610 22258
rect 12686 22206 12738 22258
rect 13694 22206 13746 22258
rect 2270 22094 2322 22146
rect 9774 22094 9826 22146
rect 10334 22094 10386 22146
rect 11454 22094 11506 22146
rect 12350 22094 12402 22146
rect 12798 22094 12850 22146
rect 13806 22094 13858 22146
rect 14254 22150 14306 22202
rect 14590 22206 14642 22258
rect 15934 22206 15986 22258
rect 19406 22206 19458 22258
rect 22094 22206 22146 22258
rect 23102 22206 23154 22258
rect 23998 22206 24050 22258
rect 24894 22206 24946 22258
rect 29038 22206 29090 22258
rect 29374 22206 29426 22258
rect 29934 22206 29986 22258
rect 30606 22206 30658 22258
rect 31390 22206 31442 22258
rect 31502 22206 31554 22258
rect 32062 22206 32114 22258
rect 32622 22206 32674 22258
rect 33294 22206 33346 22258
rect 36990 22206 37042 22258
rect 37662 22206 37714 22258
rect 39454 22206 39506 22258
rect 40462 22206 40514 22258
rect 41358 22206 41410 22258
rect 44830 22206 44882 22258
rect 45838 22206 45890 22258
rect 46174 22206 46226 22258
rect 47406 22206 47458 22258
rect 48078 22206 48130 22258
rect 48526 22206 48578 22258
rect 48638 22206 48690 22258
rect 48974 22206 49026 22258
rect 49310 22206 49362 22258
rect 14366 22094 14418 22146
rect 15038 22094 15090 22146
rect 16158 22094 16210 22146
rect 16718 22094 16770 22146
rect 20302 22094 20354 22146
rect 21646 22094 21698 22146
rect 21870 22094 21922 22146
rect 24222 22094 24274 22146
rect 24446 22094 24498 22146
rect 25118 22094 25170 22146
rect 25342 22094 25394 22146
rect 25902 22094 25954 22146
rect 28030 22094 28082 22146
rect 32286 22094 32338 22146
rect 35310 22094 35362 22146
rect 38222 22094 38274 22146
rect 39118 22094 39170 22146
rect 39342 22094 39394 22146
rect 40574 22094 40626 22146
rect 40798 22094 40850 22146
rect 46286 22094 46338 22146
rect 47070 22094 47122 22146
rect 47742 22094 47794 22146
rect 49982 22094 50034 22146
rect 50206 22094 50258 22146
rect 51326 22094 51378 22146
rect 51438 22094 51490 22146
rect 57598 22094 57650 22146
rect 15520 21926 15572 21978
rect 15624 21926 15676 21978
rect 15728 21926 15780 21978
rect 29827 21926 29879 21978
rect 29931 21926 29983 21978
rect 30035 21926 30087 21978
rect 44134 21926 44186 21978
rect 44238 21926 44290 21978
rect 44342 21926 44394 21978
rect 58441 21926 58493 21978
rect 58545 21926 58597 21978
rect 58649 21926 58701 21978
rect 1934 21758 1986 21810
rect 2830 21758 2882 21810
rect 3166 21758 3218 21810
rect 4846 21758 4898 21810
rect 9998 21758 10050 21810
rect 14702 21758 14754 21810
rect 15262 21758 15314 21810
rect 18398 21758 18450 21810
rect 18958 21758 19010 21810
rect 22766 21758 22818 21810
rect 22990 21758 23042 21810
rect 25790 21758 25842 21810
rect 25902 21758 25954 21810
rect 26126 21758 26178 21810
rect 31614 21758 31666 21810
rect 32398 21758 32450 21810
rect 33630 21758 33682 21810
rect 33854 21758 33906 21810
rect 34414 21758 34466 21810
rect 37774 21758 37826 21810
rect 38110 21758 38162 21810
rect 39790 21758 39842 21810
rect 41246 21758 41298 21810
rect 46174 21758 46226 21810
rect 46846 21758 46898 21810
rect 51326 21758 51378 21810
rect 53678 21758 53730 21810
rect 54350 21758 54402 21810
rect 55694 21758 55746 21810
rect 57934 21758 57986 21810
rect 2158 21646 2210 21698
rect 2494 21646 2546 21698
rect 8654 21646 8706 21698
rect 10110 21646 10162 21698
rect 14030 21646 14082 21698
rect 14366 21646 14418 21698
rect 15486 21646 15538 21698
rect 15598 21646 15650 21698
rect 15934 21646 15986 21698
rect 16046 21646 16098 21698
rect 17502 21646 17554 21698
rect 18062 21646 18114 21698
rect 18510 21646 18562 21698
rect 19070 21646 19122 21698
rect 35422 21646 35474 21698
rect 36094 21646 36146 21698
rect 36878 21646 36930 21698
rect 38446 21646 38498 21698
rect 43822 21646 43874 21698
rect 44382 21646 44434 21698
rect 47406 21646 47458 21698
rect 47518 21646 47570 21698
rect 47966 21646 48018 21698
rect 48078 21646 48130 21698
rect 50654 21646 50706 21698
rect 50990 21646 51042 21698
rect 51102 21646 51154 21698
rect 51998 21646 52050 21698
rect 54462 21646 54514 21698
rect 55918 21646 55970 21698
rect 57262 21646 57314 21698
rect 4174 21534 4226 21586
rect 4622 21534 4674 21586
rect 8206 21534 8258 21586
rect 10446 21534 10498 21586
rect 14926 21534 14978 21586
rect 16606 21534 16658 21586
rect 19518 21534 19570 21586
rect 23438 21534 23490 21586
rect 26238 21534 26290 21586
rect 27246 21534 27298 21586
rect 28142 21534 28194 21586
rect 28590 21534 28642 21586
rect 29710 21534 29762 21586
rect 31950 21534 32002 21586
rect 32174 21534 32226 21586
rect 32510 21534 32562 21586
rect 33070 21534 33122 21586
rect 33406 21534 33458 21586
rect 34638 21534 34690 21586
rect 35086 21534 35138 21586
rect 36206 21534 36258 21586
rect 36766 21534 36818 21586
rect 37102 21534 37154 21586
rect 39118 21534 39170 21586
rect 40126 21534 40178 21586
rect 41022 21534 41074 21586
rect 41358 21534 41410 21586
rect 41582 21534 41634 21586
rect 42366 21534 42418 21586
rect 42926 21534 42978 21586
rect 44158 21534 44210 21586
rect 44494 21534 44546 21586
rect 45166 21534 45218 21586
rect 45838 21534 45890 21586
rect 45950 21534 46002 21586
rect 46286 21534 46338 21586
rect 46734 21534 46786 21586
rect 48302 21534 48354 21586
rect 49758 21534 49810 21586
rect 50430 21534 50482 21586
rect 52222 21534 52274 21586
rect 53118 21534 53170 21586
rect 57374 21534 57426 21586
rect 57822 21534 57874 21586
rect 4062 21422 4114 21474
rect 7758 21422 7810 21474
rect 11230 21422 11282 21474
rect 13358 21422 13410 21474
rect 20302 21422 20354 21474
rect 22430 21422 22482 21474
rect 22878 21422 22930 21474
rect 23774 21422 23826 21474
rect 26798 21422 26850 21474
rect 30270 21422 30322 21474
rect 33630 21422 33682 21474
rect 36318 21422 36370 21474
rect 37438 21422 37490 21474
rect 39342 21422 39394 21474
rect 44830 21422 44882 21474
rect 45390 21422 45442 21474
rect 46062 21422 46114 21474
rect 48862 21422 48914 21474
rect 55582 21422 55634 21474
rect 3838 21310 3890 21362
rect 8542 21310 8594 21362
rect 8878 21310 8930 21362
rect 9998 21310 10050 21362
rect 16046 21310 16098 21362
rect 18398 21310 18450 21362
rect 18958 21310 19010 21362
rect 46846 21310 46898 21362
rect 47518 21310 47570 21362
rect 54238 21310 54290 21362
rect 8367 21142 8419 21194
rect 8471 21142 8523 21194
rect 8575 21142 8627 21194
rect 22674 21142 22726 21194
rect 22778 21142 22830 21194
rect 22882 21142 22934 21194
rect 36981 21142 37033 21194
rect 37085 21142 37137 21194
rect 37189 21142 37241 21194
rect 51288 21142 51340 21194
rect 51392 21142 51444 21194
rect 51496 21142 51548 21194
rect 9102 20974 9154 21026
rect 9438 20974 9490 21026
rect 16270 20974 16322 21026
rect 20302 20974 20354 21026
rect 4622 20862 4674 20914
rect 8542 20862 8594 20914
rect 8878 20862 8930 20914
rect 10670 20862 10722 20914
rect 17390 20862 17442 20914
rect 19518 20862 19570 20914
rect 21870 20862 21922 20914
rect 26462 20862 26514 20914
rect 32062 20862 32114 20914
rect 32622 20862 32674 20914
rect 33854 20862 33906 20914
rect 34974 20862 35026 20914
rect 37438 20862 37490 20914
rect 41470 20862 41522 20914
rect 46398 20862 46450 20914
rect 48526 20862 48578 20914
rect 51550 20862 51602 20914
rect 53454 20862 53506 20914
rect 53902 20862 53954 20914
rect 57038 20862 57090 20914
rect 58046 20862 58098 20914
rect 1822 20762 1874 20814
rect 5630 20750 5682 20802
rect 10894 20750 10946 20802
rect 11342 20750 11394 20802
rect 11454 20750 11506 20802
rect 14142 20750 14194 20802
rect 14814 20750 14866 20802
rect 15038 20750 15090 20802
rect 15374 20750 15426 20802
rect 16270 20750 16322 20802
rect 16606 20750 16658 20802
rect 20078 20750 20130 20802
rect 20638 20750 20690 20802
rect 21982 20750 22034 20802
rect 28478 20750 28530 20802
rect 29150 20750 29202 20802
rect 30270 20750 30322 20802
rect 30494 20750 30546 20802
rect 31838 20750 31890 20802
rect 32734 20750 32786 20802
rect 33182 20750 33234 20802
rect 33518 20750 33570 20802
rect 36094 20750 36146 20802
rect 36318 20750 36370 20802
rect 36430 20750 36482 20802
rect 37326 20750 37378 20802
rect 38110 20750 38162 20802
rect 39454 20750 39506 20802
rect 40574 20750 40626 20802
rect 41246 20750 41298 20802
rect 41918 20750 41970 20802
rect 43934 20750 43986 20802
rect 46062 20750 46114 20802
rect 47182 20750 47234 20802
rect 47854 20750 47906 20802
rect 49310 20750 49362 20802
rect 49646 20750 49698 20802
rect 50318 20750 50370 20802
rect 50654 20750 50706 20802
rect 50878 20750 50930 20802
rect 53118 20750 53170 20802
rect 54126 20750 54178 20802
rect 55806 20750 55858 20802
rect 56926 20750 56978 20802
rect 2494 20638 2546 20690
rect 6414 20638 6466 20690
rect 12238 20638 12290 20690
rect 15934 20638 15986 20690
rect 19854 20638 19906 20690
rect 22654 20638 22706 20690
rect 29262 20638 29314 20690
rect 32174 20638 32226 20690
rect 35422 20638 35474 20690
rect 40014 20638 40066 20690
rect 40350 20638 40402 20690
rect 40910 20638 40962 20690
rect 41582 20638 41634 20690
rect 42030 20638 42082 20690
rect 44158 20638 44210 20690
rect 44942 20638 44994 20690
rect 46622 20638 46674 20690
rect 46734 20638 46786 20690
rect 47630 20638 47682 20690
rect 50990 20638 51042 20690
rect 52894 20638 52946 20690
rect 54798 20638 54850 20690
rect 55358 20638 55410 20690
rect 55470 20638 55522 20690
rect 56142 20638 56194 20690
rect 5070 20526 5122 20578
rect 11230 20526 11282 20578
rect 11902 20526 11954 20578
rect 12686 20526 12738 20578
rect 13694 20526 13746 20578
rect 14366 20526 14418 20578
rect 15038 20526 15090 20578
rect 20190 20526 20242 20578
rect 32510 20526 32562 20578
rect 34414 20526 34466 20578
rect 40798 20526 40850 20578
rect 47406 20526 47458 20578
rect 49198 20526 49250 20578
rect 49422 20526 49474 20578
rect 49534 20526 49586 20578
rect 50430 20526 50482 20578
rect 51214 20526 51266 20578
rect 51998 20526 52050 20578
rect 55694 20526 55746 20578
rect 56030 20526 56082 20578
rect 15520 20358 15572 20410
rect 15624 20358 15676 20410
rect 15728 20358 15780 20410
rect 29827 20358 29879 20410
rect 29931 20358 29983 20410
rect 30035 20358 30087 20410
rect 44134 20358 44186 20410
rect 44238 20358 44290 20410
rect 44342 20358 44394 20410
rect 58441 20358 58493 20410
rect 58545 20358 58597 20410
rect 58649 20358 58701 20410
rect 1934 20190 1986 20242
rect 3278 20190 3330 20242
rect 18510 20190 18562 20242
rect 19294 20190 19346 20242
rect 30494 20190 30546 20242
rect 31054 20190 31106 20242
rect 40798 20190 40850 20242
rect 50878 20190 50930 20242
rect 51326 20190 51378 20242
rect 54126 20190 54178 20242
rect 2270 20078 2322 20130
rect 3166 20078 3218 20130
rect 4622 20078 4674 20130
rect 4958 20078 5010 20130
rect 5630 20078 5682 20130
rect 8654 20078 8706 20130
rect 11678 20078 11730 20130
rect 14702 20078 14754 20130
rect 17502 20078 17554 20130
rect 17726 20078 17778 20130
rect 18174 20078 18226 20130
rect 19742 20078 19794 20130
rect 21758 20078 21810 20130
rect 24334 20078 24386 20130
rect 24670 20078 24722 20130
rect 26014 20078 26066 20130
rect 31390 20078 31442 20130
rect 34414 20078 34466 20130
rect 35982 20078 36034 20130
rect 37326 20078 37378 20130
rect 38670 20078 38722 20130
rect 39230 20078 39282 20130
rect 41022 20078 41074 20130
rect 42366 20078 42418 20130
rect 47854 20078 47906 20130
rect 50318 20078 50370 20130
rect 53006 20078 53058 20130
rect 53902 20078 53954 20130
rect 55694 20078 55746 20130
rect 55918 20078 55970 20130
rect 3502 19966 3554 20018
rect 3726 19966 3778 20018
rect 5294 19966 5346 20018
rect 8094 19966 8146 20018
rect 8318 19966 8370 20018
rect 10782 19966 10834 20018
rect 11454 19966 11506 20018
rect 12462 19966 12514 20018
rect 13918 19966 13970 20018
rect 18958 19966 19010 20018
rect 19406 19966 19458 20018
rect 22318 19966 22370 20018
rect 22990 19966 23042 20018
rect 23326 19966 23378 20018
rect 25230 19966 25282 20018
rect 28702 19966 28754 20018
rect 29374 19966 29426 20018
rect 30158 19966 30210 20018
rect 33182 19966 33234 20018
rect 34638 19966 34690 20018
rect 35310 19966 35362 20018
rect 36430 19966 36482 20018
rect 36654 19966 36706 20018
rect 37662 19966 37714 20018
rect 38222 19966 38274 20018
rect 38446 19966 38498 20018
rect 38782 19966 38834 20018
rect 39678 19966 39730 20018
rect 41134 19966 41186 20018
rect 42030 19966 42082 20018
rect 43822 19966 43874 20018
rect 44494 19966 44546 20018
rect 46622 19966 46674 20018
rect 48078 19966 48130 20018
rect 48750 19966 48802 20018
rect 48974 19966 49026 20018
rect 49086 19966 49138 20018
rect 49534 19966 49586 20018
rect 49758 19966 49810 20018
rect 50206 19966 50258 20018
rect 50542 19966 50594 20018
rect 52446 19966 52498 20018
rect 52894 19966 52946 20018
rect 53118 19966 53170 20018
rect 56030 19966 56082 20018
rect 56702 19966 56754 20018
rect 57038 19966 57090 20018
rect 2606 19854 2658 19906
rect 6190 19854 6242 19906
rect 6638 19854 6690 19906
rect 7198 19854 7250 19906
rect 9886 19854 9938 19906
rect 10334 19854 10386 19906
rect 10558 19854 10610 19906
rect 11118 19854 11170 19906
rect 11790 19854 11842 19906
rect 12910 19854 12962 19906
rect 13694 19854 13746 19906
rect 16830 19854 16882 19906
rect 20190 19854 20242 19906
rect 20974 19854 21026 19906
rect 28142 19854 28194 19906
rect 28590 19854 28642 19906
rect 29934 19854 29986 19906
rect 32510 19854 32562 19906
rect 40126 19854 40178 19906
rect 41806 19854 41858 19906
rect 43374 19854 43426 19906
rect 44718 19854 44770 19906
rect 46062 19854 46114 19906
rect 51774 19854 51826 19906
rect 54238 19854 54290 19906
rect 56590 19854 56642 19906
rect 2718 19742 2770 19794
rect 3726 19742 3778 19794
rect 6862 19742 6914 19794
rect 7198 19742 7250 19794
rect 8878 19742 8930 19794
rect 9102 19742 9154 19794
rect 17838 19742 17890 19794
rect 19182 19742 19234 19794
rect 31950 19742 32002 19794
rect 32286 19742 32338 19794
rect 33070 19742 33122 19794
rect 50766 19742 50818 19794
rect 51774 19742 51826 19794
rect 8367 19574 8419 19626
rect 8471 19574 8523 19626
rect 8575 19574 8627 19626
rect 22674 19574 22726 19626
rect 22778 19574 22830 19626
rect 22882 19574 22934 19626
rect 36981 19574 37033 19626
rect 37085 19574 37137 19626
rect 37189 19574 37241 19626
rect 51288 19574 51340 19626
rect 51392 19574 51444 19626
rect 51496 19574 51548 19626
rect 8542 19406 8594 19458
rect 8990 19406 9042 19458
rect 11454 19406 11506 19458
rect 16830 19406 16882 19458
rect 17390 19406 17442 19458
rect 21646 19406 21698 19458
rect 23438 19406 23490 19458
rect 32734 19406 32786 19458
rect 34414 19406 34466 19458
rect 43934 19406 43986 19458
rect 52110 19406 52162 19458
rect 53230 19406 53282 19458
rect 53566 19406 53618 19458
rect 53902 19406 53954 19458
rect 57486 19406 57538 19458
rect 4622 19294 4674 19346
rect 7198 19294 7250 19346
rect 9998 19294 10050 19346
rect 11678 19294 11730 19346
rect 16830 19294 16882 19346
rect 19854 19294 19906 19346
rect 22766 19294 22818 19346
rect 23998 19294 24050 19346
rect 24446 19294 24498 19346
rect 24894 19294 24946 19346
rect 25454 19294 25506 19346
rect 28590 19294 28642 19346
rect 29262 19294 29314 19346
rect 30270 19294 30322 19346
rect 30606 19294 30658 19346
rect 31502 19294 31554 19346
rect 31950 19294 32002 19346
rect 32846 19294 32898 19346
rect 34078 19294 34130 19346
rect 35982 19294 36034 19346
rect 37998 19294 38050 19346
rect 40126 19294 40178 19346
rect 40686 19294 40738 19346
rect 42030 19294 42082 19346
rect 45166 19294 45218 19346
rect 50206 19294 50258 19346
rect 51550 19294 51602 19346
rect 52670 19294 52722 19346
rect 55022 19294 55074 19346
rect 56254 19294 56306 19346
rect 56926 19294 56978 19346
rect 1710 19182 1762 19234
rect 5742 19182 5794 19234
rect 6526 19182 6578 19234
rect 6862 19182 6914 19234
rect 8094 19182 8146 19234
rect 9214 19182 9266 19234
rect 9438 19182 9490 19234
rect 10670 19182 10722 19234
rect 11118 19182 11170 19234
rect 11566 19182 11618 19234
rect 12574 19182 12626 19234
rect 13470 19182 13522 19234
rect 13806 19182 13858 19234
rect 14030 19182 14082 19234
rect 17278 19182 17330 19234
rect 19070 19182 19122 19234
rect 19518 19182 19570 19234
rect 20078 19182 20130 19234
rect 22878 19182 22930 19234
rect 23774 19182 23826 19234
rect 25790 19182 25842 19234
rect 26462 19182 26514 19234
rect 28142 19182 28194 19234
rect 28478 19182 28530 19234
rect 29038 19182 29090 19234
rect 31278 19182 31330 19234
rect 33070 19182 33122 19234
rect 33854 19182 33906 19234
rect 35310 19182 35362 19234
rect 35758 19182 35810 19234
rect 36206 19182 36258 19234
rect 37214 19182 37266 19234
rect 41134 19182 41186 19234
rect 42254 19182 42306 19234
rect 43262 19182 43314 19234
rect 47854 19182 47906 19234
rect 48190 19182 48242 19234
rect 48862 19182 48914 19234
rect 49534 19182 49586 19234
rect 50766 19182 50818 19234
rect 51774 19182 51826 19234
rect 52894 19182 52946 19234
rect 55134 19182 55186 19234
rect 55470 19182 55522 19234
rect 55694 19182 55746 19234
rect 56814 19182 56866 19234
rect 2494 19070 2546 19122
rect 6078 19070 6130 19122
rect 6302 19070 6354 19122
rect 7534 19070 7586 19122
rect 8318 19070 8370 19122
rect 9886 19070 9938 19122
rect 10334 19070 10386 19122
rect 10446 19070 10498 19122
rect 12798 19070 12850 19122
rect 14590 19070 14642 19122
rect 14702 19070 14754 19122
rect 15822 19070 15874 19122
rect 17614 19070 17666 19122
rect 26910 19070 26962 19122
rect 29486 19070 29538 19122
rect 29710 19070 29762 19122
rect 34638 19070 34690 19122
rect 36430 19070 36482 19122
rect 46286 19070 46338 19122
rect 46622 19070 46674 19122
rect 46958 19070 47010 19122
rect 47294 19070 47346 19122
rect 47406 19070 47458 19122
rect 47966 19070 48018 19122
rect 49758 19070 49810 19122
rect 50878 19070 50930 19122
rect 53790 19070 53842 19122
rect 54798 19070 54850 19122
rect 5070 18958 5122 19010
rect 6414 18958 6466 19010
rect 7310 18958 7362 19010
rect 13918 18958 13970 19010
rect 14366 18958 14418 19010
rect 15486 18958 15538 19010
rect 15934 18958 15986 19010
rect 16158 18958 16210 19010
rect 17726 18958 17778 19010
rect 17950 18958 18002 19010
rect 18734 18958 18786 19010
rect 20414 18958 20466 19010
rect 26126 18958 26178 19010
rect 26350 18958 26402 19010
rect 35534 18958 35586 19010
rect 41358 18958 41410 19010
rect 45726 18958 45778 19010
rect 45950 18958 46002 19010
rect 47630 18958 47682 19010
rect 49086 18958 49138 19010
rect 51102 18958 51154 19010
rect 15520 18790 15572 18842
rect 15624 18790 15676 18842
rect 15728 18790 15780 18842
rect 29827 18790 29879 18842
rect 29931 18790 29983 18842
rect 30035 18790 30087 18842
rect 44134 18790 44186 18842
rect 44238 18790 44290 18842
rect 44342 18790 44394 18842
rect 58441 18790 58493 18842
rect 58545 18790 58597 18842
rect 58649 18790 58701 18842
rect 2046 18622 2098 18674
rect 3054 18622 3106 18674
rect 3502 18622 3554 18674
rect 4510 18622 4562 18674
rect 8654 18622 8706 18674
rect 12126 18622 12178 18674
rect 13694 18622 13746 18674
rect 24446 18622 24498 18674
rect 24670 18622 24722 18674
rect 30046 18622 30098 18674
rect 33294 18622 33346 18674
rect 33966 18622 34018 18674
rect 34190 18622 34242 18674
rect 36318 18622 36370 18674
rect 37774 18622 37826 18674
rect 38782 18622 38834 18674
rect 41470 18622 41522 18674
rect 42702 18622 42754 18674
rect 47854 18622 47906 18674
rect 50542 18622 50594 18674
rect 51102 18622 51154 18674
rect 3390 18510 3442 18562
rect 3614 18510 3666 18562
rect 5182 18510 5234 18562
rect 5854 18510 5906 18562
rect 6862 18510 6914 18562
rect 8542 18510 8594 18562
rect 13022 18510 13074 18562
rect 13470 18510 13522 18562
rect 14702 18510 14754 18562
rect 19742 18510 19794 18562
rect 21198 18510 21250 18562
rect 22766 18510 22818 18562
rect 26686 18510 26738 18562
rect 28590 18510 28642 18562
rect 30942 18510 30994 18562
rect 31054 18510 31106 18562
rect 31502 18510 31554 18562
rect 34862 18510 34914 18562
rect 34974 18510 35026 18562
rect 37886 18510 37938 18562
rect 46510 18510 46562 18562
rect 47182 18510 47234 18562
rect 49982 18510 50034 18562
rect 50430 18510 50482 18562
rect 51998 18510 52050 18562
rect 1822 18398 1874 18450
rect 2830 18398 2882 18450
rect 4174 18398 4226 18450
rect 4846 18398 4898 18450
rect 5518 18398 5570 18450
rect 6190 18398 6242 18450
rect 6526 18398 6578 18450
rect 7646 18398 7698 18450
rect 8206 18398 8258 18450
rect 8878 18398 8930 18450
rect 10222 18398 10274 18450
rect 10334 18398 10386 18450
rect 11230 18398 11282 18450
rect 11678 18398 11730 18450
rect 12686 18398 12738 18450
rect 13358 18398 13410 18450
rect 13918 18398 13970 18450
rect 17950 18398 18002 18450
rect 18510 18398 18562 18450
rect 18846 18398 18898 18450
rect 19294 18398 19346 18450
rect 20414 18398 20466 18450
rect 21086 18398 21138 18450
rect 21422 18398 21474 18450
rect 22206 18398 22258 18450
rect 23102 18398 23154 18450
rect 23662 18398 23714 18450
rect 24110 18398 24162 18450
rect 24782 18398 24834 18450
rect 25902 18398 25954 18450
rect 26126 18398 26178 18450
rect 26462 18398 26514 18450
rect 26798 18398 26850 18450
rect 27918 18398 27970 18450
rect 28366 18398 28418 18450
rect 29150 18398 29202 18450
rect 29262 18398 29314 18450
rect 29374 18398 29426 18450
rect 29822 18398 29874 18450
rect 31278 18398 31330 18450
rect 32174 18398 32226 18450
rect 32398 18398 32450 18450
rect 33070 18398 33122 18450
rect 33182 18398 33234 18450
rect 33630 18398 33682 18450
rect 33854 18398 33906 18450
rect 34414 18398 34466 18450
rect 34638 18398 34690 18450
rect 36766 18398 36818 18450
rect 37102 18398 37154 18450
rect 37326 18398 37378 18450
rect 37550 18398 37602 18450
rect 40462 18398 40514 18450
rect 41806 18398 41858 18450
rect 42030 18398 42082 18450
rect 42366 18398 42418 18450
rect 43822 18398 43874 18450
rect 44382 18398 44434 18450
rect 44718 18398 44770 18450
rect 46286 18398 46338 18450
rect 46846 18398 46898 18450
rect 47518 18398 47570 18450
rect 48974 18398 49026 18450
rect 49870 18398 49922 18450
rect 50206 18398 50258 18450
rect 50766 18398 50818 18450
rect 53006 18398 53058 18450
rect 55134 18398 55186 18450
rect 56030 18398 56082 18450
rect 57150 18398 57202 18450
rect 7310 18286 7362 18338
rect 10670 18286 10722 18338
rect 16830 18286 16882 18338
rect 17614 18286 17666 18338
rect 19630 18286 19682 18338
rect 21982 18286 22034 18338
rect 25230 18286 25282 18338
rect 30382 18286 30434 18338
rect 30606 18286 30658 18338
rect 35534 18286 35586 18338
rect 35870 18286 35922 18338
rect 37214 18286 37266 18338
rect 38334 18286 38386 18338
rect 41022 18286 41074 18338
rect 44158 18286 44210 18338
rect 45166 18286 45218 18338
rect 45726 18286 45778 18338
rect 49534 18286 49586 18338
rect 51550 18286 51602 18338
rect 53678 18286 53730 18338
rect 55582 18286 55634 18338
rect 56814 18286 56866 18338
rect 3950 18174 4002 18226
rect 9774 18174 9826 18226
rect 11454 18174 11506 18226
rect 40798 18174 40850 18226
rect 41022 18174 41074 18226
rect 56702 18174 56754 18226
rect 8367 18006 8419 18058
rect 8471 18006 8523 18058
rect 8575 18006 8627 18058
rect 22674 18006 22726 18058
rect 22778 18006 22830 18058
rect 22882 18006 22934 18058
rect 36981 18006 37033 18058
rect 37085 18006 37137 18058
rect 37189 18006 37241 18058
rect 51288 18006 51340 18058
rect 51392 18006 51444 18058
rect 51496 18006 51548 18058
rect 10334 17838 10386 17890
rect 10558 17838 10610 17890
rect 16606 17838 16658 17890
rect 30718 17838 30770 17890
rect 34974 17838 35026 17890
rect 35310 17838 35362 17890
rect 35758 17838 35810 17890
rect 50542 17838 50594 17890
rect 53342 17838 53394 17890
rect 55582 17838 55634 17890
rect 55918 17838 55970 17890
rect 4062 17726 4114 17778
rect 11902 17726 11954 17778
rect 12910 17726 12962 17778
rect 16158 17726 16210 17778
rect 17278 17726 17330 17778
rect 18622 17726 18674 17778
rect 20190 17726 20242 17778
rect 28030 17726 28082 17778
rect 30046 17726 30098 17778
rect 32286 17726 32338 17778
rect 33966 17726 34018 17778
rect 37102 17726 37154 17778
rect 40350 17726 40402 17778
rect 41470 17726 41522 17778
rect 43934 17726 43986 17778
rect 49310 17726 49362 17778
rect 51774 17726 51826 17778
rect 55246 17726 55298 17778
rect 56702 17726 56754 17778
rect 57822 17726 57874 17778
rect 1710 17614 1762 17666
rect 2606 17614 2658 17666
rect 4286 17614 4338 17666
rect 5854 17614 5906 17666
rect 6414 17614 6466 17666
rect 7086 17614 7138 17666
rect 7534 17614 7586 17666
rect 8542 17614 8594 17666
rect 9662 17614 9714 17666
rect 10110 17614 10162 17666
rect 11790 17614 11842 17666
rect 12126 17614 12178 17666
rect 12574 17614 12626 17666
rect 13470 17614 13522 17666
rect 14030 17614 14082 17666
rect 14478 17614 14530 17666
rect 14926 17614 14978 17666
rect 17726 17614 17778 17666
rect 19294 17614 19346 17666
rect 19518 17614 19570 17666
rect 20526 17614 20578 17666
rect 20862 17614 20914 17666
rect 26574 17614 26626 17666
rect 27358 17614 27410 17666
rect 27918 17614 27970 17666
rect 29150 17614 29202 17666
rect 29598 17614 29650 17666
rect 30830 17614 30882 17666
rect 31278 17614 31330 17666
rect 31614 17614 31666 17666
rect 32734 17614 32786 17666
rect 33182 17614 33234 17666
rect 34750 17614 34802 17666
rect 35534 17614 35586 17666
rect 36318 17614 36370 17666
rect 37550 17614 37602 17666
rect 38222 17614 38274 17666
rect 42926 17614 42978 17666
rect 45614 17614 45666 17666
rect 45950 17614 46002 17666
rect 48750 17614 48802 17666
rect 49534 17614 49586 17666
rect 50766 17614 50818 17666
rect 51102 17614 51154 17666
rect 53118 17614 53170 17666
rect 53342 17614 53394 17666
rect 54462 17614 54514 17666
rect 54910 17614 54962 17666
rect 55582 17614 55634 17666
rect 56926 17614 56978 17666
rect 2046 17502 2098 17554
rect 2382 17502 2434 17554
rect 3950 17502 4002 17554
rect 4958 17502 5010 17554
rect 9438 17502 9490 17554
rect 13582 17502 13634 17554
rect 14702 17502 14754 17554
rect 15150 17502 15202 17554
rect 15262 17502 15314 17554
rect 15822 17502 15874 17554
rect 16046 17502 16098 17554
rect 16494 17502 16546 17554
rect 16606 17502 16658 17554
rect 20638 17502 20690 17554
rect 21534 17502 21586 17554
rect 30606 17502 30658 17554
rect 34190 17502 34242 17554
rect 42030 17502 42082 17554
rect 44830 17502 44882 17554
rect 46510 17502 46562 17554
rect 47854 17502 47906 17554
rect 49086 17502 49138 17554
rect 54686 17502 54738 17554
rect 56254 17502 56306 17554
rect 57710 17502 57762 17554
rect 3166 17390 3218 17442
rect 3726 17390 3778 17442
rect 4622 17390 4674 17442
rect 5630 17390 5682 17442
rect 7758 17390 7810 17442
rect 9102 17390 9154 17442
rect 11006 17390 11058 17442
rect 13806 17390 13858 17442
rect 14366 17390 14418 17442
rect 17838 17390 17890 17442
rect 18062 17390 18114 17442
rect 31054 17390 31106 17442
rect 31502 17390 31554 17442
rect 34414 17390 34466 17442
rect 34638 17390 34690 17442
rect 35870 17390 35922 17442
rect 36094 17390 36146 17442
rect 45166 17390 45218 17442
rect 45726 17390 45778 17442
rect 46846 17390 46898 17442
rect 47518 17390 47570 17442
rect 48414 17390 48466 17442
rect 48862 17390 48914 17442
rect 49870 17390 49922 17442
rect 50206 17390 50258 17442
rect 51214 17390 51266 17442
rect 51438 17390 51490 17442
rect 57934 17390 57986 17442
rect 15520 17222 15572 17274
rect 15624 17222 15676 17274
rect 15728 17222 15780 17274
rect 29827 17222 29879 17274
rect 29931 17222 29983 17274
rect 30035 17222 30087 17274
rect 44134 17222 44186 17274
rect 44238 17222 44290 17274
rect 44342 17222 44394 17274
rect 58441 17222 58493 17274
rect 58545 17222 58597 17274
rect 58649 17222 58701 17274
rect 2046 17054 2098 17106
rect 6414 17054 6466 17106
rect 11454 17054 11506 17106
rect 12798 17054 12850 17106
rect 13022 17054 13074 17106
rect 13358 17054 13410 17106
rect 14030 17054 14082 17106
rect 14366 17054 14418 17106
rect 20862 17054 20914 17106
rect 24222 17054 24274 17106
rect 24446 17054 24498 17106
rect 30270 17054 30322 17106
rect 31390 17054 31442 17106
rect 32174 17054 32226 17106
rect 33070 17054 33122 17106
rect 33630 17054 33682 17106
rect 34750 17054 34802 17106
rect 35086 17054 35138 17106
rect 35646 17054 35698 17106
rect 42366 17054 42418 17106
rect 43150 17054 43202 17106
rect 45278 17054 45330 17106
rect 45950 17054 46002 17106
rect 47742 17054 47794 17106
rect 50430 17054 50482 17106
rect 55918 17054 55970 17106
rect 2382 16942 2434 16994
rect 2718 16942 2770 16994
rect 3838 16942 3890 16994
rect 8318 16942 8370 16994
rect 9550 16942 9602 16994
rect 10894 16942 10946 16994
rect 12686 16942 12738 16994
rect 15262 16942 15314 16994
rect 15710 16942 15762 16994
rect 16830 16942 16882 16994
rect 18174 16942 18226 16994
rect 20974 16942 21026 16994
rect 21310 16942 21362 16994
rect 29038 16942 29090 16994
rect 30494 16942 30546 16994
rect 30606 16942 30658 16994
rect 31726 16942 31778 16994
rect 33406 16942 33458 16994
rect 33854 16942 33906 16994
rect 35982 16942 36034 16994
rect 41246 16942 41298 16994
rect 43038 16942 43090 16994
rect 43598 16942 43650 16994
rect 43934 16942 43986 16994
rect 45614 16942 45666 16994
rect 46958 16942 47010 16994
rect 47294 16942 47346 16994
rect 1710 16830 1762 16882
rect 3054 16830 3106 16882
rect 7758 16830 7810 16882
rect 8542 16830 8594 16882
rect 8766 16830 8818 16882
rect 12014 16830 12066 16882
rect 13470 16830 13522 16882
rect 14702 16830 14754 16882
rect 15038 16830 15090 16882
rect 16270 16830 16322 16882
rect 16606 16830 16658 16882
rect 17502 16830 17554 16882
rect 20638 16830 20690 16882
rect 21758 16830 21810 16882
rect 22206 16830 22258 16882
rect 22654 16830 22706 16882
rect 23102 16830 23154 16882
rect 24782 16830 24834 16882
rect 25678 16830 25730 16882
rect 27358 16830 27410 16882
rect 28366 16830 28418 16882
rect 29486 16830 29538 16882
rect 32398 16830 32450 16882
rect 33966 16830 34018 16882
rect 34414 16830 34466 16882
rect 35870 16830 35922 16882
rect 36206 16830 36258 16882
rect 36430 16830 36482 16882
rect 36654 16830 36706 16882
rect 36878 16830 36930 16882
rect 37102 16830 37154 16882
rect 37438 16830 37490 16882
rect 38110 16830 38162 16882
rect 41134 16830 41186 16882
rect 41470 16830 41522 16882
rect 42702 16830 42754 16882
rect 43374 16830 43426 16882
rect 46174 16830 46226 16882
rect 47630 16830 47682 16882
rect 48974 16830 49026 16882
rect 49198 16830 49250 16882
rect 49646 16830 49698 16882
rect 51214 16830 51266 16882
rect 52782 16830 52834 16882
rect 54686 16830 54738 16882
rect 55134 16830 55186 16882
rect 56814 16830 56866 16882
rect 57150 16830 57202 16882
rect 5966 16718 6018 16770
rect 6974 16718 7026 16770
rect 7646 16718 7698 16770
rect 9774 16718 9826 16770
rect 11006 16718 11058 16770
rect 11118 16718 11170 16770
rect 15150 16718 15202 16770
rect 16718 16718 16770 16770
rect 20302 16718 20354 16770
rect 23438 16718 23490 16770
rect 24558 16718 24610 16770
rect 25342 16718 25394 16770
rect 25566 16718 25618 16770
rect 27806 16718 27858 16770
rect 29934 16718 29986 16770
rect 40238 16718 40290 16770
rect 49086 16718 49138 16770
rect 49982 16718 50034 16770
rect 51438 16718 51490 16770
rect 51886 16718 51938 16770
rect 53118 16718 53170 16770
rect 53566 16718 53618 16770
rect 54350 16718 54402 16770
rect 55694 16718 55746 16770
rect 56030 16718 56082 16770
rect 8206 16606 8258 16658
rect 10110 16606 10162 16658
rect 13358 16606 13410 16658
rect 16270 16606 16322 16658
rect 27358 16606 27410 16658
rect 47742 16606 47794 16658
rect 56926 16606 56978 16658
rect 8367 16438 8419 16490
rect 8471 16438 8523 16490
rect 8575 16438 8627 16490
rect 22674 16438 22726 16490
rect 22778 16438 22830 16490
rect 22882 16438 22934 16490
rect 36981 16438 37033 16490
rect 37085 16438 37137 16490
rect 37189 16438 37241 16490
rect 51288 16438 51340 16490
rect 51392 16438 51444 16490
rect 51496 16438 51548 16490
rect 12686 16270 12738 16322
rect 24782 16270 24834 16322
rect 27358 16270 27410 16322
rect 28366 16270 28418 16322
rect 42366 16270 42418 16322
rect 48974 16270 49026 16322
rect 49870 16270 49922 16322
rect 50990 16270 51042 16322
rect 51326 16270 51378 16322
rect 55582 16270 55634 16322
rect 2494 16158 2546 16210
rect 4622 16158 4674 16210
rect 6974 16158 7026 16210
rect 9774 16158 9826 16210
rect 14366 16158 14418 16210
rect 15598 16158 15650 16210
rect 17726 16158 17778 16210
rect 19630 16158 19682 16210
rect 21758 16158 21810 16210
rect 25118 16158 25170 16210
rect 27582 16158 27634 16210
rect 29374 16158 29426 16210
rect 31278 16158 31330 16210
rect 34414 16158 34466 16210
rect 34974 16158 35026 16210
rect 35310 16158 35362 16210
rect 38110 16158 38162 16210
rect 38894 16158 38946 16210
rect 42478 16158 42530 16210
rect 43262 16158 43314 16210
rect 44158 16158 44210 16210
rect 48414 16158 48466 16210
rect 49310 16158 49362 16210
rect 50878 16158 50930 16210
rect 51326 16158 51378 16210
rect 51774 16158 51826 16210
rect 53006 16158 53058 16210
rect 56030 16158 56082 16210
rect 1822 16046 1874 16098
rect 6302 16046 6354 16098
rect 7198 16046 7250 16098
rect 8542 16046 8594 16098
rect 8990 16046 9042 16098
rect 10782 16046 10834 16098
rect 11342 16046 11394 16098
rect 12014 16046 12066 16098
rect 12574 16046 12626 16098
rect 14926 16046 14978 16098
rect 18286 16046 18338 16098
rect 20526 16046 20578 16098
rect 20862 16046 20914 16098
rect 23326 16046 23378 16098
rect 25342 16046 25394 16098
rect 27694 16046 27746 16098
rect 28254 16046 28306 16098
rect 29710 16046 29762 16098
rect 30046 16046 30098 16098
rect 30382 16046 30434 16098
rect 30830 16046 30882 16098
rect 32286 16046 32338 16098
rect 33182 16046 33234 16098
rect 36206 16046 36258 16098
rect 36990 16046 37042 16098
rect 37662 16046 37714 16098
rect 39902 16046 39954 16098
rect 40462 16046 40514 16098
rect 42254 16046 42306 16098
rect 43486 16046 43538 16098
rect 45278 16046 45330 16098
rect 45726 16046 45778 16098
rect 46174 16046 46226 16098
rect 46510 16046 46562 16098
rect 47070 16046 47122 16098
rect 47854 16046 47906 16098
rect 48190 16046 48242 16098
rect 48638 16046 48690 16098
rect 49534 16046 49586 16098
rect 50094 16046 50146 16098
rect 55582 16046 55634 16098
rect 5070 15934 5122 15986
rect 8094 15934 8146 15986
rect 8766 15934 8818 15986
rect 9214 15934 9266 15986
rect 9326 15934 9378 15986
rect 10558 15934 10610 15986
rect 12238 15934 12290 15986
rect 12686 15934 12738 15986
rect 18398 15934 18450 15986
rect 22206 15934 22258 15986
rect 26014 15934 26066 15986
rect 31726 15934 31778 15986
rect 32062 15934 32114 15986
rect 32622 15934 32674 15986
rect 36542 15934 36594 15986
rect 37214 15934 37266 15986
rect 39566 15934 39618 15986
rect 41022 15934 41074 15986
rect 45502 15934 45554 15986
rect 46286 15934 46338 15986
rect 46734 15934 46786 15986
rect 46846 15934 46898 15986
rect 47966 15934 48018 15986
rect 50318 15934 50370 15986
rect 50430 15934 50482 15986
rect 52670 15934 52722 15986
rect 52894 15934 52946 15986
rect 55246 15934 55298 15986
rect 56254 15934 56306 15986
rect 57934 15934 57986 15986
rect 6078 15822 6130 15874
rect 8318 15822 8370 15874
rect 8878 15822 8930 15874
rect 10222 15822 10274 15874
rect 11454 15822 11506 15874
rect 11678 15822 11730 15874
rect 13918 15822 13970 15874
rect 18622 15822 18674 15874
rect 18958 15822 19010 15874
rect 20078 15822 20130 15874
rect 20638 15822 20690 15874
rect 23550 15822 23602 15874
rect 26126 15822 26178 15874
rect 26350 15822 26402 15874
rect 28366 15822 28418 15874
rect 29822 15822 29874 15874
rect 31950 15822 32002 15874
rect 32510 15822 32562 15874
rect 32958 15822 33010 15874
rect 33630 15822 33682 15874
rect 33966 15822 34018 15874
rect 35758 15822 35810 15874
rect 36318 15822 36370 15874
rect 37438 15822 37490 15874
rect 38446 15822 38498 15874
rect 41358 15822 41410 15874
rect 47406 15822 47458 15874
rect 57822 15822 57874 15874
rect 15520 15654 15572 15706
rect 15624 15654 15676 15706
rect 15728 15654 15780 15706
rect 29827 15654 29879 15706
rect 29931 15654 29983 15706
rect 30035 15654 30087 15706
rect 44134 15654 44186 15706
rect 44238 15654 44290 15706
rect 44342 15654 44394 15706
rect 58441 15654 58493 15706
rect 58545 15654 58597 15706
rect 58649 15654 58701 15706
rect 5742 15486 5794 15538
rect 11454 15486 11506 15538
rect 15486 15486 15538 15538
rect 15934 15486 15986 15538
rect 16382 15486 16434 15538
rect 17614 15486 17666 15538
rect 18062 15486 18114 15538
rect 20414 15486 20466 15538
rect 21982 15486 22034 15538
rect 22206 15486 22258 15538
rect 25342 15486 25394 15538
rect 28702 15486 28754 15538
rect 28926 15486 28978 15538
rect 30718 15486 30770 15538
rect 33742 15486 33794 15538
rect 41022 15486 41074 15538
rect 42366 15486 42418 15538
rect 43150 15486 43202 15538
rect 43710 15486 43762 15538
rect 44606 15486 44658 15538
rect 47406 15486 47458 15538
rect 48078 15486 48130 15538
rect 56926 15486 56978 15538
rect 57486 15486 57538 15538
rect 5518 15374 5570 15426
rect 6526 15374 6578 15426
rect 7422 15374 7474 15426
rect 9886 15374 9938 15426
rect 10558 15374 10610 15426
rect 20750 15374 20802 15426
rect 22318 15374 22370 15426
rect 23662 15374 23714 15426
rect 26910 15374 26962 15426
rect 27246 15374 27298 15426
rect 27358 15374 27410 15426
rect 27582 15374 27634 15426
rect 28030 15374 28082 15426
rect 30270 15374 30322 15426
rect 35310 15374 35362 15426
rect 35982 15374 36034 15426
rect 36318 15374 36370 15426
rect 37438 15374 37490 15426
rect 40910 15374 40962 15426
rect 41470 15374 41522 15426
rect 41806 15374 41858 15426
rect 42926 15374 42978 15426
rect 43822 15374 43874 15426
rect 44270 15374 44322 15426
rect 48190 15374 48242 15426
rect 49198 15374 49250 15426
rect 50654 15374 50706 15426
rect 52446 15374 52498 15426
rect 55806 15374 55858 15426
rect 56030 15374 56082 15426
rect 56702 15374 56754 15426
rect 57710 15374 57762 15426
rect 1822 15262 1874 15314
rect 5966 15262 6018 15314
rect 6750 15262 6802 15314
rect 7870 15262 7922 15314
rect 10110 15262 10162 15314
rect 10782 15262 10834 15314
rect 14590 15262 14642 15314
rect 15038 15262 15090 15314
rect 21422 15262 21474 15314
rect 22766 15262 22818 15314
rect 23102 15262 23154 15314
rect 23214 15262 23266 15314
rect 23326 15262 23378 15314
rect 24110 15262 24162 15314
rect 24558 15262 24610 15314
rect 25454 15262 25506 15314
rect 26014 15262 26066 15314
rect 26462 15262 26514 15314
rect 27918 15262 27970 15314
rect 28254 15262 28306 15314
rect 28478 15262 28530 15314
rect 29374 15262 29426 15314
rect 29598 15262 29650 15314
rect 32286 15262 32338 15314
rect 33630 15262 33682 15314
rect 34414 15262 34466 15314
rect 36766 15262 36818 15314
rect 41246 15262 41298 15314
rect 42142 15262 42194 15314
rect 44942 15262 44994 15314
rect 45166 15262 45218 15314
rect 46062 15262 46114 15314
rect 46398 15262 46450 15314
rect 46622 15262 46674 15314
rect 51550 15262 51602 15314
rect 53006 15262 53058 15314
rect 54798 15262 54850 15314
rect 2494 15150 2546 15202
rect 4622 15150 4674 15202
rect 5182 15150 5234 15202
rect 7982 15150 8034 15202
rect 8990 15150 9042 15202
rect 13806 15150 13858 15202
rect 16830 15150 16882 15202
rect 11678 15094 11730 15146
rect 19070 15150 19122 15202
rect 21534 15150 21586 15202
rect 34526 15150 34578 15202
rect 39566 15150 39618 15202
rect 43262 15150 43314 15202
rect 43598 15150 43650 15202
rect 48862 15150 48914 15202
rect 50990 15150 51042 15202
rect 51662 15150 51714 15202
rect 53230 15150 53282 15202
rect 55134 15150 55186 15202
rect 55694 15150 55746 15202
rect 57038 15150 57090 15202
rect 57598 15150 57650 15202
rect 5854 15038 5906 15090
rect 14814 15038 14866 15090
rect 15598 15038 15650 15090
rect 25342 15038 25394 15090
rect 28590 15038 28642 15090
rect 33742 15038 33794 15090
rect 42478 15038 42530 15090
rect 45502 15038 45554 15090
rect 46958 15038 47010 15090
rect 48078 15038 48130 15090
rect 53790 15038 53842 15090
rect 54686 15038 54738 15090
rect 8367 14870 8419 14922
rect 8471 14870 8523 14922
rect 8575 14870 8627 14922
rect 22674 14870 22726 14922
rect 22778 14870 22830 14922
rect 22882 14870 22934 14922
rect 36981 14870 37033 14922
rect 37085 14870 37137 14922
rect 37189 14870 37241 14922
rect 51288 14870 51340 14922
rect 51392 14870 51444 14922
rect 51496 14870 51548 14922
rect 4174 14702 4226 14754
rect 4510 14702 4562 14754
rect 6862 14702 6914 14754
rect 7310 14702 7362 14754
rect 28366 14702 28418 14754
rect 55022 14702 55074 14754
rect 3166 14590 3218 14642
rect 3502 14590 3554 14642
rect 4958 14590 5010 14642
rect 6862 14590 6914 14642
rect 7310 14590 7362 14642
rect 8430 14590 8482 14642
rect 12350 14590 12402 14642
rect 14590 14590 14642 14642
rect 17054 14590 17106 14642
rect 18398 14590 18450 14642
rect 20526 14590 20578 14642
rect 24894 14590 24946 14642
rect 25342 14590 25394 14642
rect 27358 14590 27410 14642
rect 33630 14590 33682 14642
rect 35646 14590 35698 14642
rect 44942 14590 44994 14642
rect 49422 14590 49474 14642
rect 49870 14590 49922 14642
rect 50654 14590 50706 14642
rect 50990 14590 51042 14642
rect 52782 14590 52834 14642
rect 56142 14590 56194 14642
rect 1822 14478 1874 14530
rect 3390 14478 3442 14530
rect 3838 14478 3890 14530
rect 4174 14478 4226 14530
rect 4846 14478 4898 14530
rect 7646 14478 7698 14530
rect 8766 14478 8818 14530
rect 9886 14478 9938 14530
rect 10670 14478 10722 14530
rect 11230 14478 11282 14530
rect 12126 14478 12178 14530
rect 12798 14478 12850 14530
rect 15598 14478 15650 14530
rect 16606 14478 16658 14530
rect 17726 14478 17778 14530
rect 21310 14478 21362 14530
rect 21758 14478 21810 14530
rect 22206 14478 22258 14530
rect 22654 14478 22706 14530
rect 24222 14478 24274 14530
rect 24670 14478 24722 14530
rect 25454 14478 25506 14530
rect 25902 14478 25954 14530
rect 28254 14478 28306 14530
rect 29374 14478 29426 14530
rect 32958 14478 33010 14530
rect 35534 14478 35586 14530
rect 37102 14478 37154 14530
rect 38670 14478 38722 14530
rect 40014 14478 40066 14530
rect 40350 14478 40402 14530
rect 40910 14478 40962 14530
rect 41134 14478 41186 14530
rect 41806 14478 41858 14530
rect 44270 14478 44322 14530
rect 45390 14478 45442 14530
rect 46174 14478 46226 14530
rect 46846 14478 46898 14530
rect 47294 14478 47346 14530
rect 48750 14478 48802 14530
rect 51326 14478 51378 14530
rect 51774 14478 51826 14530
rect 51998 14478 52050 14530
rect 52558 14478 52610 14530
rect 52894 14478 52946 14530
rect 53118 14478 53170 14530
rect 55806 14478 55858 14530
rect 57598 14478 57650 14530
rect 2382 14366 2434 14418
rect 2718 14366 2770 14418
rect 3054 14366 3106 14418
rect 10782 14366 10834 14418
rect 11006 14366 11058 14418
rect 12574 14366 12626 14418
rect 14142 14366 14194 14418
rect 15038 14366 15090 14418
rect 15262 14366 15314 14418
rect 15934 14366 15986 14418
rect 16270 14366 16322 14418
rect 22766 14366 22818 14418
rect 23550 14366 23602 14418
rect 26798 14366 26850 14418
rect 27918 14366 27970 14418
rect 29150 14366 29202 14418
rect 29710 14366 29762 14418
rect 30270 14366 30322 14418
rect 31726 14366 31778 14418
rect 32062 14366 32114 14418
rect 34862 14366 34914 14418
rect 34974 14366 35026 14418
rect 36430 14366 36482 14418
rect 38894 14366 38946 14418
rect 39230 14366 39282 14418
rect 39342 14366 39394 14418
rect 39790 14366 39842 14418
rect 40238 14366 40290 14418
rect 40798 14366 40850 14418
rect 43934 14366 43986 14418
rect 46286 14366 46338 14418
rect 48078 14366 48130 14418
rect 48302 14366 48354 14418
rect 51102 14366 51154 14418
rect 54686 14366 54738 14418
rect 56142 14366 56194 14418
rect 2046 14254 2098 14306
rect 6078 14254 6130 14306
rect 6414 14254 6466 14306
rect 11566 14254 11618 14306
rect 13694 14254 13746 14306
rect 15150 14254 15202 14306
rect 16382 14254 16434 14306
rect 22990 14254 23042 14306
rect 23214 14254 23266 14306
rect 23438 14254 23490 14306
rect 25230 14254 25282 14306
rect 26462 14254 26514 14306
rect 28366 14254 28418 14306
rect 29262 14254 29314 14306
rect 29934 14254 29986 14306
rect 30158 14254 30210 14306
rect 32510 14254 32562 14306
rect 33070 14254 33122 14306
rect 33294 14254 33346 14306
rect 34078 14254 34130 14306
rect 34638 14254 34690 14306
rect 39566 14254 39618 14306
rect 47406 14254 47458 14306
rect 48190 14254 48242 14306
rect 48862 14254 48914 14306
rect 49086 14254 49138 14306
rect 54910 14254 54962 14306
rect 15520 14086 15572 14138
rect 15624 14086 15676 14138
rect 15728 14086 15780 14138
rect 29827 14086 29879 14138
rect 29931 14086 29983 14138
rect 30035 14086 30087 14138
rect 44134 14086 44186 14138
rect 44238 14086 44290 14138
rect 44342 14086 44394 14138
rect 58441 14086 58493 14138
rect 58545 14086 58597 14138
rect 58649 14086 58701 14138
rect 3502 13918 3554 13970
rect 7646 13918 7698 13970
rect 8766 13918 8818 13970
rect 14030 13918 14082 13970
rect 15598 13918 15650 13970
rect 16494 13918 16546 13970
rect 24782 13918 24834 13970
rect 25230 13918 25282 13970
rect 27358 13918 27410 13970
rect 28030 13918 28082 13970
rect 30718 13918 30770 13970
rect 33182 13918 33234 13970
rect 35086 13918 35138 13970
rect 35646 13918 35698 13970
rect 37326 13918 37378 13970
rect 40350 13918 40402 13970
rect 49758 13918 49810 13970
rect 53902 13918 53954 13970
rect 55918 13918 55970 13970
rect 2382 13806 2434 13858
rect 2718 13806 2770 13858
rect 2942 13806 2994 13858
rect 3726 13806 3778 13858
rect 7310 13806 7362 13858
rect 8318 13806 8370 13858
rect 8990 13806 9042 13858
rect 11790 13806 11842 13858
rect 12462 13806 12514 13858
rect 13358 13806 13410 13858
rect 13470 13806 13522 13858
rect 14366 13806 14418 13858
rect 21646 13806 21698 13858
rect 23886 13806 23938 13858
rect 29486 13806 29538 13858
rect 30942 13806 30994 13858
rect 31502 13806 31554 13858
rect 31950 13806 32002 13858
rect 33070 13806 33122 13858
rect 36430 13806 36482 13858
rect 41246 13806 41298 13858
rect 43486 13806 43538 13858
rect 46286 13806 46338 13858
rect 47294 13806 47346 13858
rect 48750 13806 48802 13858
rect 51102 13806 51154 13858
rect 53006 13806 53058 13858
rect 56030 13806 56082 13858
rect 2046 13694 2098 13746
rect 4734 13694 4786 13746
rect 6302 13694 6354 13746
rect 6750 13694 6802 13746
rect 7982 13694 8034 13746
rect 9550 13694 9602 13746
rect 10558 13694 10610 13746
rect 12126 13694 12178 13746
rect 12798 13694 12850 13746
rect 12910 13694 12962 13746
rect 13694 13694 13746 13746
rect 14702 13694 14754 13746
rect 15374 13694 15426 13746
rect 16046 13694 16098 13746
rect 16606 13694 16658 13746
rect 16830 13694 16882 13746
rect 17390 13694 17442 13746
rect 17950 13694 18002 13746
rect 18174 13694 18226 13746
rect 21422 13694 21474 13746
rect 22094 13694 22146 13746
rect 23438 13694 23490 13746
rect 25566 13694 25618 13746
rect 25902 13694 25954 13746
rect 26462 13694 26514 13746
rect 28590 13694 28642 13746
rect 30494 13694 30546 13746
rect 31614 13694 31666 13746
rect 33294 13694 33346 13746
rect 33742 13694 33794 13746
rect 36766 13694 36818 13746
rect 37326 13694 37378 13746
rect 42478 13694 42530 13746
rect 44606 13694 44658 13746
rect 47854 13694 47906 13746
rect 49086 13694 49138 13746
rect 49646 13694 49698 13746
rect 51662 13694 51714 13746
rect 52334 13694 52386 13746
rect 53566 13694 53618 13746
rect 54910 13694 54962 13746
rect 55358 13694 55410 13746
rect 56702 13694 56754 13746
rect 57262 13694 57314 13746
rect 57598 13694 57650 13746
rect 2158 13582 2210 13634
rect 3950 13582 4002 13634
rect 4174 13582 4226 13634
rect 8878 13582 8930 13634
rect 10110 13582 10162 13634
rect 10670 13582 10722 13634
rect 11566 13582 11618 13634
rect 12574 13582 12626 13634
rect 14926 13582 14978 13634
rect 18062 13582 18114 13634
rect 18622 13582 18674 13634
rect 19070 13582 19122 13634
rect 19742 13582 19794 13634
rect 20190 13582 20242 13634
rect 20638 13582 20690 13634
rect 20974 13582 21026 13634
rect 22430 13582 22482 13634
rect 23102 13582 23154 13634
rect 27022 13582 27074 13634
rect 30046 13582 30098 13634
rect 32286 13582 32338 13634
rect 32510 13582 32562 13634
rect 33966 13582 34018 13634
rect 34190 13582 34242 13634
rect 34526 13582 34578 13634
rect 39790 13582 39842 13634
rect 41134 13582 41186 13634
rect 46062 13582 46114 13634
rect 50318 13582 50370 13634
rect 53342 13582 53394 13634
rect 54686 13582 54738 13634
rect 57822 13582 57874 13634
rect 3054 13470 3106 13522
rect 3390 13470 3442 13522
rect 6526 13470 6578 13522
rect 9774 13470 9826 13522
rect 10894 13470 10946 13522
rect 15038 13470 15090 13522
rect 15710 13470 15762 13522
rect 16270 13470 16322 13522
rect 17614 13470 17666 13522
rect 19182 13470 19234 13522
rect 19966 13470 20018 13522
rect 30606 13470 30658 13522
rect 31502 13470 31554 13522
rect 40014 13470 40066 13522
rect 55918 13470 55970 13522
rect 8367 13302 8419 13354
rect 8471 13302 8523 13354
rect 8575 13302 8627 13354
rect 22674 13302 22726 13354
rect 22778 13302 22830 13354
rect 22882 13302 22934 13354
rect 36981 13302 37033 13354
rect 37085 13302 37137 13354
rect 37189 13302 37241 13354
rect 51288 13302 51340 13354
rect 51392 13302 51444 13354
rect 51496 13302 51548 13354
rect 15262 13134 15314 13186
rect 40238 13134 40290 13186
rect 41358 13134 41410 13186
rect 41694 13134 41746 13186
rect 50766 13134 50818 13186
rect 5070 13022 5122 13074
rect 6526 13022 6578 13074
rect 9550 13022 9602 13074
rect 17166 13022 17218 13074
rect 19294 13022 19346 13074
rect 22766 13022 22818 13074
rect 24894 13022 24946 13074
rect 31054 13022 31106 13074
rect 34862 13022 34914 13074
rect 39342 13022 39394 13074
rect 39902 13022 39954 13074
rect 41134 13022 41186 13074
rect 43598 13022 43650 13074
rect 45502 13022 45554 13074
rect 48974 13022 49026 13074
rect 49870 13022 49922 13074
rect 52110 13022 52162 13074
rect 55470 13022 55522 13074
rect 58046 13022 58098 13074
rect 3502 12910 3554 12962
rect 4398 12910 4450 12962
rect 4846 12910 4898 12962
rect 8094 12910 8146 12962
rect 12462 12910 12514 12962
rect 15262 12910 15314 12962
rect 15822 12910 15874 12962
rect 16382 12910 16434 12962
rect 20302 12910 20354 12962
rect 23550 12910 23602 12962
rect 24446 12910 24498 12962
rect 24670 12910 24722 12962
rect 25678 12910 25730 12962
rect 26014 12910 26066 12962
rect 26238 12910 26290 12962
rect 26462 12910 26514 12962
rect 26686 12910 26738 12962
rect 29150 12910 29202 12962
rect 29374 12910 29426 12962
rect 29934 12910 29986 12962
rect 30270 12910 30322 12962
rect 31166 12910 31218 12962
rect 32734 12910 32786 12962
rect 33630 12910 33682 12962
rect 34974 12910 35026 12962
rect 37438 12910 37490 12962
rect 37886 12910 37938 12962
rect 38558 12910 38610 12962
rect 40238 12910 40290 12962
rect 44270 12910 44322 12962
rect 45278 12910 45330 12962
rect 46286 12910 46338 12962
rect 46846 12910 46898 12962
rect 47518 12910 47570 12962
rect 49534 12910 49586 12962
rect 50206 12910 50258 12962
rect 50430 12910 50482 12962
rect 51214 12910 51266 12962
rect 51438 12910 51490 12962
rect 56590 12910 56642 12962
rect 2046 12798 2098 12850
rect 2382 12798 2434 12850
rect 3726 12798 3778 12850
rect 5742 12798 5794 12850
rect 6638 12798 6690 12850
rect 8542 12798 8594 12850
rect 8878 12798 8930 12850
rect 9214 12798 9266 12850
rect 11678 12798 11730 12850
rect 13470 12798 13522 12850
rect 13806 12798 13858 12850
rect 15598 12798 15650 12850
rect 19966 12798 20018 12850
rect 25118 12798 25170 12850
rect 25342 12798 25394 12850
rect 26910 12798 26962 12850
rect 27022 12798 27074 12850
rect 27470 12798 27522 12850
rect 30158 12798 30210 12850
rect 30942 12798 30994 12850
rect 32398 12798 32450 12850
rect 35646 12798 35698 12850
rect 45166 12798 45218 12850
rect 48638 12798 48690 12850
rect 49758 12798 49810 12850
rect 50654 12798 50706 12850
rect 57374 12798 57426 12850
rect 2718 12686 2770 12738
rect 3054 12686 3106 12738
rect 5630 12686 5682 12738
rect 13022 12686 13074 12738
rect 14254 12686 14306 12738
rect 14814 12686 14866 12738
rect 15038 12686 15090 12738
rect 20078 12686 20130 12738
rect 20862 12686 20914 12738
rect 21758 12686 21810 12738
rect 22206 12686 22258 12738
rect 22990 12686 23042 12738
rect 23886 12686 23938 12738
rect 25678 12686 25730 12738
rect 27358 12686 27410 12738
rect 28030 12686 28082 12738
rect 29262 12686 29314 12738
rect 29598 12686 29650 12738
rect 30718 12686 30770 12738
rect 33966 12686 34018 12738
rect 43934 12686 43986 12738
rect 46174 12686 46226 12738
rect 15520 12518 15572 12570
rect 15624 12518 15676 12570
rect 15728 12518 15780 12570
rect 29827 12518 29879 12570
rect 29931 12518 29983 12570
rect 30035 12518 30087 12570
rect 44134 12518 44186 12570
rect 44238 12518 44290 12570
rect 44342 12518 44394 12570
rect 58441 12518 58493 12570
rect 58545 12518 58597 12570
rect 58649 12518 58701 12570
rect 5518 12350 5570 12402
rect 7870 12350 7922 12402
rect 8094 12350 8146 12402
rect 10782 12350 10834 12402
rect 11230 12350 11282 12402
rect 17390 12350 17442 12402
rect 23998 12350 24050 12402
rect 28254 12350 28306 12402
rect 28926 12350 28978 12402
rect 32062 12350 32114 12402
rect 32286 12350 32338 12402
rect 33406 12350 33458 12402
rect 33630 12350 33682 12402
rect 37326 12350 37378 12402
rect 40014 12350 40066 12402
rect 44046 12350 44098 12402
rect 45614 12350 45666 12402
rect 47182 12350 47234 12402
rect 47854 12350 47906 12402
rect 48302 12350 48354 12402
rect 48862 12350 48914 12402
rect 55470 12350 55522 12402
rect 56702 12350 56754 12402
rect 57598 12350 57650 12402
rect 5182 12238 5234 12290
rect 7758 12238 7810 12290
rect 8318 12238 8370 12290
rect 9550 12238 9602 12290
rect 9886 12238 9938 12290
rect 10446 12238 10498 12290
rect 12350 12238 12402 12290
rect 15598 12238 15650 12290
rect 15822 12238 15874 12290
rect 18174 12238 18226 12290
rect 19854 12238 19906 12290
rect 22430 12238 22482 12290
rect 24558 12238 24610 12290
rect 27134 12238 27186 12290
rect 29934 12238 29986 12290
rect 31278 12238 31330 12290
rect 33854 12238 33906 12290
rect 36990 12238 37042 12290
rect 39342 12238 39394 12290
rect 39566 12238 39618 12290
rect 40126 12238 40178 12290
rect 44382 12238 44434 12290
rect 44718 12238 44770 12290
rect 52334 12238 52386 12290
rect 56590 12238 56642 12290
rect 56814 12238 56866 12290
rect 57262 12238 57314 12290
rect 57374 12238 57426 12290
rect 1934 12126 1986 12178
rect 6302 12126 6354 12178
rect 6638 12126 6690 12178
rect 6974 12126 7026 12178
rect 7198 12126 7250 12178
rect 7534 12126 7586 12178
rect 11566 12126 11618 12178
rect 16494 12126 16546 12178
rect 17390 12126 17442 12178
rect 17838 12126 17890 12178
rect 19070 12126 19122 12178
rect 22542 12126 22594 12178
rect 22990 12126 23042 12178
rect 23438 12126 23490 12178
rect 23550 12126 23602 12178
rect 23662 12126 23714 12178
rect 24334 12126 24386 12178
rect 25566 12126 25618 12178
rect 26238 12126 26290 12178
rect 27246 12126 27298 12178
rect 27918 12126 27970 12178
rect 28254 12126 28306 12178
rect 28478 12126 28530 12178
rect 30942 12126 30994 12178
rect 31390 12126 31442 12178
rect 31950 12126 32002 12178
rect 33182 12126 33234 12178
rect 33966 12126 34018 12178
rect 36318 12126 36370 12178
rect 36766 12126 36818 12178
rect 37662 12126 37714 12178
rect 39230 12126 39282 12178
rect 39678 12126 39730 12178
rect 40350 12126 40402 12178
rect 41134 12126 41186 12178
rect 42478 12126 42530 12178
rect 43822 12126 43874 12178
rect 45054 12126 45106 12178
rect 45390 12126 45442 12178
rect 45838 12126 45890 12178
rect 46174 12126 46226 12178
rect 46398 12126 46450 12178
rect 46622 12126 46674 12178
rect 47294 12126 47346 12178
rect 49422 12126 49474 12178
rect 50766 12126 50818 12178
rect 53566 12126 53618 12178
rect 2718 12014 2770 12066
rect 4846 11987 4898 12039
rect 6078 12014 6130 12066
rect 7086 12014 7138 12066
rect 9102 12014 9154 12066
rect 14478 12014 14530 12066
rect 16606 12014 16658 12066
rect 18846 12014 18898 12066
rect 21982 12014 22034 12066
rect 25342 12014 25394 12066
rect 26126 12014 26178 12066
rect 27582 12014 27634 12066
rect 31054 12014 31106 12066
rect 34414 12014 34466 12066
rect 34862 12014 34914 12066
rect 37886 12014 37938 12066
rect 41022 12014 41074 12066
rect 45726 12014 45778 12066
rect 46286 12014 46338 12066
rect 49758 12014 49810 12066
rect 51550 12014 51602 12066
rect 52110 12014 52162 12066
rect 55582 12014 55634 12066
rect 17614 11902 17666 11954
rect 23214 11902 23266 11954
rect 42702 11902 42754 11954
rect 47182 11902 47234 11954
rect 54910 11902 54962 11954
rect 55246 11902 55298 11954
rect 8367 11734 8419 11786
rect 8471 11734 8523 11786
rect 8575 11734 8627 11786
rect 22674 11734 22726 11786
rect 22778 11734 22830 11786
rect 22882 11734 22934 11786
rect 36981 11734 37033 11786
rect 37085 11734 37137 11786
rect 37189 11734 37241 11786
rect 51288 11734 51340 11786
rect 51392 11734 51444 11786
rect 51496 11734 51548 11786
rect 2046 11566 2098 11618
rect 3166 11566 3218 11618
rect 4174 11566 4226 11618
rect 7646 11566 7698 11618
rect 9214 11566 9266 11618
rect 10670 11566 10722 11618
rect 18622 11566 18674 11618
rect 20750 11566 20802 11618
rect 30270 11566 30322 11618
rect 35758 11566 35810 11618
rect 40910 11566 40962 11618
rect 41246 11566 41298 11618
rect 45726 11566 45778 11618
rect 51550 11566 51602 11618
rect 7982 11454 8034 11506
rect 11902 11454 11954 11506
rect 12686 11454 12738 11506
rect 15038 11454 15090 11506
rect 17166 11454 17218 11506
rect 19070 11454 19122 11506
rect 20526 11454 20578 11506
rect 27022 11454 27074 11506
rect 27806 11454 27858 11506
rect 31054 11454 31106 11506
rect 33518 11454 33570 11506
rect 35870 11454 35922 11506
rect 37102 11454 37154 11506
rect 39230 11454 39282 11506
rect 39566 11454 39618 11506
rect 39902 11454 39954 11506
rect 43486 11454 43538 11506
rect 46734 11454 46786 11506
rect 47966 11454 48018 11506
rect 50990 11454 51042 11506
rect 57934 11454 57986 11506
rect 1934 11342 1986 11394
rect 2494 11342 2546 11394
rect 3054 11342 3106 11394
rect 3390 11342 3442 11394
rect 3614 11342 3666 11394
rect 4062 11342 4114 11394
rect 4734 11342 4786 11394
rect 5854 11342 5906 11394
rect 6750 11342 6802 11394
rect 8318 11342 8370 11394
rect 9214 11342 9266 11394
rect 9438 11342 9490 11394
rect 10222 11342 10274 11394
rect 10558 11342 10610 11394
rect 10894 11342 10946 11394
rect 11454 11342 11506 11394
rect 12350 11342 12402 11394
rect 14366 11342 14418 11394
rect 17838 11342 17890 11394
rect 18174 11342 18226 11394
rect 18734 11342 18786 11394
rect 19742 11342 19794 11394
rect 19966 11342 20018 11394
rect 21310 11342 21362 11394
rect 21982 11342 22034 11394
rect 22206 11342 22258 11394
rect 22542 11342 22594 11394
rect 23326 11342 23378 11394
rect 23774 11342 23826 11394
rect 24222 11342 24274 11394
rect 24558 11342 24610 11394
rect 25230 11342 25282 11394
rect 26350 11342 26402 11394
rect 26574 11342 26626 11394
rect 26910 11342 26962 11394
rect 27134 11342 27186 11394
rect 29598 11342 29650 11394
rect 29822 11342 29874 11394
rect 31166 11342 31218 11394
rect 31502 11342 31554 11394
rect 31950 11342 32002 11394
rect 32062 11342 32114 11394
rect 32398 11342 32450 11394
rect 33294 11342 33346 11394
rect 34526 11342 34578 11394
rect 35758 11342 35810 11394
rect 36542 11342 36594 11394
rect 38558 11342 38610 11394
rect 40238 11342 40290 11394
rect 40910 11342 40962 11394
rect 45390 11342 45442 11394
rect 45726 11342 45778 11394
rect 47070 11342 47122 11394
rect 48190 11342 48242 11394
rect 49422 11342 49474 11394
rect 49758 11342 49810 11394
rect 49982 11342 50034 11394
rect 50542 11342 50594 11394
rect 54798 11342 54850 11394
rect 55246 11342 55298 11394
rect 2270 11230 2322 11282
rect 4510 11230 4562 11282
rect 5966 11230 6018 11282
rect 7086 11230 7138 11282
rect 7870 11230 7922 11282
rect 8654 11230 8706 11282
rect 9774 11230 9826 11282
rect 13470 11230 13522 11282
rect 17950 11230 18002 11282
rect 22878 11230 22930 11282
rect 25678 11230 25730 11282
rect 26014 11230 26066 11282
rect 29710 11230 29762 11282
rect 30718 11230 30770 11282
rect 31726 11230 31778 11282
rect 32734 11230 32786 11282
rect 33966 11230 34018 11282
rect 37326 11230 37378 11282
rect 45166 11230 45218 11282
rect 47630 11230 47682 11282
rect 49534 11230 49586 11282
rect 50654 11230 50706 11282
rect 51774 11230 51826 11282
rect 54574 11230 54626 11282
rect 56142 11230 56194 11282
rect 57486 11230 57538 11282
rect 2382 11118 2434 11170
rect 2830 11118 2882 11170
rect 3950 11118 4002 11170
rect 6302 11118 6354 11170
rect 8542 11118 8594 11170
rect 8990 11118 9042 11170
rect 10334 11118 10386 11170
rect 13806 11118 13858 11170
rect 20526 11118 20578 11170
rect 22766 11118 22818 11170
rect 27358 11118 27410 11170
rect 28366 11118 28418 11170
rect 30942 11118 30994 11170
rect 32510 11118 32562 11170
rect 34302 11118 34354 11170
rect 41806 11118 41858 11170
rect 42142 11118 42194 11170
rect 42590 11118 42642 11170
rect 43038 11118 43090 11170
rect 45950 11118 46002 11170
rect 48526 11118 48578 11170
rect 51662 11118 51714 11170
rect 56254 11118 56306 11170
rect 15520 10950 15572 11002
rect 15624 10950 15676 11002
rect 15728 10950 15780 11002
rect 29827 10950 29879 11002
rect 29931 10950 29983 11002
rect 30035 10950 30087 11002
rect 44134 10950 44186 11002
rect 44238 10950 44290 11002
rect 44342 10950 44394 11002
rect 58441 10950 58493 11002
rect 58545 10950 58597 11002
rect 58649 10950 58701 11002
rect 2046 10782 2098 10834
rect 5742 10782 5794 10834
rect 16382 10782 16434 10834
rect 25342 10782 25394 10834
rect 25566 10782 25618 10834
rect 26126 10782 26178 10834
rect 26910 10782 26962 10834
rect 32174 10782 32226 10834
rect 33070 10782 33122 10834
rect 35870 10782 35922 10834
rect 36430 10782 36482 10834
rect 36878 10782 36930 10834
rect 42926 10782 42978 10834
rect 43262 10782 43314 10834
rect 45166 10782 45218 10834
rect 53902 10782 53954 10834
rect 1710 10670 1762 10722
rect 3278 10670 3330 10722
rect 7870 10670 7922 10722
rect 12686 10670 12738 10722
rect 13582 10670 13634 10722
rect 14702 10670 14754 10722
rect 20078 10670 20130 10722
rect 22766 10670 22818 10722
rect 27358 10670 27410 10722
rect 31054 10670 31106 10722
rect 35310 10670 35362 10722
rect 36318 10670 36370 10722
rect 37102 10670 37154 10722
rect 37214 10670 37266 10722
rect 39566 10670 39618 10722
rect 42702 10670 42754 10722
rect 46398 10670 46450 10722
rect 48750 10670 48802 10722
rect 55358 10670 55410 10722
rect 2494 10558 2546 10610
rect 6638 10558 6690 10610
rect 7422 10558 7474 10610
rect 8318 10558 8370 10610
rect 8990 10558 9042 10610
rect 9886 10558 9938 10610
rect 10446 10558 10498 10610
rect 10670 10558 10722 10610
rect 12574 10558 12626 10610
rect 14254 10558 14306 10610
rect 14926 10558 14978 10610
rect 19294 10558 19346 10610
rect 19742 10558 19794 10610
rect 21646 10558 21698 10610
rect 22990 10558 23042 10610
rect 23774 10558 23826 10610
rect 24334 10558 24386 10610
rect 25230 10558 25282 10610
rect 26126 10558 26178 10610
rect 27470 10558 27522 10610
rect 27806 10558 27858 10610
rect 28814 10558 28866 10610
rect 29710 10558 29762 10610
rect 30942 10558 30994 10610
rect 31726 10558 31778 10610
rect 33406 10558 33458 10610
rect 34302 10558 34354 10610
rect 34862 10558 34914 10610
rect 35086 10558 35138 10610
rect 35422 10558 35474 10610
rect 35758 10558 35810 10610
rect 36654 10558 36706 10610
rect 38894 10558 38946 10610
rect 39230 10558 39282 10610
rect 40126 10558 40178 10610
rect 40910 10558 40962 10610
rect 41806 10558 41858 10610
rect 42254 10558 42306 10610
rect 43150 10558 43202 10610
rect 44270 10558 44322 10610
rect 44606 10558 44658 10610
rect 44718 10558 44770 10610
rect 45054 10558 45106 10610
rect 45950 10558 46002 10610
rect 46174 10558 46226 10610
rect 47070 10558 47122 10610
rect 49310 10558 49362 10610
rect 51326 10558 51378 10610
rect 54462 10558 54514 10610
rect 57150 10558 57202 10610
rect 5406 10446 5458 10498
rect 5854 10446 5906 10498
rect 6414 10446 6466 10498
rect 10558 10446 10610 10498
rect 11006 10446 11058 10498
rect 15262 10446 15314 10498
rect 15934 10446 15986 10498
rect 16830 10446 16882 10498
rect 17838 10446 17890 10498
rect 18174 10446 18226 10498
rect 19182 10446 19234 10498
rect 19630 10446 19682 10498
rect 22206 10446 22258 10498
rect 23438 10446 23490 10498
rect 28254 10446 28306 10498
rect 29822 10446 29874 10498
rect 30830 10446 30882 10498
rect 33966 10446 34018 10498
rect 39342 10446 39394 10498
rect 41134 10446 41186 10498
rect 41470 10446 41522 10498
rect 43262 10446 43314 10498
rect 46286 10446 46338 10498
rect 46846 10446 46898 10498
rect 49534 10446 49586 10498
rect 51550 10446 51602 10498
rect 51998 10446 52050 10498
rect 55918 10446 55970 10498
rect 56814 10446 56866 10498
rect 57598 10446 57650 10498
rect 6750 10334 6802 10386
rect 10110 10334 10162 10386
rect 18398 10334 18450 10386
rect 18734 10334 18786 10386
rect 20862 10334 20914 10386
rect 28702 10334 28754 10386
rect 31726 10334 31778 10386
rect 32062 10334 32114 10386
rect 33630 10334 33682 10386
rect 33966 10334 34018 10386
rect 35870 10334 35922 10386
rect 45166 10334 45218 10386
rect 46734 10334 46786 10386
rect 8367 10166 8419 10218
rect 8471 10166 8523 10218
rect 8575 10166 8627 10218
rect 22674 10166 22726 10218
rect 22778 10166 22830 10218
rect 22882 10166 22934 10218
rect 36981 10166 37033 10218
rect 37085 10166 37137 10218
rect 37189 10166 37241 10218
rect 51288 10166 51340 10218
rect 51392 10166 51444 10218
rect 51496 10166 51548 10218
rect 11006 9998 11058 10050
rect 29598 9998 29650 10050
rect 35646 9998 35698 10050
rect 40014 9998 40066 10050
rect 48750 9998 48802 10050
rect 50654 9998 50706 10050
rect 2494 9886 2546 9938
rect 4622 9886 4674 9938
rect 5182 9886 5234 9938
rect 5854 9886 5906 9938
rect 12462 9886 12514 9938
rect 12798 9886 12850 9938
rect 17502 9886 17554 9938
rect 19630 9886 19682 9938
rect 25230 9886 25282 9938
rect 26014 9886 26066 9938
rect 27246 9886 27298 9938
rect 27918 9886 27970 9938
rect 29822 9886 29874 9938
rect 32622 9886 32674 9938
rect 34190 9886 34242 9938
rect 34862 9886 34914 9938
rect 36206 9886 36258 9938
rect 39230 9886 39282 9938
rect 39678 9886 39730 9938
rect 40126 9886 40178 9938
rect 45166 9886 45218 9938
rect 47070 9886 47122 9938
rect 54910 9886 54962 9938
rect 56590 9886 56642 9938
rect 1822 9774 1874 9826
rect 6302 9774 6354 9826
rect 7982 9774 8034 9826
rect 9662 9774 9714 9826
rect 10670 9774 10722 9826
rect 11454 9774 11506 9826
rect 14478 9774 14530 9826
rect 15150 9774 15202 9826
rect 16382 9774 16434 9826
rect 16830 9774 16882 9826
rect 20638 9774 20690 9826
rect 21982 9774 22034 9826
rect 23662 9774 23714 9826
rect 25790 9774 25842 9826
rect 26126 9774 26178 9826
rect 27022 9774 27074 9826
rect 28254 9774 28306 9826
rect 29710 9774 29762 9826
rect 30718 9774 30770 9826
rect 30942 9774 30994 9826
rect 32062 9774 32114 9826
rect 33630 9774 33682 9826
rect 34078 9774 34130 9826
rect 34302 9774 34354 9826
rect 35086 9774 35138 9826
rect 39006 9774 39058 9826
rect 40350 9774 40402 9826
rect 41022 9774 41074 9826
rect 42814 9774 42866 9826
rect 44046 9774 44098 9826
rect 44830 9774 44882 9826
rect 45054 9774 45106 9826
rect 45950 9774 46002 9826
rect 46622 9774 46674 9826
rect 47406 9774 47458 9826
rect 48526 9774 48578 9826
rect 48974 9774 49026 9826
rect 49310 9774 49362 9826
rect 49534 9774 49586 9826
rect 50542 9774 50594 9826
rect 50990 9774 51042 9826
rect 52558 9774 52610 9826
rect 53118 9774 53170 9826
rect 55134 9774 55186 9826
rect 55806 9774 55858 9826
rect 57150 9774 57202 9826
rect 6750 9662 6802 9714
rect 9438 9662 9490 9714
rect 11230 9662 11282 9714
rect 12910 9662 12962 9714
rect 13918 9662 13970 9714
rect 15822 9662 15874 9714
rect 20750 9662 20802 9714
rect 21534 9662 21586 9714
rect 22542 9662 22594 9714
rect 23550 9662 23602 9714
rect 26686 9662 26738 9714
rect 27134 9662 27186 9714
rect 31390 9662 31442 9714
rect 31726 9662 31778 9714
rect 33070 9662 33122 9714
rect 33182 9662 33234 9714
rect 40686 9662 40738 9714
rect 41694 9662 41746 9714
rect 42030 9662 42082 9714
rect 42142 9662 42194 9714
rect 43486 9662 43538 9714
rect 43710 9662 43762 9714
rect 45278 9662 45330 9714
rect 45614 9662 45666 9714
rect 45726 9662 45778 9714
rect 46510 9662 46562 9714
rect 46958 9662 47010 9714
rect 53006 9662 53058 9714
rect 57710 9662 57762 9714
rect 8766 9550 8818 9602
rect 10670 9550 10722 9602
rect 12014 9550 12066 9602
rect 20190 9550 20242 9602
rect 21646 9550 21698 9602
rect 32846 9550 32898 9602
rect 38334 9550 38386 9602
rect 40798 9550 40850 9602
rect 41470 9550 41522 9602
rect 41582 9550 41634 9602
rect 42366 9550 42418 9602
rect 42478 9550 42530 9602
rect 42702 9550 42754 9602
rect 43150 9550 43202 9602
rect 43934 9550 43986 9602
rect 48078 9550 48130 9602
rect 52894 9550 52946 9602
rect 55470 9550 55522 9602
rect 15520 9382 15572 9434
rect 15624 9382 15676 9434
rect 15728 9382 15780 9434
rect 29827 9382 29879 9434
rect 29931 9382 29983 9434
rect 30035 9382 30087 9434
rect 44134 9382 44186 9434
rect 44238 9382 44290 9434
rect 44342 9382 44394 9434
rect 58441 9382 58493 9434
rect 58545 9382 58597 9434
rect 58649 9382 58701 9434
rect 1822 9214 1874 9266
rect 2158 9214 2210 9266
rect 3054 9214 3106 9266
rect 3726 9214 3778 9266
rect 4062 9214 4114 9266
rect 4846 9214 4898 9266
rect 6750 9214 6802 9266
rect 20414 9214 20466 9266
rect 22318 9214 22370 9266
rect 29374 9214 29426 9266
rect 31166 9214 31218 9266
rect 31278 9214 31330 9266
rect 39342 9214 39394 9266
rect 39678 9214 39730 9266
rect 40910 9214 40962 9266
rect 43934 9214 43986 9266
rect 44494 9214 44546 9266
rect 44942 9214 44994 9266
rect 45278 9214 45330 9266
rect 46286 9214 46338 9266
rect 47406 9214 47458 9266
rect 53902 9214 53954 9266
rect 57486 9214 57538 9266
rect 2718 9102 2770 9154
rect 5854 9102 5906 9154
rect 7534 9102 7586 9154
rect 9886 9102 9938 9154
rect 11006 9102 11058 9154
rect 15038 9102 15090 9154
rect 16494 9102 16546 9154
rect 16830 9102 16882 9154
rect 23102 9102 23154 9154
rect 24558 9102 24610 9154
rect 27806 9102 27858 9154
rect 30494 9102 30546 9154
rect 32174 9102 32226 9154
rect 37326 9102 37378 9154
rect 40014 9102 40066 9154
rect 41246 9102 41298 9154
rect 41806 9102 41858 9154
rect 46510 9102 46562 9154
rect 50990 9102 51042 9154
rect 52334 9102 52386 9154
rect 53790 9102 53842 9154
rect 54014 9102 54066 9154
rect 54798 9102 54850 9154
rect 54910 9102 54962 9154
rect 56702 9102 56754 9154
rect 5406 8990 5458 9042
rect 7646 8990 7698 9042
rect 9550 8990 9602 9042
rect 10222 8990 10274 9042
rect 13582 8990 13634 9042
rect 13918 8990 13970 9042
rect 17502 8990 17554 9042
rect 18174 8990 18226 9042
rect 22430 8990 22482 9042
rect 22990 8990 23042 9042
rect 24110 8990 24162 9042
rect 25678 8990 25730 9042
rect 25902 8990 25954 9042
rect 26910 8990 26962 9042
rect 27694 8990 27746 9042
rect 28030 8990 28082 9042
rect 28590 8990 28642 9042
rect 29934 8990 29986 9042
rect 31054 8990 31106 9042
rect 31726 8990 31778 9042
rect 32510 8990 32562 9042
rect 33182 8990 33234 9042
rect 33742 8990 33794 9042
rect 34526 8990 34578 9042
rect 36318 8990 36370 9042
rect 36766 8990 36818 9042
rect 37214 8990 37266 9042
rect 38110 8990 38162 9042
rect 42030 8990 42082 9042
rect 42590 8990 42642 9042
rect 43038 8990 43090 9042
rect 44046 8990 44098 9042
rect 45502 8990 45554 9042
rect 45950 8990 46002 9042
rect 47630 8990 47682 9042
rect 48862 8990 48914 9042
rect 49086 8990 49138 9042
rect 49758 8990 49810 9042
rect 51662 8990 51714 9042
rect 51886 8990 51938 9042
rect 53118 8990 53170 9042
rect 55358 8990 55410 9042
rect 56590 8990 56642 9042
rect 57486 8990 57538 9042
rect 9662 8878 9714 8930
rect 13134 8878 13186 8930
rect 15486 8878 15538 8930
rect 15598 8878 15650 8930
rect 16270 8878 16322 8930
rect 20862 8878 20914 8930
rect 23438 8878 23490 8930
rect 24334 8878 24386 8930
rect 27918 8878 27970 8930
rect 29038 8878 29090 8930
rect 30606 8878 30658 8930
rect 34862 8878 34914 8930
rect 35534 8878 35586 8930
rect 35758 8878 35810 8930
rect 38334 8878 38386 8930
rect 38894 8878 38946 8930
rect 45390 8878 45442 8930
rect 46286 8878 46338 8930
rect 47518 8878 47570 8930
rect 52894 8878 52946 8930
rect 8206 8766 8258 8818
rect 8542 8766 8594 8818
rect 21086 8766 21138 8818
rect 21310 8766 21362 8818
rect 21758 8766 21810 8818
rect 26798 8766 26850 8818
rect 27358 8766 27410 8818
rect 30270 8766 30322 8818
rect 35982 8766 36034 8818
rect 38670 8766 38722 8818
rect 43374 8766 43426 8818
rect 43934 8766 43986 8818
rect 49982 8766 50034 8818
rect 54910 8766 54962 8818
rect 55582 8766 55634 8818
rect 55918 8766 55970 8818
rect 8367 8598 8419 8650
rect 8471 8598 8523 8650
rect 8575 8598 8627 8650
rect 22674 8598 22726 8650
rect 22778 8598 22830 8650
rect 22882 8598 22934 8650
rect 36981 8598 37033 8650
rect 37085 8598 37137 8650
rect 37189 8598 37241 8650
rect 51288 8598 51340 8650
rect 51392 8598 51444 8650
rect 51496 8598 51548 8650
rect 22430 8430 22482 8482
rect 33518 8430 33570 8482
rect 35982 8430 36034 8482
rect 41246 8430 41298 8482
rect 54350 8430 54402 8482
rect 55918 8430 55970 8482
rect 57150 8430 57202 8482
rect 4622 8318 4674 8370
rect 5182 8318 5234 8370
rect 7758 8318 7810 8370
rect 9774 8318 9826 8370
rect 11902 8318 11954 8370
rect 15038 8318 15090 8370
rect 18510 8318 18562 8370
rect 20078 8318 20130 8370
rect 25566 8318 25618 8370
rect 29598 8318 29650 8370
rect 30606 8318 30658 8370
rect 34750 8318 34802 8370
rect 39902 8318 39954 8370
rect 45390 8318 45442 8370
rect 46510 8318 46562 8370
rect 47294 8318 47346 8370
rect 47406 8318 47458 8370
rect 49310 8318 49362 8370
rect 50206 8318 50258 8370
rect 53230 8318 53282 8370
rect 54686 8318 54738 8370
rect 55134 8318 55186 8370
rect 56254 8318 56306 8370
rect 57374 8318 57426 8370
rect 1822 8206 1874 8258
rect 6190 8206 6242 8258
rect 8990 8206 9042 8258
rect 12462 8206 12514 8258
rect 13022 8206 13074 8258
rect 13582 8206 13634 8258
rect 16494 8206 16546 8258
rect 17166 8206 17218 8258
rect 17726 8206 17778 8258
rect 18622 8206 18674 8258
rect 20638 8206 20690 8258
rect 22206 8206 22258 8258
rect 22766 8206 22818 8258
rect 23102 8206 23154 8258
rect 23998 8206 24050 8258
rect 24334 8206 24386 8258
rect 25902 8206 25954 8258
rect 26014 8206 26066 8258
rect 26238 8206 26290 8258
rect 26350 8206 26402 8258
rect 27582 8206 27634 8258
rect 27918 8206 27970 8258
rect 30046 8206 30098 8258
rect 31950 8206 32002 8258
rect 32734 8206 32786 8258
rect 33182 8206 33234 8258
rect 36094 8206 36146 8258
rect 37774 8206 37826 8258
rect 38670 8206 38722 8258
rect 42590 8206 42642 8258
rect 45726 8206 45778 8258
rect 46062 8206 46114 8258
rect 46398 8206 46450 8258
rect 47070 8206 47122 8258
rect 48190 8206 48242 8258
rect 49534 8206 49586 8258
rect 49982 8206 50034 8258
rect 54910 8206 54962 8258
rect 55246 8206 55298 8258
rect 55470 8206 55522 8258
rect 56478 8206 56530 8258
rect 57150 8206 57202 8258
rect 58046 8206 58098 8258
rect 2494 8094 2546 8146
rect 7198 8094 7250 8146
rect 12686 8094 12738 8146
rect 13806 8094 13858 8146
rect 14254 8094 14306 8146
rect 14366 8094 14418 8146
rect 14702 8094 14754 8146
rect 15262 8094 15314 8146
rect 15598 8094 15650 8146
rect 15934 8094 15986 8146
rect 17838 8094 17890 8146
rect 19182 8094 19234 8146
rect 27022 8094 27074 8146
rect 28478 8094 28530 8146
rect 31278 8094 31330 8146
rect 32174 8094 32226 8146
rect 33742 8094 33794 8146
rect 35198 8094 35250 8146
rect 35982 8094 36034 8146
rect 37438 8094 37490 8146
rect 40238 8094 40290 8146
rect 42142 8094 42194 8146
rect 43710 8094 43762 8146
rect 43934 8094 43986 8146
rect 44830 8094 44882 8146
rect 47518 8094 47570 8146
rect 48302 8094 48354 8146
rect 48750 8094 48802 8146
rect 54574 8094 54626 8146
rect 5742 7982 5794 8034
rect 8766 7982 8818 8034
rect 12798 7982 12850 8034
rect 14030 7982 14082 8034
rect 14926 7982 14978 8034
rect 15486 7982 15538 8034
rect 21422 7982 21474 8034
rect 21758 7982 21810 8034
rect 28366 7982 28418 8034
rect 29150 7982 29202 8034
rect 30942 7982 30994 8034
rect 35534 7982 35586 8034
rect 44942 7982 44994 8034
rect 46622 7982 46674 8034
rect 53342 7982 53394 8034
rect 53454 7982 53506 8034
rect 54126 7982 54178 8034
rect 15520 7814 15572 7866
rect 15624 7814 15676 7866
rect 15728 7814 15780 7866
rect 29827 7814 29879 7866
rect 29931 7814 29983 7866
rect 30035 7814 30087 7866
rect 44134 7814 44186 7866
rect 44238 7814 44290 7866
rect 44342 7814 44394 7866
rect 58441 7814 58493 7866
rect 58545 7814 58597 7866
rect 58649 7814 58701 7866
rect 2270 7646 2322 7698
rect 2494 7646 2546 7698
rect 3838 7646 3890 7698
rect 4510 7646 4562 7698
rect 4958 7646 5010 7698
rect 6638 7646 6690 7698
rect 15038 7646 15090 7698
rect 17502 7646 17554 7698
rect 19294 7646 19346 7698
rect 25230 7646 25282 7698
rect 30830 7646 30882 7698
rect 34526 7646 34578 7698
rect 35422 7646 35474 7698
rect 36094 7646 36146 7698
rect 36318 7646 36370 7698
rect 37326 7646 37378 7698
rect 37774 7646 37826 7698
rect 38670 7646 38722 7698
rect 40014 7646 40066 7698
rect 41134 7646 41186 7698
rect 44830 7646 44882 7698
rect 47630 7646 47682 7698
rect 47854 7646 47906 7698
rect 55022 7646 55074 7698
rect 2830 7534 2882 7586
rect 3166 7534 3218 7586
rect 10334 7534 10386 7586
rect 14030 7534 14082 7586
rect 18958 7534 19010 7586
rect 27806 7534 27858 7586
rect 28814 7534 28866 7586
rect 30942 7534 30994 7586
rect 31278 7534 31330 7586
rect 34190 7534 34242 7586
rect 36430 7534 36482 7586
rect 36878 7534 36930 7586
rect 38782 7534 38834 7586
rect 39342 7534 39394 7586
rect 41582 7534 41634 7586
rect 43262 7534 43314 7586
rect 46958 7534 47010 7586
rect 50318 7534 50370 7586
rect 54126 7534 54178 7586
rect 3502 7422 3554 7474
rect 5406 7422 5458 7474
rect 5630 7422 5682 7474
rect 5966 7422 6018 7474
rect 6190 7422 6242 7474
rect 6862 7422 6914 7474
rect 7198 7422 7250 7474
rect 8206 7422 8258 7474
rect 9662 7422 9714 7474
rect 13582 7422 13634 7474
rect 16382 7422 16434 7474
rect 18062 7422 18114 7474
rect 18846 7422 18898 7474
rect 20414 7422 20466 7474
rect 22318 7422 22370 7474
rect 22990 7422 23042 7474
rect 23550 7422 23602 7474
rect 26798 7422 26850 7474
rect 27022 7422 27074 7474
rect 28366 7422 28418 7474
rect 28702 7422 28754 7474
rect 29822 7422 29874 7474
rect 30382 7422 30434 7474
rect 33518 7422 33570 7474
rect 33742 7422 33794 7474
rect 35310 7422 35362 7474
rect 35534 7422 35586 7474
rect 35982 7422 36034 7474
rect 39118 7422 39170 7474
rect 40126 7422 40178 7474
rect 40910 7422 40962 7474
rect 41470 7422 41522 7474
rect 42366 7422 42418 7474
rect 43486 7422 43538 7474
rect 43822 7422 43874 7474
rect 44606 7422 44658 7474
rect 44942 7422 44994 7474
rect 46398 7422 46450 7474
rect 47518 7422 47570 7474
rect 48078 7422 48130 7474
rect 48190 7422 48242 7474
rect 49534 7422 49586 7474
rect 50542 7422 50594 7474
rect 51550 7422 51602 7474
rect 53006 7422 53058 7474
rect 54350 7422 54402 7474
rect 54910 7422 54962 7474
rect 56926 7422 56978 7474
rect 57262 7422 57314 7474
rect 3950 7310 4002 7362
rect 5518 7310 5570 7362
rect 6750 7310 6802 7362
rect 7310 7310 7362 7362
rect 7758 7310 7810 7362
rect 9102 7310 9154 7362
rect 12462 7310 12514 7362
rect 13246 7310 13298 7362
rect 14478 7310 14530 7362
rect 15934 7310 15986 7362
rect 16718 7310 16770 7362
rect 18398 7310 18450 7362
rect 19854 7310 19906 7362
rect 20862 7310 20914 7362
rect 25790 7310 25842 7362
rect 29150 7310 29202 7362
rect 32286 7310 32338 7362
rect 33854 7310 33906 7362
rect 34974 7310 35026 7362
rect 42814 7310 42866 7362
rect 44382 7310 44434 7362
rect 46174 7310 46226 7362
rect 49198 7310 49250 7362
rect 51438 7310 51490 7362
rect 56814 7310 56866 7362
rect 14702 7198 14754 7250
rect 15374 7198 15426 7250
rect 15710 7198 15762 7250
rect 23214 7198 23266 7250
rect 30830 7198 30882 7250
rect 38670 7198 38722 7250
rect 49534 7198 49586 7250
rect 50878 7198 50930 7250
rect 53118 7198 53170 7250
rect 8367 7030 8419 7082
rect 8471 7030 8523 7082
rect 8575 7030 8627 7082
rect 22674 7030 22726 7082
rect 22778 7030 22830 7082
rect 22882 7030 22934 7082
rect 36981 7030 37033 7082
rect 37085 7030 37137 7082
rect 37189 7030 37241 7082
rect 51288 7030 51340 7082
rect 51392 7030 51444 7082
rect 51496 7030 51548 7082
rect 19966 6862 20018 6914
rect 20190 6862 20242 6914
rect 20638 6862 20690 6914
rect 28254 6862 28306 6914
rect 35422 6862 35474 6914
rect 36318 6862 36370 6914
rect 39790 6862 39842 6914
rect 49310 6862 49362 6914
rect 50878 6862 50930 6914
rect 51886 6862 51938 6914
rect 58046 6862 58098 6914
rect 2606 6750 2658 6802
rect 4734 6750 4786 6802
rect 6414 6750 6466 6802
rect 14366 6750 14418 6802
rect 23102 6750 23154 6802
rect 28590 6750 28642 6802
rect 35086 6750 35138 6802
rect 35982 6750 36034 6802
rect 43038 6750 43090 6802
rect 45950 6750 46002 6802
rect 49534 6750 49586 6802
rect 50094 6750 50146 6802
rect 50430 6750 50482 6802
rect 55806 6750 55858 6802
rect 57262 6750 57314 6802
rect 1934 6638 1986 6690
rect 5742 6638 5794 6690
rect 6302 6638 6354 6690
rect 7534 6638 7586 6690
rect 7870 6638 7922 6690
rect 8542 6638 8594 6690
rect 12126 6638 12178 6690
rect 12238 6638 12290 6690
rect 12574 6638 12626 6690
rect 13470 6638 13522 6690
rect 14030 6638 14082 6690
rect 15486 6638 15538 6690
rect 16270 6638 16322 6690
rect 16830 6638 16882 6690
rect 18622 6638 18674 6690
rect 19070 6638 19122 6690
rect 20526 6638 20578 6690
rect 22766 6638 22818 6690
rect 26126 6638 26178 6690
rect 26686 6638 26738 6690
rect 28030 6638 28082 6690
rect 31054 6638 31106 6690
rect 31278 6638 31330 6690
rect 32622 6638 32674 6690
rect 33406 6638 33458 6690
rect 33966 6638 34018 6690
rect 34302 6638 34354 6690
rect 34862 6638 34914 6690
rect 35758 6638 35810 6690
rect 38558 6638 38610 6690
rect 38894 6638 38946 6690
rect 39902 6638 39954 6690
rect 42366 6638 42418 6690
rect 43598 6638 43650 6690
rect 44046 6638 44098 6690
rect 44158 6638 44210 6690
rect 45838 6638 45890 6690
rect 46958 6638 47010 6690
rect 47742 6638 47794 6690
rect 48862 6638 48914 6690
rect 51774 6638 51826 6690
rect 53006 6638 53058 6690
rect 53566 6638 53618 6690
rect 54014 6638 54066 6690
rect 54350 6638 54402 6690
rect 57150 6638 57202 6690
rect 58158 6638 58210 6690
rect 6526 6526 6578 6578
rect 17502 6526 17554 6578
rect 17838 6526 17890 6578
rect 20750 6526 20802 6578
rect 21870 6526 21922 6578
rect 25230 6526 25282 6578
rect 27358 6526 27410 6578
rect 28478 6526 28530 6578
rect 29150 6526 29202 6578
rect 30830 6526 30882 6578
rect 31166 6526 31218 6578
rect 31614 6526 31666 6578
rect 31950 6526 32002 6578
rect 32286 6526 32338 6578
rect 32398 6526 32450 6578
rect 32846 6526 32898 6578
rect 33294 6526 33346 6578
rect 37550 6526 37602 6578
rect 41694 6526 41746 6578
rect 43710 6526 43762 6578
rect 45726 6526 45778 6578
rect 47854 6526 47906 6578
rect 50318 6526 50370 6578
rect 50878 6526 50930 6578
rect 51326 6526 51378 6578
rect 53678 6526 53730 6578
rect 57598 6526 57650 6578
rect 10782 6414 10834 6466
rect 11342 6414 11394 6466
rect 11902 6414 11954 6466
rect 12910 6414 12962 6466
rect 15150 6414 15202 6466
rect 23326 6414 23378 6466
rect 24334 6414 24386 6466
rect 29710 6414 29762 6466
rect 34078 6414 34130 6466
rect 37662 6414 37714 6466
rect 40798 6414 40850 6466
rect 42142 6414 42194 6466
rect 48078 6414 48130 6466
rect 54126 6414 54178 6466
rect 55694 6414 55746 6466
rect 55918 6414 55970 6466
rect 56142 6414 56194 6466
rect 58046 6414 58098 6466
rect 15520 6246 15572 6298
rect 15624 6246 15676 6298
rect 15728 6246 15780 6298
rect 29827 6246 29879 6298
rect 29931 6246 29983 6298
rect 30035 6246 30087 6298
rect 44134 6246 44186 6298
rect 44238 6246 44290 6298
rect 44342 6246 44394 6298
rect 58441 6246 58493 6298
rect 58545 6246 58597 6298
rect 58649 6246 58701 6298
rect 1934 6078 1986 6130
rect 2494 6078 2546 6130
rect 4734 6078 4786 6130
rect 5294 6078 5346 6130
rect 8206 6078 8258 6130
rect 8990 6078 9042 6130
rect 9774 6078 9826 6130
rect 10222 6078 10274 6130
rect 13918 6078 13970 6130
rect 14478 6078 14530 6130
rect 14814 6078 14866 6130
rect 22766 6078 22818 6130
rect 24670 6078 24722 6130
rect 27246 6078 27298 6130
rect 32398 6078 32450 6130
rect 33182 6078 33234 6130
rect 34750 6078 34802 6130
rect 38110 6078 38162 6130
rect 38222 6078 38274 6130
rect 39006 6078 39058 6130
rect 53566 6078 53618 6130
rect 54126 6078 54178 6130
rect 57822 6078 57874 6130
rect 3278 5966 3330 6018
rect 4622 5966 4674 6018
rect 6638 5966 6690 6018
rect 8654 5966 8706 6018
rect 10446 5966 10498 6018
rect 10782 5966 10834 6018
rect 11118 5966 11170 6018
rect 11230 5966 11282 6018
rect 11902 5966 11954 6018
rect 12238 5966 12290 6018
rect 12350 5966 12402 6018
rect 13022 5966 13074 6018
rect 19854 5966 19906 6018
rect 21646 5966 21698 6018
rect 23662 5966 23714 6018
rect 25230 5966 25282 6018
rect 27806 5966 27858 6018
rect 28814 5966 28866 6018
rect 31838 5966 31890 6018
rect 33966 5966 34018 6018
rect 34190 5966 34242 6018
rect 37326 5966 37378 6018
rect 38670 5966 38722 6018
rect 41246 5966 41298 6018
rect 43598 5966 43650 6018
rect 50990 5966 51042 6018
rect 51886 5966 51938 6018
rect 54014 5966 54066 6018
rect 54686 5966 54738 6018
rect 54798 5966 54850 6018
rect 55806 5966 55858 6018
rect 58046 5966 58098 6018
rect 3614 5854 3666 5906
rect 5518 5854 5570 5906
rect 5966 5854 6018 5906
rect 6302 5854 6354 5906
rect 7758 5854 7810 5906
rect 12574 5854 12626 5906
rect 12798 5854 12850 5906
rect 13358 5854 13410 5906
rect 13806 5854 13858 5906
rect 14030 5854 14082 5906
rect 15822 5854 15874 5906
rect 16158 5854 16210 5906
rect 17838 5854 17890 5906
rect 18958 5854 19010 5906
rect 22094 5854 22146 5906
rect 22542 5854 22594 5906
rect 25342 5854 25394 5906
rect 26014 5854 26066 5906
rect 26574 5854 26626 5906
rect 27470 5854 27522 5906
rect 28926 5854 28978 5906
rect 29710 5854 29762 5906
rect 31390 5854 31442 5906
rect 32286 5854 32338 5906
rect 32958 5854 33010 5906
rect 33294 5854 33346 5906
rect 33854 5854 33906 5906
rect 34302 5854 34354 5906
rect 35534 5854 35586 5906
rect 36542 5854 36594 5906
rect 39790 5854 39842 5906
rect 40238 5854 40290 5906
rect 42478 5854 42530 5906
rect 44270 5854 44322 5906
rect 44718 5854 44770 5906
rect 46286 5854 46338 5906
rect 46510 5854 46562 5906
rect 47182 5854 47234 5906
rect 47630 5854 47682 5906
rect 48862 5854 48914 5906
rect 49310 5854 49362 5906
rect 50430 5854 50482 5906
rect 53230 5854 53282 5906
rect 54462 5854 54514 5906
rect 56030 5854 56082 5906
rect 56590 5854 56642 5906
rect 57038 5854 57090 5906
rect 57486 5854 57538 5906
rect 58158 5854 58210 5906
rect 13134 5742 13186 5794
rect 16718 5742 16770 5794
rect 18286 5742 18338 5794
rect 31054 5742 31106 5794
rect 35086 5742 35138 5794
rect 41022 5742 41074 5794
rect 45838 5742 45890 5794
rect 47854 5742 47906 5794
rect 49758 5742 49810 5794
rect 50094 5742 50146 5794
rect 50206 5742 50258 5794
rect 50878 5742 50930 5794
rect 51662 5742 51714 5794
rect 55694 5742 55746 5794
rect 5966 5630 6018 5682
rect 11230 5630 11282 5682
rect 26350 5630 26402 5682
rect 38334 5630 38386 5682
rect 48190 5630 48242 5682
rect 50766 5630 50818 5682
rect 54126 5630 54178 5682
rect 8367 5462 8419 5514
rect 8471 5462 8523 5514
rect 8575 5462 8627 5514
rect 22674 5462 22726 5514
rect 22778 5462 22830 5514
rect 22882 5462 22934 5514
rect 36981 5462 37033 5514
rect 37085 5462 37137 5514
rect 37189 5462 37241 5514
rect 51288 5462 51340 5514
rect 51392 5462 51444 5514
rect 51496 5462 51548 5514
rect 5070 5294 5122 5346
rect 9102 5294 9154 5346
rect 12910 5294 12962 5346
rect 26238 5294 26290 5346
rect 26798 5294 26850 5346
rect 29262 5294 29314 5346
rect 29598 5294 29650 5346
rect 30606 5294 30658 5346
rect 32622 5294 32674 5346
rect 41134 5294 41186 5346
rect 47966 5294 48018 5346
rect 48974 5294 49026 5346
rect 49422 5294 49474 5346
rect 49758 5294 49810 5346
rect 51102 5294 51154 5346
rect 55246 5294 55298 5346
rect 3502 5182 3554 5234
rect 4958 5182 5010 5234
rect 5854 5182 5906 5234
rect 8206 5182 8258 5234
rect 8878 5182 8930 5234
rect 9214 5182 9266 5234
rect 9886 5182 9938 5234
rect 12014 5182 12066 5234
rect 12462 5182 12514 5234
rect 15486 5182 15538 5234
rect 17054 5182 17106 5234
rect 20302 5182 20354 5234
rect 23326 5182 23378 5234
rect 25342 5182 25394 5234
rect 25678 5182 25730 5234
rect 30158 5182 30210 5234
rect 31726 5182 31778 5234
rect 33518 5182 33570 5234
rect 34526 5182 34578 5234
rect 35086 5182 35138 5234
rect 35534 5182 35586 5234
rect 35758 5182 35810 5234
rect 37102 5182 37154 5234
rect 43486 5182 43538 5234
rect 43710 5182 43762 5234
rect 53454 5182 53506 5234
rect 6638 5070 6690 5122
rect 9550 5070 9602 5122
rect 10446 5070 10498 5122
rect 10670 5070 10722 5122
rect 10782 5070 10834 5122
rect 11006 5070 11058 5122
rect 16718 5070 16770 5122
rect 17390 5070 17442 5122
rect 18286 5070 18338 5122
rect 19182 5070 19234 5122
rect 19518 5070 19570 5122
rect 22318 5070 22370 5122
rect 22654 5070 22706 5122
rect 23774 5070 23826 5122
rect 24222 5070 24274 5122
rect 25902 5070 25954 5122
rect 27582 5070 27634 5122
rect 28366 5070 28418 5122
rect 29374 5070 29426 5122
rect 31278 5070 31330 5122
rect 31502 5070 31554 5122
rect 32286 5070 32338 5122
rect 32510 5070 32562 5122
rect 33070 5070 33122 5122
rect 33966 5070 34018 5122
rect 34414 5070 34466 5122
rect 38782 5070 38834 5122
rect 39902 5070 39954 5122
rect 40686 5070 40738 5122
rect 41918 5070 41970 5122
rect 44830 5070 44882 5122
rect 46622 5070 46674 5122
rect 48526 5070 48578 5122
rect 48750 5070 48802 5122
rect 49758 5070 49810 5122
rect 51438 5070 51490 5122
rect 51662 5070 51714 5122
rect 51774 5070 51826 5122
rect 51998 5070 52050 5122
rect 53118 5070 53170 5122
rect 54014 5070 54066 5122
rect 54350 5070 54402 5122
rect 55918 5070 55970 5122
rect 56590 5070 56642 5122
rect 56926 5070 56978 5122
rect 4846 4958 4898 5010
rect 7870 4958 7922 5010
rect 9774 4958 9826 5010
rect 10222 4958 10274 5010
rect 11342 4958 11394 5010
rect 12798 4958 12850 5010
rect 13694 4958 13746 5010
rect 15150 4958 15202 5010
rect 16494 4958 16546 5010
rect 28590 4958 28642 5010
rect 30494 4958 30546 5010
rect 37550 4958 37602 5010
rect 39230 4958 39282 5010
rect 39678 4958 39730 5010
rect 40350 4958 40402 5010
rect 41022 4958 41074 5010
rect 41134 4958 41186 5010
rect 41694 4958 41746 5010
rect 42366 4958 42418 5010
rect 47182 4958 47234 5010
rect 49086 4958 49138 5010
rect 51102 4958 51154 5010
rect 51214 4958 51266 5010
rect 52670 4958 52722 5010
rect 54238 4958 54290 5010
rect 3950 4846 4002 4898
rect 4398 4846 4450 4898
rect 6414 4846 6466 4898
rect 11230 4846 11282 4898
rect 13582 4846 13634 4898
rect 32622 4846 32674 4898
rect 34190 4846 34242 4898
rect 34526 4846 34578 4898
rect 36094 4846 36146 4898
rect 42702 4846 42754 4898
rect 43710 4846 43762 4898
rect 45166 4846 45218 4898
rect 15520 4678 15572 4730
rect 15624 4678 15676 4730
rect 15728 4678 15780 4730
rect 29827 4678 29879 4730
rect 29931 4678 29983 4730
rect 30035 4678 30087 4730
rect 44134 4678 44186 4730
rect 44238 4678 44290 4730
rect 44342 4678 44394 4730
rect 58441 4678 58493 4730
rect 58545 4678 58597 4730
rect 58649 4678 58701 4730
rect 8990 4510 9042 4562
rect 10110 4510 10162 4562
rect 11342 4510 11394 4562
rect 15934 4510 15986 4562
rect 17726 4510 17778 4562
rect 24334 4510 24386 4562
rect 25454 4510 25506 4562
rect 33630 4510 33682 4562
rect 34078 4510 34130 4562
rect 35086 4510 35138 4562
rect 40238 4510 40290 4562
rect 46734 4510 46786 4562
rect 8094 4398 8146 4450
rect 8430 4398 8482 4450
rect 9886 4398 9938 4450
rect 10894 4398 10946 4450
rect 12126 4398 12178 4450
rect 12910 4398 12962 4450
rect 14030 4398 14082 4450
rect 14702 4398 14754 4450
rect 15038 4398 15090 4450
rect 18510 4398 18562 4450
rect 20414 4398 20466 4450
rect 20974 4398 21026 4450
rect 23998 4398 24050 4450
rect 24670 4398 24722 4450
rect 27134 4398 27186 4450
rect 28814 4398 28866 4450
rect 29486 4398 29538 4450
rect 30606 4398 30658 4450
rect 33854 4398 33906 4450
rect 38894 4398 38946 4450
rect 40126 4398 40178 4450
rect 43262 4398 43314 4450
rect 44606 4398 44658 4450
rect 51998 4398 52050 4450
rect 52222 4398 52274 4450
rect 4398 4286 4450 4338
rect 7646 4286 7698 4338
rect 10558 4286 10610 4338
rect 11454 4286 11506 4338
rect 11902 4286 11954 4338
rect 12686 4286 12738 4338
rect 13246 4286 13298 4338
rect 13806 4286 13858 4338
rect 15374 4286 15426 4338
rect 16718 4286 16770 4338
rect 17502 4286 17554 4338
rect 18062 4286 18114 4338
rect 19406 4286 19458 4338
rect 20862 4286 20914 4338
rect 21982 4286 22034 4338
rect 22766 4286 22818 4338
rect 25230 4286 25282 4338
rect 26238 4286 26290 4338
rect 26574 4286 26626 4338
rect 27806 4286 27858 4338
rect 28926 4286 28978 4338
rect 29822 4286 29874 4338
rect 30942 4286 30994 4338
rect 31950 4286 32002 4338
rect 33294 4286 33346 4338
rect 34190 4286 34242 4338
rect 38222 4286 38274 4338
rect 39342 4286 39394 4338
rect 40462 4286 40514 4338
rect 41134 4286 41186 4338
rect 42478 4286 42530 4338
rect 45390 4286 45442 4338
rect 47406 4286 47458 4338
rect 5070 4174 5122 4226
rect 7198 4174 7250 4226
rect 8878 4174 8930 4226
rect 10222 4174 10274 4226
rect 13694 4174 13746 4226
rect 16270 4174 16322 4226
rect 20974 4174 21026 4226
rect 22878 4174 22930 4226
rect 25566 4174 25618 4226
rect 26686 4174 26738 4226
rect 27582 4174 27634 4226
rect 28478 4174 28530 4226
rect 29934 4174 29986 4226
rect 32510 4174 32562 4226
rect 34638 4174 34690 4226
rect 37886 4174 37938 4226
rect 39118 4174 39170 4226
rect 41470 4174 41522 4226
rect 43934 4174 43986 4226
rect 47070 4174 47122 4226
rect 47854 4174 47906 4226
rect 51886 4174 51938 4226
rect 7758 4062 7810 4114
rect 11566 4062 11618 4114
rect 12238 4062 12290 4114
rect 8367 3894 8419 3946
rect 8471 3894 8523 3946
rect 8575 3894 8627 3946
rect 22674 3894 22726 3946
rect 22778 3894 22830 3946
rect 22882 3894 22934 3946
rect 36981 3894 37033 3946
rect 37085 3894 37137 3946
rect 37189 3894 37241 3946
rect 51288 3894 51340 3946
rect 51392 3894 51444 3946
rect 51496 3894 51548 3946
rect 16046 3726 16098 3778
rect 16382 3726 16434 3778
rect 28590 3726 28642 3778
rect 28926 3726 28978 3778
rect 29374 3726 29426 3778
rect 29710 3726 29762 3778
rect 38110 3726 38162 3778
rect 40798 3726 40850 3778
rect 6302 3614 6354 3666
rect 6750 3614 6802 3666
rect 7198 3614 7250 3666
rect 7646 3614 7698 3666
rect 9326 3614 9378 3666
rect 11454 3614 11506 3666
rect 13470 3614 13522 3666
rect 15822 3614 15874 3666
rect 16942 3614 16994 3666
rect 19070 3614 19122 3666
rect 20974 3614 21026 3666
rect 21758 3614 21810 3666
rect 23998 3614 24050 3666
rect 27806 3614 27858 3666
rect 29934 3614 29986 3666
rect 33406 3614 33458 3666
rect 34638 3614 34690 3666
rect 38558 3614 38610 3666
rect 41134 3614 41186 3666
rect 41918 3614 41970 3666
rect 47406 3614 47458 3666
rect 56590 3614 56642 3666
rect 57374 3614 57426 3666
rect 3166 3502 3218 3554
rect 4734 3502 4786 3554
rect 8094 3502 8146 3554
rect 12126 3502 12178 3554
rect 13694 3502 13746 3554
rect 14702 3502 14754 3554
rect 19854 3502 19906 3554
rect 21086 3502 21138 3554
rect 22430 3502 22482 3554
rect 22990 3502 23042 3554
rect 25006 3502 25058 3554
rect 28366 3502 28418 3554
rect 30606 3502 30658 3554
rect 35086 3502 35138 3554
rect 37662 3502 37714 3554
rect 38334 3502 38386 3554
rect 41470 3502 41522 3554
rect 42590 3502 42642 3554
rect 43486 3502 43538 3554
rect 43822 3502 43874 3554
rect 45054 3502 45106 3554
rect 45838 3502 45890 3554
rect 47518 3502 47570 3554
rect 47966 3502 48018 3554
rect 52782 3502 52834 3554
rect 56926 3502 56978 3554
rect 2718 3390 2770 3442
rect 2942 3390 2994 3442
rect 4958 3390 5010 3442
rect 5854 3390 5906 3442
rect 7870 3390 7922 3442
rect 8878 3390 8930 3442
rect 15262 3390 15314 3442
rect 25678 3390 25730 3442
rect 30942 3390 30994 3442
rect 31278 3390 31330 3442
rect 32510 3390 32562 3442
rect 32846 3390 32898 3442
rect 34190 3390 34242 3442
rect 37326 3390 37378 3442
rect 41022 3390 41074 3442
rect 42142 3390 42194 3442
rect 43710 3390 43762 3442
rect 45950 3390 46002 3442
rect 51998 3390 52050 3442
rect 52222 3390 52274 3442
rect 30270 3278 30322 3330
rect 33742 3278 33794 3330
rect 45054 3278 45106 3330
rect 15520 3110 15572 3162
rect 15624 3110 15676 3162
rect 15728 3110 15780 3162
rect 29827 3110 29879 3162
rect 29931 3110 29983 3162
rect 30035 3110 30087 3162
rect 44134 3110 44186 3162
rect 44238 3110 44290 3162
rect 44342 3110 44394 3162
rect 58441 3110 58493 3162
rect 58545 3110 58597 3162
rect 58649 3110 58701 3162
<< metal2 >>
rect 2912 39200 3024 40000
rect 5152 39200 5264 40000
rect 7392 39200 7504 40000
rect 7756 39228 8148 39284
rect 1820 36484 1876 36494
rect 1820 36390 1876 36428
rect 2492 36370 2548 36382
rect 2492 36318 2494 36370
rect 2546 36318 2548 36370
rect 1708 35698 1764 35710
rect 1708 35646 1710 35698
rect 1762 35646 1764 35698
rect 1708 35588 1764 35646
rect 1484 35364 1540 35374
rect 1372 34916 1428 34926
rect 1148 33796 1204 33806
rect 1036 29316 1092 29326
rect 1036 10836 1092 29260
rect 1148 14420 1204 33740
rect 1148 14354 1204 14364
rect 1260 28868 1316 28878
rect 1260 12852 1316 28812
rect 1372 16772 1428 34860
rect 1484 26068 1540 35308
rect 1708 35028 1764 35532
rect 2156 35586 2212 35598
rect 2156 35534 2158 35586
rect 2210 35534 2212 35586
rect 2156 35364 2212 35534
rect 2156 35298 2212 35308
rect 1708 34962 1764 34972
rect 1820 34914 1876 34926
rect 1820 34862 1822 34914
rect 1874 34862 1876 34914
rect 1820 34356 1876 34862
rect 2268 34916 2324 34926
rect 2268 34822 2324 34860
rect 2492 34356 2548 36318
rect 2604 36148 2660 36158
rect 2604 34914 2660 36092
rect 2940 35810 2996 39200
rect 2940 35758 2942 35810
rect 2994 35758 2996 35810
rect 2940 35746 2996 35758
rect 3500 37268 3556 37278
rect 2604 34862 2606 34914
rect 2658 34862 2660 34914
rect 2604 34692 2660 34862
rect 2604 34626 2660 34636
rect 3164 34914 3220 34926
rect 3164 34862 3166 34914
rect 3218 34862 3220 34914
rect 2716 34356 2772 34366
rect 2492 34354 2772 34356
rect 2492 34302 2718 34354
rect 2770 34302 2772 34354
rect 2492 34300 2772 34302
rect 1708 34132 1764 34142
rect 1596 34130 1764 34132
rect 1596 34078 1710 34130
rect 1762 34078 1764 34130
rect 1596 34076 1764 34078
rect 1596 33460 1652 34076
rect 1708 34066 1764 34076
rect 1708 33908 1764 33918
rect 1820 33908 1876 34300
rect 2716 34290 2772 34300
rect 3052 34244 3108 34254
rect 3052 34150 3108 34188
rect 2380 34132 2436 34142
rect 1764 33852 1876 33908
rect 2156 34018 2212 34030
rect 2156 33966 2158 34018
rect 2210 33966 2212 34018
rect 1708 33842 1764 33852
rect 1708 33460 1764 33470
rect 1596 33404 1708 33460
rect 1596 32788 1652 33404
rect 1708 33394 1764 33404
rect 1820 33348 1876 33358
rect 1820 33254 1876 33292
rect 2156 32788 2212 33966
rect 1596 32722 1652 32732
rect 2044 32732 2212 32788
rect 1820 32676 1876 32686
rect 1820 32582 1876 32620
rect 1932 32674 1988 32686
rect 1932 32622 1934 32674
rect 1986 32622 1988 32674
rect 1932 32452 1988 32622
rect 1820 32396 1988 32452
rect 1484 26002 1540 26012
rect 1596 32116 1652 32126
rect 1820 32116 1876 32396
rect 1820 32060 1988 32116
rect 1596 21924 1652 32060
rect 1820 31780 1876 31790
rect 1820 31686 1876 31724
rect 1708 30996 1764 31006
rect 1708 30548 1764 30940
rect 1708 30482 1764 30492
rect 1708 30100 1764 30110
rect 1708 28308 1764 30044
rect 1708 28242 1764 28252
rect 1820 29426 1876 29438
rect 1820 29374 1822 29426
rect 1874 29374 1876 29426
rect 1820 28420 1876 29374
rect 1932 29316 1988 32060
rect 2044 30772 2100 32732
rect 2380 32674 2436 34076
rect 2716 33908 2772 33918
rect 2492 33234 2548 33246
rect 2492 33182 2494 33234
rect 2546 33182 2548 33234
rect 2492 32786 2548 33182
rect 2492 32734 2494 32786
rect 2546 32734 2548 32786
rect 2492 32722 2548 32734
rect 2380 32622 2382 32674
rect 2434 32622 2436 32674
rect 2380 32610 2436 32622
rect 2716 32674 2772 33852
rect 2716 32622 2718 32674
rect 2770 32622 2772 32674
rect 2716 32610 2772 32622
rect 3052 33124 3108 33134
rect 2156 32564 2212 32574
rect 2156 32562 2324 32564
rect 2156 32510 2158 32562
rect 2210 32510 2324 32562
rect 2156 32508 2324 32510
rect 2156 32498 2212 32508
rect 2268 32340 2324 32508
rect 2268 32274 2324 32284
rect 2940 32562 2996 32574
rect 2940 32510 2942 32562
rect 2994 32510 2996 32562
rect 2940 32004 2996 32510
rect 2940 31938 2996 31948
rect 2828 31892 2884 31902
rect 2268 31778 2324 31790
rect 2268 31726 2270 31778
rect 2322 31726 2324 31778
rect 2268 31220 2324 31726
rect 2268 31154 2324 31164
rect 2716 31554 2772 31566
rect 2716 31502 2718 31554
rect 2770 31502 2772 31554
rect 2268 30882 2324 30894
rect 2268 30830 2270 30882
rect 2322 30830 2324 30882
rect 2044 30716 2212 30772
rect 2044 30548 2100 30558
rect 2044 30098 2100 30492
rect 2044 30046 2046 30098
rect 2098 30046 2100 30098
rect 2044 30034 2100 30046
rect 1932 29250 1988 29260
rect 2156 29092 2212 30716
rect 2268 30436 2324 30830
rect 2268 30370 2324 30380
rect 2492 30324 2548 30334
rect 2380 30268 2492 30324
rect 2380 30212 2436 30268
rect 2492 30258 2548 30268
rect 2156 29026 2212 29036
rect 2268 30156 2436 30212
rect 2268 28980 2324 30156
rect 2492 30100 2548 30110
rect 2716 30100 2772 31502
rect 2828 30994 2884 31836
rect 2828 30942 2830 30994
rect 2882 30942 2884 30994
rect 2828 30930 2884 30942
rect 2940 31554 2996 31566
rect 2940 31502 2942 31554
rect 2994 31502 2996 31554
rect 2940 30436 2996 31502
rect 2548 30044 2772 30100
rect 2828 30380 2996 30436
rect 2492 30034 2548 30044
rect 2380 29988 2436 29998
rect 2380 29428 2436 29932
rect 2380 29362 2436 29372
rect 2604 29314 2660 29326
rect 2604 29262 2606 29314
rect 2658 29262 2660 29314
rect 2604 29204 2660 29262
rect 2604 29138 2660 29148
rect 2268 28924 2548 28980
rect 1708 28084 1764 28094
rect 1820 28084 1876 28364
rect 1708 28082 1876 28084
rect 1708 28030 1710 28082
rect 1762 28030 1876 28082
rect 1708 28028 1876 28030
rect 1932 28644 1988 28654
rect 2156 28644 2212 28654
rect 1932 28642 2212 28644
rect 1932 28590 1934 28642
rect 1986 28590 2158 28642
rect 2210 28590 2212 28642
rect 1932 28588 2212 28590
rect 1708 27074 1764 28028
rect 1708 27022 1710 27074
rect 1762 27022 1764 27074
rect 1708 27010 1764 27022
rect 1820 27188 1876 27198
rect 1820 26290 1876 27132
rect 1820 26238 1822 26290
rect 1874 26238 1876 26290
rect 1820 26226 1876 26238
rect 1596 21858 1652 21868
rect 1708 24276 1764 24286
rect 1372 16706 1428 16716
rect 1484 21252 1540 21262
rect 1484 14308 1540 21196
rect 1708 20468 1764 24220
rect 1932 23492 1988 28588
rect 2156 28578 2212 28588
rect 2492 28532 2548 28924
rect 2828 28642 2884 30380
rect 2940 30210 2996 30222
rect 2940 30158 2942 30210
rect 2994 30158 2996 30210
rect 2940 29540 2996 30158
rect 3052 29988 3108 33068
rect 3164 32116 3220 34862
rect 3500 34916 3556 37212
rect 5180 36820 5236 39200
rect 7420 39060 7476 39200
rect 7756 39060 7812 39228
rect 7420 39004 7812 39060
rect 5180 36764 5796 36820
rect 4620 36596 4676 36606
rect 4620 36502 4676 36540
rect 5404 36596 5460 36606
rect 4172 36484 4228 36494
rect 3836 35698 3892 35710
rect 3836 35646 3838 35698
rect 3890 35646 3892 35698
rect 3836 35364 3892 35646
rect 4172 35700 4228 36428
rect 4956 35924 5012 35934
rect 4956 35810 5012 35868
rect 4956 35758 4958 35810
rect 5010 35758 5012 35810
rect 4956 35746 5012 35758
rect 4172 35606 4228 35644
rect 5068 35700 5124 35710
rect 3836 35298 3892 35308
rect 5068 35026 5124 35644
rect 5068 34974 5070 35026
rect 5122 34974 5124 35026
rect 5068 34962 5124 34974
rect 3500 34822 3556 34860
rect 4060 34916 4116 34926
rect 4060 34822 4116 34860
rect 5180 34916 5236 34926
rect 5236 34860 5348 34916
rect 5180 34850 5236 34860
rect 4620 34692 4676 34702
rect 4620 34690 4900 34692
rect 4620 34638 4622 34690
rect 4674 34638 4900 34690
rect 4620 34636 4900 34638
rect 4620 34626 4676 34636
rect 4060 34356 4116 34366
rect 4060 34354 4564 34356
rect 4060 34302 4062 34354
rect 4114 34302 4564 34354
rect 4060 34300 4564 34302
rect 4060 34290 4116 34300
rect 3500 34242 3556 34254
rect 3500 34190 3502 34242
rect 3554 34190 3556 34242
rect 3388 34130 3444 34142
rect 3388 34078 3390 34130
rect 3442 34078 3444 34130
rect 3164 32050 3220 32060
rect 3276 33348 3332 33358
rect 3276 32562 3332 33292
rect 3388 32676 3444 34078
rect 3500 33796 3556 34190
rect 3500 33730 3556 33740
rect 3724 34130 3780 34142
rect 3724 34078 3726 34130
rect 3778 34078 3780 34130
rect 3724 33012 3780 34078
rect 4172 34130 4228 34142
rect 4172 34078 4174 34130
rect 4226 34078 4228 34130
rect 4060 33908 4116 33918
rect 4060 33814 4116 33852
rect 3724 32946 3780 32956
rect 4172 32900 4228 34078
rect 4396 34132 4452 34142
rect 4396 34038 4452 34076
rect 4508 33460 4564 34300
rect 4620 34242 4676 34254
rect 4620 34190 4622 34242
rect 4674 34190 4676 34242
rect 4620 33796 4676 34190
rect 4620 33730 4676 33740
rect 4732 34130 4788 34142
rect 4732 34078 4734 34130
rect 4786 34078 4788 34130
rect 4620 33460 4676 33470
rect 4508 33458 4676 33460
rect 4508 33406 4622 33458
rect 4674 33406 4676 33458
rect 4508 33404 4676 33406
rect 4620 33348 4676 33404
rect 4620 33282 4676 33292
rect 4172 32834 4228 32844
rect 3444 32620 3556 32676
rect 3388 32610 3444 32620
rect 3276 32510 3278 32562
rect 3330 32510 3332 32562
rect 3276 31892 3332 32510
rect 3276 31826 3332 31836
rect 3276 31668 3332 31678
rect 3164 31554 3220 31566
rect 3164 31502 3166 31554
rect 3218 31502 3220 31554
rect 3164 30772 3220 31502
rect 3164 30706 3220 30716
rect 3276 30436 3332 31612
rect 3052 29922 3108 29932
rect 3164 30380 3332 30436
rect 2940 29474 2996 29484
rect 3052 29204 3108 29214
rect 3052 28754 3108 29148
rect 3052 28702 3054 28754
rect 3106 28702 3108 28754
rect 3052 28690 3108 28702
rect 2828 28590 2830 28642
rect 2882 28590 2884 28642
rect 2828 28578 2884 28590
rect 3164 28532 3220 30380
rect 3500 30212 3556 32620
rect 3948 32564 4004 32574
rect 3836 32004 3892 32014
rect 3836 31778 3892 31948
rect 3836 31726 3838 31778
rect 3890 31726 3892 31778
rect 3836 31714 3892 31726
rect 3948 31778 4004 32508
rect 3948 31726 3950 31778
rect 4002 31726 4004 31778
rect 3948 31714 4004 31726
rect 4060 32450 4116 32462
rect 4060 32398 4062 32450
rect 4114 32398 4116 32450
rect 4060 31554 4116 32398
rect 4060 31502 4062 31554
rect 4114 31502 4116 31554
rect 4060 31490 4116 31502
rect 4172 32340 4228 32350
rect 4172 31108 4228 32284
rect 4620 31892 4676 31902
rect 4284 31668 4340 31678
rect 4284 31666 4564 31668
rect 4284 31614 4286 31666
rect 4338 31614 4564 31666
rect 4284 31612 4564 31614
rect 4284 31602 4340 31612
rect 4172 31052 4452 31108
rect 3612 30884 3668 30894
rect 3612 30882 4340 30884
rect 3612 30830 3614 30882
rect 3666 30830 4340 30882
rect 3612 30828 4340 30830
rect 3612 30818 3668 30828
rect 3612 30212 3668 30222
rect 3388 30210 3668 30212
rect 3388 30158 3614 30210
rect 3666 30158 3668 30210
rect 3388 30156 3668 30158
rect 3276 28644 3332 28654
rect 3276 28550 3332 28588
rect 2380 28530 2548 28532
rect 2380 28478 2494 28530
rect 2546 28478 2548 28530
rect 2380 28476 2548 28478
rect 2380 28420 2436 28476
rect 2492 28466 2548 28476
rect 2940 28476 3220 28532
rect 3388 28532 3444 30156
rect 3612 30146 3668 30156
rect 3724 29986 3780 29998
rect 3724 29934 3726 29986
rect 3778 29934 3780 29986
rect 3724 29876 3780 29934
rect 3948 29988 4004 29998
rect 4284 29988 4340 30828
rect 4396 30210 4452 31052
rect 4396 30158 4398 30210
rect 4450 30158 4452 30210
rect 4396 30146 4452 30158
rect 4508 30212 4564 31612
rect 4620 31666 4676 31836
rect 4620 31614 4622 31666
rect 4674 31614 4676 31666
rect 4620 31602 4676 31614
rect 4732 31668 4788 34078
rect 4732 31602 4788 31612
rect 4508 30146 4564 30156
rect 4620 30772 4676 30782
rect 4844 30772 4900 34636
rect 5180 33122 5236 33134
rect 5180 33070 5182 33122
rect 5234 33070 5236 33122
rect 5180 32004 5236 33070
rect 4676 30716 4900 30772
rect 4956 31666 5012 31678
rect 4956 31614 4958 31666
rect 5010 31614 5012 31666
rect 4956 31108 5012 31614
rect 5180 31556 5236 31948
rect 5292 31948 5348 34860
rect 5404 34354 5460 36540
rect 5628 35364 5684 35374
rect 5628 35026 5684 35308
rect 5628 34974 5630 35026
rect 5682 34974 5684 35026
rect 5628 34962 5684 34974
rect 5404 34302 5406 34354
rect 5458 34302 5460 34354
rect 5404 34290 5460 34302
rect 5740 34020 5796 36764
rect 5852 36482 5908 36494
rect 5852 36430 5854 36482
rect 5906 36430 5908 36482
rect 5852 35700 5908 36430
rect 6636 36372 6692 36382
rect 6636 36278 6692 36316
rect 7868 36372 7924 36382
rect 6972 35812 7028 35822
rect 5852 35634 5908 35644
rect 6860 35756 6972 35812
rect 6636 34356 6692 34366
rect 6636 34262 6692 34300
rect 5852 34020 5908 34030
rect 5740 34018 5908 34020
rect 5740 33966 5854 34018
rect 5906 33966 5908 34018
rect 5740 33964 5908 33966
rect 5852 33954 5908 33964
rect 6188 33460 6244 33470
rect 6188 33366 6244 33404
rect 5852 33122 5908 33134
rect 6636 33124 6692 33134
rect 5852 33070 5854 33122
rect 5906 33070 5908 33122
rect 5852 31948 5908 33070
rect 6300 33122 6692 33124
rect 6300 33070 6638 33122
rect 6690 33070 6692 33122
rect 6300 33068 6692 33070
rect 6300 32676 6356 33068
rect 6636 33058 6692 33068
rect 6748 32900 6804 32910
rect 6636 32676 6692 32686
rect 6076 32620 6356 32676
rect 6524 32674 6692 32676
rect 6524 32622 6638 32674
rect 6690 32622 6692 32674
rect 6524 32620 6692 32622
rect 5292 31892 5460 31948
rect 5740 31892 5908 31948
rect 5964 32452 6020 32462
rect 5180 31490 5236 31500
rect 4508 29988 4564 29998
rect 4284 29986 4564 29988
rect 4284 29934 4510 29986
rect 4562 29934 4564 29986
rect 4284 29932 4564 29934
rect 3948 29894 4004 29932
rect 4508 29922 4564 29932
rect 3724 28868 3780 29820
rect 3724 28802 3780 28812
rect 3948 28868 4004 28878
rect 3724 28644 3780 28654
rect 3724 28550 3780 28588
rect 2044 28364 2436 28420
rect 2044 27970 2100 28364
rect 2716 28084 2772 28094
rect 2940 28084 2996 28476
rect 3388 28420 3444 28476
rect 2716 28082 2996 28084
rect 2716 28030 2718 28082
rect 2770 28030 2996 28082
rect 2716 28028 2996 28030
rect 3052 28364 3444 28420
rect 3500 28530 3556 28542
rect 3500 28478 3502 28530
rect 3554 28478 3556 28530
rect 3052 28082 3108 28364
rect 3052 28030 3054 28082
rect 3106 28030 3108 28082
rect 2716 28018 2772 28028
rect 3052 28018 3108 28030
rect 2044 27918 2046 27970
rect 2098 27918 2100 27970
rect 2044 27906 2100 27918
rect 2380 27858 2436 27870
rect 3276 27860 3332 27870
rect 2380 27806 2382 27858
rect 2434 27806 2436 27858
rect 2380 26908 2436 27806
rect 3164 27858 3332 27860
rect 3164 27806 3278 27858
rect 3330 27806 3332 27858
rect 3164 27804 3332 27806
rect 2268 26852 2436 26908
rect 2492 26962 2548 26974
rect 2492 26910 2494 26962
rect 2546 26910 2548 26962
rect 2492 26908 2548 26910
rect 2492 26852 3108 26908
rect 2044 26402 2100 26414
rect 2044 26350 2046 26402
rect 2098 26350 2100 26402
rect 2044 25732 2100 26350
rect 2044 25666 2100 25676
rect 2044 25506 2100 25518
rect 2044 25454 2046 25506
rect 2098 25454 2100 25506
rect 2044 24948 2100 25454
rect 2156 24948 2212 24958
rect 2044 24892 2156 24948
rect 2156 24854 2212 24892
rect 2268 24164 2324 26852
rect 2492 26740 2548 26750
rect 2492 26514 2548 26684
rect 2492 26462 2494 26514
rect 2546 26462 2548 26514
rect 2492 26450 2548 26462
rect 3052 26514 3108 26852
rect 3052 26462 3054 26514
rect 3106 26462 3108 26514
rect 3052 26450 3108 26462
rect 2828 26292 2884 26302
rect 2268 24098 2324 24108
rect 2380 26290 2884 26292
rect 2380 26238 2830 26290
rect 2882 26238 2884 26290
rect 2380 26236 2884 26238
rect 2044 23940 2100 23950
rect 2044 23938 2324 23940
rect 2044 23886 2046 23938
rect 2098 23886 2324 23938
rect 2044 23884 2324 23886
rect 2044 23874 2100 23884
rect 1820 23154 1876 23166
rect 1820 23102 1822 23154
rect 1874 23102 1876 23154
rect 1820 21812 1876 23102
rect 1820 20814 1876 21756
rect 1820 20762 1822 20814
rect 1874 20762 1876 20814
rect 1820 20750 1876 20762
rect 1932 21812 1988 23436
rect 2156 23716 2212 23726
rect 2156 21924 2212 23660
rect 2268 23604 2324 23884
rect 2380 23938 2436 26236
rect 2828 26226 2884 26236
rect 3164 25620 3220 27804
rect 3276 27794 3332 27804
rect 3500 26402 3556 28478
rect 3948 28530 4004 28812
rect 3948 28478 3950 28530
rect 4002 28478 4004 28530
rect 3948 28466 4004 28478
rect 4060 28532 4116 28542
rect 4396 28532 4452 28542
rect 4060 28530 4228 28532
rect 4060 28478 4062 28530
rect 4114 28478 4228 28530
rect 4060 28476 4228 28478
rect 4060 28466 4116 28476
rect 4060 28196 4116 28206
rect 4060 27858 4116 28140
rect 4172 27972 4228 28476
rect 4396 28438 4452 28476
rect 4508 28420 4564 28430
rect 4620 28420 4676 30716
rect 4956 30324 5012 31052
rect 4956 30258 5012 30268
rect 5068 30996 5124 31006
rect 4732 30100 4788 30110
rect 4732 30006 4788 30044
rect 4956 30098 5012 30110
rect 4956 30046 4958 30098
rect 5010 30046 5012 30098
rect 4732 29314 4788 29326
rect 4732 29262 4734 29314
rect 4786 29262 4788 29314
rect 4732 28868 4788 29262
rect 4956 29092 5012 30046
rect 4956 29026 5012 29036
rect 4732 28802 4788 28812
rect 5068 28754 5124 30940
rect 5068 28702 5070 28754
rect 5122 28702 5124 28754
rect 5068 28690 5124 28702
rect 5180 30548 5236 30558
rect 4732 28644 4788 28654
rect 4732 28550 4788 28588
rect 4508 28418 4676 28420
rect 4508 28366 4510 28418
rect 4562 28366 4676 28418
rect 4508 28364 4676 28366
rect 4284 27972 4340 27982
rect 4172 27970 4340 27972
rect 4172 27918 4286 27970
rect 4338 27918 4340 27970
rect 4172 27916 4340 27918
rect 4060 27806 4062 27858
rect 4114 27806 4116 27858
rect 4060 27794 4116 27806
rect 3500 26350 3502 26402
rect 3554 26350 3556 26402
rect 3276 26292 3332 26302
rect 3276 26198 3332 26236
rect 2604 25564 3220 25620
rect 2492 24722 2548 24734
rect 2492 24670 2494 24722
rect 2546 24670 2548 24722
rect 2492 24500 2548 24670
rect 2492 24434 2548 24444
rect 2604 24052 2660 25564
rect 2716 25396 2772 25406
rect 2716 25394 3220 25396
rect 2716 25342 2718 25394
rect 2770 25342 3220 25394
rect 2716 25340 3220 25342
rect 2716 25330 2772 25340
rect 3164 24946 3220 25340
rect 3164 24894 3166 24946
rect 3218 24894 3220 24946
rect 3164 24882 3220 24894
rect 3388 25172 3444 25182
rect 3388 24834 3444 25116
rect 3388 24782 3390 24834
rect 3442 24782 3444 24834
rect 3388 24770 3444 24782
rect 2380 23886 2382 23938
rect 2434 23886 2436 23938
rect 2380 23874 2436 23886
rect 2492 23996 2660 24052
rect 3052 24722 3108 24734
rect 3052 24670 3054 24722
rect 3106 24670 3108 24722
rect 2268 23538 2324 23548
rect 2492 23380 2548 23996
rect 3052 23938 3108 24670
rect 3164 24724 3220 24734
rect 3220 24668 3332 24724
rect 3164 24658 3220 24668
rect 3276 24276 3332 24668
rect 3052 23886 3054 23938
rect 3106 23886 3108 23938
rect 3052 23874 3108 23886
rect 3164 24164 3220 24174
rect 2604 23826 2660 23838
rect 2604 23774 2606 23826
rect 2658 23774 2660 23826
rect 2604 23604 2660 23774
rect 2716 23716 2772 23726
rect 2828 23716 2884 23726
rect 2716 23714 2828 23716
rect 2716 23662 2718 23714
rect 2770 23662 2828 23714
rect 2716 23660 2828 23662
rect 2716 23650 2772 23660
rect 2604 23492 2772 23548
rect 2268 23324 2548 23380
rect 2268 22372 2324 23324
rect 2492 23044 2548 23054
rect 2492 22950 2548 22988
rect 2268 22316 2548 22372
rect 2268 22148 2324 22158
rect 2268 22146 2436 22148
rect 2268 22094 2270 22146
rect 2322 22094 2436 22146
rect 2268 22092 2436 22094
rect 2268 22082 2324 22092
rect 2380 21924 2436 22092
rect 2492 22036 2548 22316
rect 2604 22260 2660 22270
rect 2604 22166 2660 22204
rect 2492 21980 2660 22036
rect 2156 21868 2324 21924
rect 2380 21868 2548 21924
rect 1932 21810 2212 21812
rect 1932 21758 1934 21810
rect 1986 21758 2212 21810
rect 1932 21756 2212 21758
rect 1932 20692 1988 21756
rect 2156 21698 2212 21756
rect 2156 21646 2158 21698
rect 2210 21646 2212 21698
rect 2156 21634 2212 21646
rect 2268 21700 2324 21868
rect 2492 21700 2548 21868
rect 2268 21644 2436 21700
rect 1708 20402 1764 20412
rect 1820 20636 1988 20692
rect 2268 21364 2324 21374
rect 1820 20244 1876 20636
rect 2044 20468 2100 20478
rect 2100 20412 2212 20468
rect 2044 20402 2100 20412
rect 1932 20244 1988 20254
rect 1820 20242 1988 20244
rect 1820 20190 1934 20242
rect 1986 20190 1988 20242
rect 1820 20188 1988 20190
rect 1932 20178 1988 20188
rect 1708 20020 1764 20030
rect 1764 19964 1876 20020
rect 1708 19954 1764 19964
rect 1708 19236 1764 19246
rect 1708 19142 1764 19180
rect 1820 18450 1876 19964
rect 2044 19908 2100 19918
rect 1820 18398 1822 18450
rect 1874 18398 1876 18450
rect 1820 18386 1876 18398
rect 1932 19236 1988 19246
rect 1708 18228 1764 18238
rect 1708 17668 1764 18172
rect 1708 17574 1764 17612
rect 1708 16882 1764 16894
rect 1708 16830 1710 16882
rect 1762 16830 1764 16882
rect 1708 15988 1764 16830
rect 1820 16884 1876 16894
rect 1820 16098 1876 16828
rect 1820 16046 1822 16098
rect 1874 16046 1876 16098
rect 1820 16034 1876 16046
rect 1708 15922 1764 15932
rect 1820 15316 1876 15326
rect 1932 15316 1988 19180
rect 2044 18674 2100 19852
rect 2044 18622 2046 18674
rect 2098 18622 2100 18674
rect 2044 18610 2100 18622
rect 2044 17556 2100 17566
rect 2156 17556 2212 20412
rect 2268 20130 2324 21308
rect 2268 20078 2270 20130
rect 2322 20078 2324 20130
rect 2268 20066 2324 20078
rect 2044 17554 2212 17556
rect 2044 17502 2046 17554
rect 2098 17502 2212 17554
rect 2044 17500 2212 17502
rect 2380 17554 2436 21644
rect 2492 21606 2548 21644
rect 2604 21140 2660 21980
rect 2716 21812 2772 23492
rect 2828 22036 2884 23660
rect 2940 23714 2996 23726
rect 2940 23662 2942 23714
rect 2994 23662 2996 23714
rect 2940 22370 2996 23662
rect 3052 23044 3108 23054
rect 3052 22482 3108 22988
rect 3052 22430 3054 22482
rect 3106 22430 3108 22482
rect 3052 22418 3108 22430
rect 2940 22318 2942 22370
rect 2994 22318 2996 22370
rect 2940 22306 2996 22318
rect 2828 21970 2884 21980
rect 2828 21812 2884 21822
rect 2716 21810 2884 21812
rect 2716 21758 2830 21810
rect 2882 21758 2884 21810
rect 2716 21756 2884 21758
rect 2828 21140 2884 21756
rect 3164 21810 3220 24108
rect 3276 23826 3332 24220
rect 3500 24722 3556 26350
rect 4060 26402 4116 26414
rect 4060 26350 4062 26402
rect 4114 26350 4116 26402
rect 3836 26292 3892 26302
rect 3836 26290 4004 26292
rect 3836 26238 3838 26290
rect 3890 26238 4004 26290
rect 3836 26236 4004 26238
rect 3836 26226 3892 26236
rect 3948 25172 4004 26236
rect 4060 25620 4116 26350
rect 4060 25554 4116 25564
rect 4172 26292 4228 26302
rect 4284 26292 4340 27916
rect 4508 27860 4564 28364
rect 4732 28196 4788 28206
rect 4732 28082 4788 28140
rect 4732 28030 4734 28082
rect 4786 28030 4788 28082
rect 4732 28018 4788 28030
rect 5180 27972 5236 30492
rect 5068 27916 5236 27972
rect 5292 29426 5348 29438
rect 5292 29374 5294 29426
rect 5346 29374 5348 29426
rect 5292 28420 5348 29374
rect 5404 28420 5460 31892
rect 5516 31836 5796 31892
rect 5516 29876 5572 31836
rect 5628 31668 5684 31678
rect 5628 30210 5684 31612
rect 5740 31666 5796 31836
rect 5964 31778 6020 32396
rect 5964 31726 5966 31778
rect 6018 31726 6020 31778
rect 5964 31714 6020 31726
rect 6076 31780 6132 32620
rect 6412 32564 6468 32574
rect 6412 32470 6468 32508
rect 6188 32450 6244 32462
rect 6188 32398 6190 32450
rect 6242 32398 6244 32450
rect 6188 31948 6244 32398
rect 6524 31948 6580 32620
rect 6636 32610 6692 32620
rect 6748 32674 6804 32844
rect 6748 32622 6750 32674
rect 6802 32622 6804 32674
rect 6748 32610 6804 32622
rect 6860 31948 6916 35756
rect 6972 35746 7028 35756
rect 7644 35700 7700 35710
rect 7084 35698 7700 35700
rect 7084 35646 7646 35698
rect 7698 35646 7700 35698
rect 7084 35644 7700 35646
rect 7084 35586 7140 35644
rect 7644 35634 7700 35644
rect 7084 35534 7086 35586
rect 7138 35534 7140 35586
rect 7084 35522 7140 35534
rect 7756 34804 7812 34814
rect 6972 34802 7812 34804
rect 6972 34750 7758 34802
rect 7810 34750 7812 34802
rect 6972 34748 7812 34750
rect 6972 34354 7028 34748
rect 7756 34738 7812 34748
rect 6972 34302 6974 34354
rect 7026 34302 7028 34354
rect 6972 34290 7028 34302
rect 7868 34354 7924 36316
rect 8092 35586 8148 39228
rect 9632 39200 9744 40000
rect 11872 39200 11984 40000
rect 14112 39200 14224 40000
rect 14476 39228 14868 39284
rect 9660 36932 9716 39200
rect 8365 36876 8629 36886
rect 8421 36820 8469 36876
rect 8525 36820 8573 36876
rect 9660 36866 9716 36876
rect 10668 36932 10724 36942
rect 8365 36810 8629 36820
rect 8764 36652 9940 36708
rect 8764 36594 8820 36652
rect 8764 36542 8766 36594
rect 8818 36542 8820 36594
rect 8764 36530 8820 36542
rect 9772 36482 9828 36494
rect 9772 36430 9774 36482
rect 9826 36430 9828 36482
rect 8092 35534 8094 35586
rect 8146 35534 8148 35586
rect 8092 35522 8148 35534
rect 8876 35586 8932 35598
rect 8876 35534 8878 35586
rect 8930 35534 8932 35586
rect 8876 35476 8932 35534
rect 8876 35410 8932 35420
rect 8988 35588 9044 35598
rect 8365 35308 8629 35318
rect 8421 35252 8469 35308
rect 8525 35252 8573 35308
rect 8365 35242 8629 35252
rect 8540 34916 8596 34926
rect 8988 34916 9044 35532
rect 9772 35588 9828 36430
rect 9884 35922 9940 36652
rect 9884 35870 9886 35922
rect 9938 35870 9940 35922
rect 9884 35858 9940 35870
rect 10444 36370 10500 36382
rect 10444 36318 10446 36370
rect 10498 36318 10500 36370
rect 9772 35522 9828 35532
rect 10444 35364 10500 36318
rect 10668 35922 10724 36876
rect 10668 35870 10670 35922
rect 10722 35870 10724 35922
rect 10668 35858 10724 35870
rect 11228 36820 11284 36830
rect 11116 35588 11172 35598
rect 11116 35494 11172 35532
rect 10444 35298 10500 35308
rect 8540 34914 9044 34916
rect 8540 34862 8542 34914
rect 8594 34862 8990 34914
rect 9042 34862 9044 34914
rect 8540 34860 9044 34862
rect 8540 34850 8596 34860
rect 7868 34302 7870 34354
rect 7922 34302 7924 34354
rect 7868 34290 7924 34302
rect 8764 34354 8820 34860
rect 8988 34850 9044 34860
rect 9660 34804 9716 34814
rect 9660 34802 9940 34804
rect 9660 34750 9662 34802
rect 9714 34750 9940 34802
rect 9660 34748 9940 34750
rect 9660 34738 9716 34748
rect 8764 34302 8766 34354
rect 8818 34302 8820 34354
rect 8764 34290 8820 34302
rect 9884 34354 9940 34748
rect 9884 34302 9886 34354
rect 9938 34302 9940 34354
rect 9884 34290 9940 34302
rect 9996 34692 10052 34702
rect 7308 34130 7364 34142
rect 7308 34078 7310 34130
rect 7362 34078 7364 34130
rect 7084 33124 7140 33134
rect 7308 33124 7364 34078
rect 8204 34132 8260 34142
rect 8204 34038 8260 34076
rect 8365 33740 8629 33750
rect 8421 33684 8469 33740
rect 8525 33684 8573 33740
rect 8365 33674 8629 33684
rect 8876 33572 8932 33582
rect 8204 33460 8260 33470
rect 8204 33366 8260 33404
rect 8540 33348 8596 33358
rect 7532 33124 7588 33134
rect 7308 33122 7700 33124
rect 7308 33070 7534 33122
rect 7586 33070 7700 33122
rect 7308 33068 7700 33070
rect 7084 33030 7140 33068
rect 7532 33058 7588 33068
rect 7196 32900 7252 32910
rect 7196 32786 7252 32844
rect 7196 32734 7198 32786
rect 7250 32734 7252 32786
rect 6188 31892 6580 31948
rect 6524 31826 6580 31836
rect 6748 31892 6916 31948
rect 6972 32676 7028 32686
rect 6076 31714 6132 31724
rect 5740 31614 5742 31666
rect 5794 31614 5796 31666
rect 5740 31602 5796 31614
rect 6636 31666 6692 31678
rect 6636 31614 6638 31666
rect 6690 31614 6692 31666
rect 6188 30996 6244 31006
rect 6188 30902 6244 30940
rect 5740 30882 5796 30894
rect 5740 30830 5742 30882
rect 5794 30830 5796 30882
rect 5740 30772 5796 30830
rect 6636 30772 6692 31614
rect 5740 30716 6692 30772
rect 5628 30158 5630 30210
rect 5682 30158 5684 30210
rect 5628 30146 5684 30158
rect 5964 30212 6020 30222
rect 5964 30118 6020 30156
rect 6412 30100 6468 30110
rect 6412 30006 6468 30044
rect 6636 30098 6692 30716
rect 6748 30660 6804 31892
rect 6972 31666 7028 32620
rect 7196 32340 7252 32734
rect 7196 32274 7252 32284
rect 7644 32004 7700 33068
rect 7644 31938 7700 31948
rect 7756 33012 7812 33022
rect 7196 31892 7252 31902
rect 7196 31798 7252 31836
rect 7532 31892 7588 31902
rect 7532 31798 7588 31836
rect 6972 31614 6974 31666
rect 7026 31614 7028 31666
rect 6972 30996 7028 31614
rect 6972 30940 7252 30996
rect 6860 30882 6916 30894
rect 6860 30830 6862 30882
rect 6914 30830 6916 30882
rect 6860 30772 6916 30830
rect 7196 30772 7252 30940
rect 6860 30716 7028 30772
rect 6748 30604 6916 30660
rect 6636 30046 6638 30098
rect 6690 30046 6692 30098
rect 6636 30034 6692 30046
rect 6748 30324 6804 30334
rect 6748 30098 6804 30268
rect 6748 30046 6750 30098
rect 6802 30046 6804 30098
rect 5740 29988 5796 29998
rect 5516 29810 5572 29820
rect 5628 29986 5796 29988
rect 5628 29934 5742 29986
rect 5794 29934 5796 29986
rect 5628 29932 5796 29934
rect 5516 29316 5572 29326
rect 5628 29316 5684 29932
rect 5740 29876 5796 29932
rect 5740 29810 5796 29820
rect 6076 29316 6132 29326
rect 5572 29260 5684 29316
rect 5740 29314 6132 29316
rect 5740 29262 6078 29314
rect 6130 29262 6132 29314
rect 5740 29260 6132 29262
rect 5516 29250 5572 29260
rect 5740 28754 5796 29260
rect 6076 29250 6132 29260
rect 5740 28702 5742 28754
rect 5794 28702 5796 28754
rect 5740 28690 5796 28702
rect 6076 29092 6132 29102
rect 5516 28644 5572 28654
rect 5516 28550 5572 28588
rect 5964 28644 6020 28654
rect 5964 28550 6020 28588
rect 6076 28642 6132 29036
rect 6748 28868 6804 30046
rect 6076 28590 6078 28642
rect 6130 28590 6132 28642
rect 6076 28578 6132 28590
rect 6636 28812 6804 28868
rect 5852 28420 5908 28430
rect 5404 28364 5572 28420
rect 4508 27804 4788 27860
rect 4732 27634 4788 27804
rect 4732 27582 4734 27634
rect 4786 27582 4788 27634
rect 4620 27186 4676 27198
rect 4620 27134 4622 27186
rect 4674 27134 4676 27186
rect 4620 26404 4676 27134
rect 4620 26310 4676 26348
rect 4508 26292 4564 26302
rect 4172 26290 4564 26292
rect 4172 26238 4174 26290
rect 4226 26238 4510 26290
rect 4562 26238 4564 26290
rect 4172 26236 4564 26238
rect 3948 25106 4004 25116
rect 4060 24836 4116 24846
rect 4060 24742 4116 24780
rect 3500 24670 3502 24722
rect 3554 24670 3556 24722
rect 3276 23774 3278 23826
rect 3330 23774 3332 23826
rect 3276 23762 3332 23774
rect 3388 23828 3444 23838
rect 3388 23734 3444 23772
rect 3388 23044 3444 23054
rect 3276 22372 3332 22382
rect 3388 22372 3444 22988
rect 3276 22370 3444 22372
rect 3276 22318 3278 22370
rect 3330 22318 3444 22370
rect 3276 22316 3444 22318
rect 3500 22372 3556 24670
rect 3948 24724 4004 24734
rect 3948 24630 4004 24668
rect 4060 24500 4116 24510
rect 4060 24406 4116 24444
rect 4060 23940 4116 23950
rect 4172 23940 4228 26236
rect 4508 26226 4564 26236
rect 4060 23938 4228 23940
rect 4060 23886 4062 23938
rect 4114 23886 4228 23938
rect 4060 23884 4228 23886
rect 4284 26068 4340 26078
rect 4060 23874 4116 23884
rect 3724 23714 3780 23726
rect 3724 23662 3726 23714
rect 3778 23662 3780 23714
rect 3724 23044 3780 23662
rect 3724 22978 3780 22988
rect 3948 23714 4004 23726
rect 3948 23662 3950 23714
rect 4002 23662 4004 23714
rect 3948 23044 4004 23662
rect 3948 22978 4004 22988
rect 3500 22370 4228 22372
rect 3500 22318 3502 22370
rect 3554 22318 4228 22370
rect 3500 22316 4228 22318
rect 3276 22306 3332 22316
rect 3500 22306 3556 22316
rect 4172 22258 4228 22316
rect 4172 22206 4174 22258
rect 4226 22206 4228 22258
rect 4172 22194 4228 22206
rect 3164 21758 3166 21810
rect 3218 21758 3220 21810
rect 3164 21476 3220 21758
rect 4172 21586 4228 21598
rect 4172 21534 4174 21586
rect 4226 21534 4228 21586
rect 3164 21410 3220 21420
rect 4060 21474 4116 21486
rect 4060 21422 4062 21474
rect 4114 21422 4116 21474
rect 3836 21364 3892 21374
rect 3836 21270 3892 21308
rect 2604 21084 2772 21140
rect 2492 20692 2548 20702
rect 2492 20598 2548 20636
rect 2716 20020 2772 21084
rect 2828 21074 2884 21084
rect 3164 21140 3220 21150
rect 3164 20130 3220 21084
rect 3276 20692 3332 20702
rect 3276 20242 3332 20636
rect 3276 20190 3278 20242
rect 3330 20190 3332 20242
rect 3276 20178 3332 20190
rect 3724 20244 3780 20254
rect 3164 20078 3166 20130
rect 3218 20078 3220 20130
rect 3164 20066 3220 20078
rect 3388 20132 3444 20142
rect 2716 19964 2884 20020
rect 2604 19908 2660 19918
rect 2604 19814 2660 19852
rect 2716 19794 2772 19806
rect 2716 19742 2718 19794
rect 2770 19742 2772 19794
rect 2716 19348 2772 19742
rect 2716 19282 2772 19292
rect 2492 19122 2548 19134
rect 2492 19070 2494 19122
rect 2546 19070 2548 19122
rect 2492 18676 2548 19070
rect 2492 18610 2548 18620
rect 2828 18450 2884 19964
rect 3052 18676 3108 18686
rect 3388 18676 3444 20076
rect 3500 20018 3556 20030
rect 3500 19966 3502 20018
rect 3554 19966 3556 20018
rect 3500 19348 3556 19966
rect 3724 20018 3780 20188
rect 3724 19966 3726 20018
rect 3778 19966 3780 20018
rect 3724 19954 3780 19966
rect 3724 19796 3780 19806
rect 3724 19702 3780 19740
rect 4060 19796 4116 21422
rect 4172 20916 4228 21534
rect 4172 20850 4228 20860
rect 4060 19730 4116 19740
rect 3612 19348 3668 19358
rect 3500 19292 3612 19348
rect 3612 19124 3668 19292
rect 3052 18674 3444 18676
rect 3052 18622 3054 18674
rect 3106 18622 3444 18674
rect 3052 18620 3444 18622
rect 3052 18610 3108 18620
rect 3388 18562 3444 18620
rect 3500 18676 3556 18686
rect 3500 18582 3556 18620
rect 3388 18510 3390 18562
rect 3442 18510 3444 18562
rect 3388 18498 3444 18510
rect 3612 18562 3668 19068
rect 4284 18900 4340 26012
rect 4620 26068 4676 26078
rect 4620 25974 4676 26012
rect 4620 24834 4676 24846
rect 4620 24782 4622 24834
rect 4674 24782 4676 24834
rect 4396 24724 4452 24734
rect 4508 24724 4564 24734
rect 4452 24722 4564 24724
rect 4452 24670 4510 24722
rect 4562 24670 4564 24722
rect 4452 24668 4564 24670
rect 4396 23826 4452 24668
rect 4508 24658 4564 24668
rect 4620 24052 4676 24782
rect 4620 23986 4676 23996
rect 4732 23940 4788 27582
rect 5068 26908 5124 27916
rect 5180 27746 5236 27758
rect 5180 27694 5182 27746
rect 5234 27694 5236 27746
rect 5180 27634 5236 27694
rect 5180 27582 5182 27634
rect 5234 27582 5236 27634
rect 5180 27570 5236 27582
rect 5292 27076 5348 28364
rect 5292 27010 5348 27020
rect 5068 26852 5460 26908
rect 4956 26292 5012 26302
rect 4844 25620 4900 25630
rect 4844 25526 4900 25564
rect 4844 24948 4900 24958
rect 4956 24948 5012 26236
rect 4844 24946 5012 24948
rect 4844 24894 4846 24946
rect 4898 24894 5012 24946
rect 4844 24892 5012 24894
rect 4844 24882 4900 24892
rect 4732 23884 4900 23940
rect 4396 23774 4398 23826
rect 4450 23774 4452 23826
rect 4396 20132 4452 23774
rect 4508 23716 4564 23726
rect 4508 23622 4564 23660
rect 4732 23714 4788 23726
rect 4732 23662 4734 23714
rect 4786 23662 4788 23714
rect 4620 23044 4676 23054
rect 4620 22596 4676 22988
rect 4620 22530 4676 22540
rect 4508 22372 4564 22382
rect 4508 22278 4564 22316
rect 4732 22260 4788 23662
rect 4732 22194 4788 22204
rect 4844 22036 4900 23884
rect 4732 21980 4900 22036
rect 5180 23154 5236 23166
rect 5180 23102 5182 23154
rect 5234 23102 5236 23154
rect 4620 21588 4676 21598
rect 4620 21494 4676 21532
rect 4732 21252 4788 21980
rect 4844 21812 4900 21822
rect 5180 21812 5236 23102
rect 4900 21756 5236 21812
rect 4844 21718 4900 21756
rect 4732 21186 4788 21196
rect 4620 20916 4676 20926
rect 4620 20822 4676 20860
rect 5292 20916 5348 20926
rect 5068 20578 5124 20590
rect 5068 20526 5070 20578
rect 5122 20526 5124 20578
rect 4396 20066 4452 20076
rect 4508 20468 4564 20478
rect 4284 18834 4340 18844
rect 4508 18676 4564 20412
rect 3612 18510 3614 18562
rect 3666 18510 3668 18562
rect 3612 18498 3668 18510
rect 3836 18674 4564 18676
rect 3836 18622 4510 18674
rect 4562 18622 4564 18674
rect 3836 18620 4564 18622
rect 2828 18398 2830 18450
rect 2882 18398 2884 18450
rect 2828 18004 2884 18398
rect 2828 17938 2884 17948
rect 3500 18004 3556 18014
rect 2380 17502 2382 17554
rect 2434 17502 2436 17554
rect 2044 17490 2100 17500
rect 2380 17490 2436 17502
rect 2604 17666 2660 17678
rect 2604 17614 2606 17666
rect 2658 17614 2660 17666
rect 2604 17444 2660 17614
rect 3500 17556 3556 17948
rect 3500 17490 3556 17500
rect 3164 17444 3220 17454
rect 2604 17442 3220 17444
rect 2604 17390 3166 17442
rect 3218 17390 3220 17442
rect 2604 17388 3220 17390
rect 2044 17332 2100 17342
rect 2044 17106 2100 17276
rect 2044 17054 2046 17106
rect 2098 17054 2100 17106
rect 2044 17042 2100 17054
rect 2604 17108 2660 17388
rect 3164 17378 3220 17388
rect 3724 17444 3780 17454
rect 3724 17350 3780 17388
rect 3836 17220 3892 18620
rect 4508 18610 4564 18620
rect 4620 20130 4676 20142
rect 4620 20078 4622 20130
rect 4674 20078 4676 20130
rect 4620 19346 4676 20078
rect 4956 20132 5012 20142
rect 4956 20038 5012 20076
rect 5068 20020 5124 20526
rect 5068 19954 5124 19964
rect 5180 20244 5236 20254
rect 4620 19294 4622 19346
rect 4674 19294 4676 19346
rect 4172 18450 4228 18462
rect 4172 18398 4174 18450
rect 4226 18398 4228 18450
rect 3948 18226 4004 18238
rect 3948 18174 3950 18226
rect 4002 18174 4004 18226
rect 3948 17780 4004 18174
rect 4060 17780 4116 17790
rect 3948 17778 4116 17780
rect 3948 17726 4062 17778
rect 4114 17726 4116 17778
rect 3948 17724 4116 17726
rect 4060 17714 4116 17724
rect 3948 17556 4004 17566
rect 3948 17462 4004 17500
rect 4172 17444 4228 18398
rect 4284 17668 4340 17678
rect 4620 17668 4676 19294
rect 5068 19012 5124 19022
rect 5180 19012 5236 20188
rect 5292 20018 5348 20860
rect 5292 19966 5294 20018
rect 5346 19966 5348 20018
rect 5292 19954 5348 19966
rect 5068 19010 5236 19012
rect 5068 18958 5070 19010
rect 5122 18958 5236 19010
rect 5068 18956 5236 18958
rect 5068 18946 5124 18956
rect 5180 18562 5236 18956
rect 5180 18510 5182 18562
rect 5234 18510 5236 18562
rect 4844 18452 4900 18462
rect 4844 18358 4900 18396
rect 5180 18116 5236 18510
rect 5180 18050 5236 18060
rect 4284 17666 4676 17668
rect 4284 17614 4286 17666
rect 4338 17614 4676 17666
rect 4284 17612 4676 17614
rect 4284 17602 4340 17612
rect 4956 17554 5012 17566
rect 4956 17502 4958 17554
rect 5010 17502 5012 17554
rect 4620 17444 4676 17454
rect 4172 17378 4228 17388
rect 4284 17442 4676 17444
rect 4284 17390 4622 17442
rect 4674 17390 4676 17442
rect 4284 17388 4676 17390
rect 2604 17042 2660 17052
rect 3724 17164 3892 17220
rect 2380 16994 2436 17006
rect 2380 16942 2382 16994
rect 2434 16942 2436 16994
rect 1484 14242 1540 14252
rect 1708 15314 1988 15316
rect 1708 15262 1822 15314
rect 1874 15262 1988 15314
rect 1708 15260 1988 15262
rect 2156 16772 2212 16782
rect 1708 12852 1764 15260
rect 1820 15250 1876 15260
rect 1820 15092 1876 15102
rect 1820 14530 1876 15036
rect 1820 14478 1822 14530
rect 1874 14478 1876 14530
rect 1820 14466 1876 14478
rect 2044 14308 2100 14318
rect 2044 14214 2100 14252
rect 2044 13972 2100 13982
rect 2044 13746 2100 13916
rect 2156 13860 2212 16716
rect 2380 16212 2436 16942
rect 2716 16996 2772 17006
rect 2716 16902 2772 16940
rect 3052 16884 3108 16894
rect 3052 16790 3108 16828
rect 3724 16772 3780 17164
rect 4284 17108 4340 17388
rect 4620 17378 4676 17388
rect 3836 17052 4340 17108
rect 3836 16994 3892 17052
rect 3836 16942 3838 16994
rect 3890 16942 3892 16994
rect 3836 16930 3892 16942
rect 3724 16716 3892 16772
rect 2492 16212 2548 16222
rect 2380 16210 2548 16212
rect 2380 16158 2494 16210
rect 2546 16158 2548 16210
rect 2380 16156 2548 16158
rect 2492 16146 2548 16156
rect 2492 15202 2548 15214
rect 2492 15150 2494 15202
rect 2546 15150 2548 15202
rect 2492 15148 2548 15150
rect 2492 15092 3220 15148
rect 2380 14980 2436 14990
rect 2380 14420 2436 14924
rect 3164 14642 3220 15092
rect 3164 14590 3166 14642
rect 3218 14590 3220 14642
rect 3164 14578 3220 14590
rect 3500 14644 3556 14654
rect 3500 14550 3556 14588
rect 3388 14532 3444 14542
rect 3388 14438 3444 14476
rect 3836 14532 3892 16716
rect 4956 16324 5012 17502
rect 4956 16258 5012 16268
rect 4620 16210 4676 16222
rect 4620 16158 4622 16210
rect 4674 16158 4676 16210
rect 4620 16100 4676 16158
rect 4620 16034 4676 16044
rect 5068 15988 5124 15998
rect 5068 15894 5124 15932
rect 4956 15428 5012 15438
rect 4620 15204 4676 15214
rect 4956 15204 5012 15372
rect 4620 15202 5012 15204
rect 4620 15150 4622 15202
rect 4674 15150 5012 15202
rect 4620 15148 5012 15150
rect 4620 15138 4676 15148
rect 3948 14812 4228 14868
rect 3948 14756 4004 14812
rect 3948 14690 4004 14700
rect 4172 14754 4228 14812
rect 4172 14702 4174 14754
rect 4226 14702 4228 14754
rect 4172 14690 4228 14702
rect 4508 14756 4564 14766
rect 4060 14644 4116 14654
rect 4060 14532 4116 14588
rect 4172 14532 4228 14542
rect 3836 14530 4004 14532
rect 3836 14478 3838 14530
rect 3890 14478 4004 14530
rect 3836 14476 4004 14478
rect 3836 14466 3892 14476
rect 2156 13794 2212 13804
rect 2268 14418 2436 14420
rect 2268 14366 2382 14418
rect 2434 14366 2436 14418
rect 2268 14364 2436 14366
rect 2044 13694 2046 13746
rect 2098 13694 2100 13746
rect 2044 13682 2100 13694
rect 2268 13748 2324 14364
rect 2380 14354 2436 14364
rect 2716 14420 2772 14430
rect 3052 14420 3108 14430
rect 2716 14326 2772 14364
rect 2828 14418 3108 14420
rect 2828 14366 3054 14418
rect 3106 14366 3108 14418
rect 2828 14364 3108 14366
rect 2380 13860 2436 13870
rect 2716 13860 2772 13870
rect 2380 13858 2716 13860
rect 2380 13806 2382 13858
rect 2434 13806 2716 13858
rect 2380 13804 2716 13806
rect 2380 13794 2436 13804
rect 2716 13766 2772 13804
rect 2268 13682 2324 13692
rect 2156 13634 2212 13646
rect 2156 13582 2158 13634
rect 2210 13582 2212 13634
rect 1260 12786 1316 12796
rect 1596 12796 1764 12852
rect 2044 12850 2100 12862
rect 2044 12798 2046 12850
rect 2098 12798 2100 12850
rect 1036 10770 1092 10780
rect 1596 10500 1652 12796
rect 1708 12628 1764 12638
rect 1708 10724 1764 12572
rect 1932 12180 1988 12190
rect 1708 10630 1764 10668
rect 1820 12178 1988 12180
rect 1820 12126 1934 12178
rect 1986 12126 1988 12178
rect 1820 12124 1988 12126
rect 1596 10444 1764 10500
rect 1708 9268 1764 10444
rect 1820 10052 1876 12124
rect 1932 12114 1988 12124
rect 2044 11844 2100 12798
rect 1932 11788 2100 11844
rect 1932 11732 1988 11788
rect 1932 11666 1988 11676
rect 2044 11620 2100 11630
rect 2156 11620 2212 13582
rect 2828 12964 2884 14364
rect 3052 14354 3108 14364
rect 3836 14308 3892 14318
rect 3724 14252 3836 14308
rect 3500 13972 3556 13982
rect 2492 12908 2884 12964
rect 2940 13858 2996 13870
rect 2940 13806 2942 13858
rect 2994 13806 2996 13858
rect 2940 13748 2996 13806
rect 2380 12852 2436 12862
rect 2380 12758 2436 12796
rect 2044 11618 2212 11620
rect 2044 11566 2046 11618
rect 2098 11566 2212 11618
rect 2044 11564 2212 11566
rect 2044 11554 2100 11564
rect 1932 11508 1988 11518
rect 1932 11394 1988 11452
rect 1932 11342 1934 11394
rect 1986 11342 1988 11394
rect 1932 11330 1988 11342
rect 2156 11396 2212 11406
rect 2044 10836 2100 10846
rect 2044 10742 2100 10780
rect 2156 10276 2212 11340
rect 2492 11396 2548 12908
rect 2716 12740 2772 12750
rect 2492 11302 2548 11340
rect 2604 12738 2772 12740
rect 2604 12686 2718 12738
rect 2770 12686 2772 12738
rect 2604 12684 2772 12686
rect 2156 10210 2212 10220
rect 2268 11282 2324 11294
rect 2268 11230 2270 11282
rect 2322 11230 2324 11282
rect 1820 9826 1876 9996
rect 1820 9774 1822 9826
rect 1874 9774 1876 9826
rect 1820 9762 1876 9774
rect 1820 9268 1876 9278
rect 1708 9266 1876 9268
rect 1708 9214 1822 9266
rect 1874 9214 1876 9266
rect 1708 9212 1876 9214
rect 1708 6132 1764 9212
rect 1820 9156 1876 9212
rect 2156 9268 2212 9278
rect 2156 9174 2212 9212
rect 1820 9090 1876 9100
rect 1820 8258 1876 8270
rect 1820 8206 1822 8258
rect 1874 8206 1876 8258
rect 1820 6692 1876 8206
rect 2268 7924 2324 11230
rect 2380 11170 2436 11182
rect 2380 11118 2382 11170
rect 2434 11118 2436 11170
rect 2380 9940 2436 11118
rect 2492 10610 2548 10622
rect 2492 10558 2494 10610
rect 2546 10558 2548 10610
rect 2492 10164 2548 10558
rect 2492 10098 2548 10108
rect 2492 9940 2548 9950
rect 2380 9938 2548 9940
rect 2380 9886 2494 9938
rect 2546 9886 2548 9938
rect 2380 9884 2548 9886
rect 2492 9874 2548 9884
rect 2604 9828 2660 12684
rect 2716 12674 2772 12684
rect 2716 12066 2772 12078
rect 2716 12014 2718 12066
rect 2770 12014 2772 12066
rect 2716 11172 2772 12014
rect 2828 11172 2884 11182
rect 2716 11170 2884 11172
rect 2716 11118 2830 11170
rect 2882 11118 2884 11170
rect 2716 11116 2884 11118
rect 2828 11106 2884 11116
rect 2604 9772 2884 9828
rect 2268 7858 2324 7868
rect 2380 9716 2436 9726
rect 2268 7700 2324 7710
rect 2268 7606 2324 7644
rect 1932 6692 1988 6702
rect 1820 6690 2100 6692
rect 1820 6638 1934 6690
rect 1986 6638 2100 6690
rect 1820 6636 2100 6638
rect 1932 6626 1988 6636
rect 1932 6132 1988 6142
rect 1708 6076 1932 6132
rect 1932 6038 1988 6076
rect 2044 5236 2100 6636
rect 2380 6132 2436 9660
rect 2716 9380 2772 9390
rect 2716 9156 2772 9324
rect 2716 9062 2772 9100
rect 2828 8260 2884 9772
rect 2940 9716 2996 13692
rect 3052 13522 3108 13534
rect 3388 13524 3444 13534
rect 3052 13470 3054 13522
rect 3106 13470 3108 13522
rect 3052 12964 3108 13470
rect 3052 12898 3108 12908
rect 3164 13522 3444 13524
rect 3164 13470 3390 13522
rect 3442 13470 3444 13522
rect 3164 13468 3444 13470
rect 3052 12740 3108 12750
rect 3052 12646 3108 12684
rect 3164 11618 3220 13468
rect 3388 13458 3444 13468
rect 3500 13188 3556 13916
rect 3724 13860 3780 14252
rect 3836 14242 3892 14252
rect 3724 13766 3780 13804
rect 3948 13634 4004 14476
rect 3948 13582 3950 13634
rect 4002 13582 4004 13634
rect 3948 13570 4004 13582
rect 4060 14530 4228 14532
rect 4060 14478 4174 14530
rect 4226 14478 4228 14530
rect 4060 14476 4228 14478
rect 3388 13132 3556 13188
rect 3388 11788 3444 13132
rect 3500 12962 3556 12974
rect 3500 12910 3502 12962
rect 3554 12910 3556 12962
rect 3500 12852 3556 12910
rect 3500 12786 3556 12796
rect 3724 12852 3780 12862
rect 3724 12292 3780 12796
rect 3724 12226 3780 12236
rect 3388 11732 3556 11788
rect 4060 11732 4116 14476
rect 4172 14466 4228 14476
rect 4396 14532 4452 14542
rect 4172 13636 4228 13646
rect 4172 13634 4340 13636
rect 4172 13582 4174 13634
rect 4226 13582 4340 13634
rect 4172 13580 4340 13582
rect 4172 13570 4228 13580
rect 3164 11566 3166 11618
rect 3218 11566 3220 11618
rect 3164 11554 3220 11566
rect 3052 11508 3108 11518
rect 3052 11394 3108 11452
rect 3052 11342 3054 11394
rect 3106 11342 3108 11394
rect 3052 11330 3108 11342
rect 3388 11396 3444 11406
rect 3388 11302 3444 11340
rect 3276 11172 3332 11182
rect 3276 10722 3332 11116
rect 3276 10670 3278 10722
rect 3330 10670 3332 10722
rect 3276 10658 3332 10670
rect 3388 10724 3444 10734
rect 2940 9650 2996 9660
rect 3052 10052 3108 10062
rect 3052 9266 3108 9996
rect 3052 9214 3054 9266
rect 3106 9214 3108 9266
rect 3052 9156 3108 9214
rect 3052 9090 3108 9100
rect 2604 8204 2884 8260
rect 2492 8146 2548 8158
rect 2492 8094 2494 8146
rect 2546 8094 2548 8146
rect 2492 7698 2548 8094
rect 2492 7646 2494 7698
rect 2546 7646 2548 7698
rect 2492 7634 2548 7646
rect 2604 7140 2660 8204
rect 2828 8036 2884 8046
rect 2828 7586 2884 7980
rect 3276 7924 3332 7934
rect 3164 7588 3220 7598
rect 2828 7534 2830 7586
rect 2882 7534 2884 7586
rect 2828 7522 2884 7534
rect 2940 7586 3220 7588
rect 2940 7534 3166 7586
rect 3218 7534 3220 7586
rect 2940 7532 3220 7534
rect 2492 7084 2660 7140
rect 2492 6580 2548 7084
rect 2940 7028 2996 7532
rect 3164 7522 3220 7532
rect 2604 6972 2996 7028
rect 2604 6802 2660 6972
rect 2604 6750 2606 6802
rect 2658 6750 2660 6802
rect 2604 6738 2660 6750
rect 2492 6524 2996 6580
rect 2492 6132 2548 6142
rect 2380 6130 2548 6132
rect 2380 6078 2494 6130
rect 2546 6078 2548 6130
rect 2380 6076 2548 6078
rect 2492 6066 2548 6076
rect 2044 5170 2100 5180
rect 2716 3442 2772 3454
rect 2716 3390 2718 3442
rect 2770 3390 2772 3442
rect 2716 3220 2772 3390
rect 2940 3442 2996 6524
rect 3276 6018 3332 7868
rect 3388 7252 3444 10668
rect 3500 7700 3556 11732
rect 3836 11676 4116 11732
rect 4172 12852 4228 12862
rect 3612 11620 3668 11630
rect 3612 11394 3668 11564
rect 3612 11342 3614 11394
rect 3666 11342 3668 11394
rect 3612 11284 3668 11342
rect 3612 11218 3668 11228
rect 3724 9268 3780 9278
rect 3836 9268 3892 11676
rect 4172 11618 4228 12796
rect 4172 11566 4174 11618
rect 4226 11566 4228 11618
rect 4172 11554 4228 11566
rect 4060 11508 4116 11518
rect 4060 11394 4116 11452
rect 4060 11342 4062 11394
rect 4114 11342 4116 11394
rect 4060 11330 4116 11342
rect 3948 11172 4004 11182
rect 3948 11078 4004 11116
rect 4284 10052 4340 13580
rect 4396 12962 4452 14476
rect 4508 14308 4564 14700
rect 4956 14642 5012 15148
rect 5180 15204 5236 15242
rect 5180 15138 5236 15148
rect 4956 14590 4958 14642
rect 5010 14590 5012 14642
rect 4956 14578 5012 14590
rect 4844 14532 4900 14542
rect 4844 14438 4900 14476
rect 4508 14242 4564 14252
rect 4956 14420 5012 14430
rect 4508 14084 4564 14094
rect 4564 14028 4676 14084
rect 4508 14018 4564 14028
rect 4396 12910 4398 12962
rect 4450 12910 4452 12962
rect 4396 12898 4452 12910
rect 4508 11284 4564 11294
rect 4508 11190 4564 11228
rect 4620 10612 4676 14028
rect 4732 13746 4788 13758
rect 4732 13694 4734 13746
rect 4786 13694 4788 13746
rect 4732 12404 4788 13694
rect 4844 13412 4900 13422
rect 4844 12962 4900 13356
rect 4956 13076 5012 14364
rect 5292 13636 5348 13646
rect 5068 13076 5124 13086
rect 4956 13074 5124 13076
rect 4956 13022 5070 13074
rect 5122 13022 5124 13074
rect 4956 13020 5124 13022
rect 5068 13010 5124 13020
rect 4844 12910 4846 12962
rect 4898 12910 4900 12962
rect 4844 12898 4900 12910
rect 4732 12338 4788 12348
rect 4844 12740 4900 12750
rect 4844 12180 4900 12684
rect 5180 12292 5236 12302
rect 5180 12198 5236 12236
rect 4732 12124 4900 12180
rect 4732 11844 4788 12124
rect 5180 12068 5236 12078
rect 4844 12039 5180 12068
rect 4844 11987 4846 12039
rect 4898 12012 5180 12039
rect 4898 11987 4900 12012
rect 5180 12002 5236 12012
rect 4844 11975 4900 11987
rect 5068 11844 5124 11854
rect 4732 11788 4900 11844
rect 4732 11620 4788 11630
rect 4732 11394 4788 11564
rect 4844 11508 4900 11788
rect 4844 11452 5012 11508
rect 4732 11342 4734 11394
rect 4786 11342 4788 11394
rect 4732 11330 4788 11342
rect 3724 9266 3892 9268
rect 3724 9214 3726 9266
rect 3778 9214 3892 9266
rect 3724 9212 3892 9214
rect 4060 9996 4340 10052
rect 4060 9266 4116 9996
rect 4284 9940 4340 9996
rect 4284 9874 4340 9884
rect 4508 10556 4676 10612
rect 4060 9214 4062 9266
rect 4114 9214 4116 9266
rect 3724 9202 3780 9212
rect 4060 9202 4116 9214
rect 3500 7634 3556 7644
rect 3836 7924 3892 7934
rect 3836 7698 3892 7868
rect 3836 7646 3838 7698
rect 3890 7646 3892 7698
rect 3836 7634 3892 7646
rect 4508 7698 4564 10556
rect 4620 9938 4676 9950
rect 4620 9886 4622 9938
rect 4674 9886 4676 9938
rect 4620 9716 4676 9886
rect 4620 9650 4676 9660
rect 4844 9380 4900 9390
rect 4844 9266 4900 9324
rect 4844 9214 4846 9266
rect 4898 9214 4900 9266
rect 4844 9202 4900 9214
rect 4620 9044 4676 9054
rect 4956 9044 5012 11452
rect 5068 9268 5124 11788
rect 5180 9940 5236 9950
rect 5292 9940 5348 13580
rect 5404 11060 5460 26852
rect 5516 20244 5572 28364
rect 6636 28420 6692 28812
rect 6748 28644 6804 28654
rect 6748 28550 6804 28588
rect 6636 28364 6804 28420
rect 5628 27076 5684 27086
rect 5628 26982 5684 27020
rect 5740 24724 5796 24734
rect 5740 24630 5796 24668
rect 5628 21812 5684 21822
rect 5628 20802 5684 21756
rect 5628 20750 5630 20802
rect 5682 20750 5684 20802
rect 5628 20738 5684 20750
rect 5516 20178 5572 20188
rect 5628 20132 5684 20142
rect 5852 20132 5908 28364
rect 6748 27860 6804 28364
rect 6860 28084 6916 30604
rect 6972 30434 7028 30716
rect 6972 30382 6974 30434
rect 7026 30382 7028 30434
rect 6972 30370 7028 30382
rect 7084 30716 7252 30772
rect 7084 29652 7140 30716
rect 7308 30434 7364 30446
rect 7308 30382 7310 30434
rect 7362 30382 7364 30434
rect 7196 29986 7252 29998
rect 7196 29934 7198 29986
rect 7250 29934 7252 29986
rect 7196 29876 7252 29934
rect 7308 29988 7364 30382
rect 7532 30212 7588 30222
rect 7756 30212 7812 32956
rect 7980 32674 8036 32686
rect 7980 32622 7982 32674
rect 8034 32622 8036 32674
rect 7980 31948 8036 32622
rect 8316 32676 8372 32686
rect 8316 32582 8372 32620
rect 8540 32562 8596 33292
rect 8876 32786 8932 33516
rect 9324 33460 9380 33470
rect 8876 32734 8878 32786
rect 8930 32734 8932 32786
rect 8876 32722 8932 32734
rect 9212 32900 9268 32910
rect 8540 32510 8542 32562
rect 8594 32510 8596 32562
rect 8540 32498 8596 32510
rect 9212 32340 9268 32844
rect 8365 32172 8629 32182
rect 8421 32116 8469 32172
rect 8525 32116 8573 32172
rect 8365 32106 8629 32116
rect 7980 31892 8372 31948
rect 8316 31668 8372 31892
rect 8316 31574 8372 31612
rect 8428 31780 8484 31790
rect 8092 31556 8148 31566
rect 7532 30210 7812 30212
rect 7532 30158 7534 30210
rect 7586 30158 7812 30210
rect 7532 30156 7812 30158
rect 7868 31554 8148 31556
rect 7868 31502 8094 31554
rect 8146 31502 8148 31554
rect 7868 31500 8148 31502
rect 7868 30210 7924 31500
rect 8092 31490 8148 31500
rect 7868 30158 7870 30210
rect 7922 30158 7924 30210
rect 7532 30146 7588 30156
rect 7868 30146 7924 30158
rect 7980 31220 8036 31230
rect 7644 29988 7700 29998
rect 7308 29986 7700 29988
rect 7308 29934 7646 29986
rect 7698 29934 7700 29986
rect 7308 29932 7700 29934
rect 7644 29922 7700 29932
rect 7196 29810 7252 29820
rect 7084 29596 7924 29652
rect 7756 29316 7812 29326
rect 7644 29260 7756 29316
rect 7644 28756 7700 29260
rect 7756 29250 7812 29260
rect 6972 28700 7700 28756
rect 6972 28530 7028 28700
rect 6972 28478 6974 28530
rect 7026 28478 7028 28530
rect 6972 28466 7028 28478
rect 7084 28532 7140 28542
rect 7084 28530 7476 28532
rect 7084 28478 7086 28530
rect 7138 28478 7476 28530
rect 7084 28476 7476 28478
rect 7084 28466 7140 28476
rect 6860 28028 7252 28084
rect 7084 27860 7140 27870
rect 6748 27858 7140 27860
rect 6748 27806 7086 27858
rect 7138 27806 7140 27858
rect 6748 27804 7140 27806
rect 6412 26962 6468 26974
rect 6412 26910 6414 26962
rect 6466 26910 6468 26962
rect 6412 26514 6468 26910
rect 6972 26908 7028 27804
rect 7084 27794 7140 27804
rect 7196 27636 7252 28028
rect 7420 28082 7476 28476
rect 7644 28530 7700 28700
rect 7644 28478 7646 28530
rect 7698 28478 7700 28530
rect 7644 28466 7700 28478
rect 7868 28532 7924 29596
rect 7980 28756 8036 31164
rect 8428 30772 8484 31724
rect 8988 31668 9044 31678
rect 8204 30716 8484 30772
rect 8876 31556 8932 31566
rect 8092 30324 8148 30334
rect 8204 30324 8260 30716
rect 8365 30604 8629 30614
rect 8421 30548 8469 30604
rect 8525 30548 8573 30604
rect 8365 30538 8629 30548
rect 8148 30268 8260 30324
rect 8092 30258 8148 30268
rect 8092 30098 8148 30110
rect 8092 30046 8094 30098
rect 8146 30046 8148 30098
rect 8092 29540 8148 30046
rect 8540 29986 8596 29998
rect 8540 29934 8542 29986
rect 8594 29934 8596 29986
rect 8540 29652 8596 29934
rect 8540 29586 8596 29596
rect 8092 29484 8372 29540
rect 8204 29316 8260 29326
rect 8204 29222 8260 29260
rect 8316 29204 8372 29484
rect 8316 29138 8372 29148
rect 8365 29036 8629 29046
rect 8421 28980 8469 29036
rect 8525 28980 8573 29036
rect 8365 28970 8629 28980
rect 8316 28868 8372 28878
rect 8316 28774 8372 28812
rect 8652 28868 8708 28878
rect 8652 28774 8708 28812
rect 7980 28700 8260 28756
rect 7980 28532 8036 28542
rect 7868 28530 8036 28532
rect 7868 28478 7982 28530
rect 8034 28478 8036 28530
rect 7868 28476 8036 28478
rect 7420 28030 7422 28082
rect 7474 28030 7476 28082
rect 6748 26852 7028 26908
rect 7084 27580 7252 27636
rect 7308 27972 7364 27982
rect 6748 26516 6804 26852
rect 6412 26462 6414 26514
rect 6466 26462 6468 26514
rect 6412 26450 6468 26462
rect 6636 26460 6804 26516
rect 6076 26292 6132 26302
rect 6076 26198 6132 26236
rect 6524 26292 6580 26302
rect 6524 26198 6580 26236
rect 6636 26068 6692 26460
rect 6748 26290 6804 26302
rect 6748 26238 6750 26290
rect 6802 26238 6804 26290
rect 6748 26180 6804 26238
rect 6748 26124 7028 26180
rect 6636 26012 6804 26068
rect 6188 25732 6244 25742
rect 5964 23042 6020 23054
rect 5964 22990 5966 23042
rect 6018 22990 6020 23042
rect 5964 22484 6020 22990
rect 6076 22484 6132 22494
rect 5964 22482 6132 22484
rect 5964 22430 6078 22482
rect 6130 22430 6132 22482
rect 5964 22428 6132 22430
rect 6076 22418 6132 22428
rect 5964 22260 6020 22270
rect 5964 22166 6020 22204
rect 6188 22148 6244 25676
rect 6524 24610 6580 24622
rect 6524 24558 6526 24610
rect 6578 24558 6580 24610
rect 6412 24500 6468 24510
rect 6300 24164 6356 24174
rect 6300 22370 6356 24108
rect 6412 23938 6468 24444
rect 6524 24052 6580 24558
rect 6636 24052 6692 24062
rect 6524 24050 6692 24052
rect 6524 23998 6638 24050
rect 6690 23998 6692 24050
rect 6524 23996 6692 23998
rect 6636 23986 6692 23996
rect 6412 23886 6414 23938
rect 6466 23886 6468 23938
rect 6412 23874 6468 23886
rect 6748 22932 6804 26012
rect 6972 24052 7028 26124
rect 7084 24164 7140 27580
rect 7196 26628 7252 26638
rect 7196 26514 7252 26572
rect 7196 26462 7198 26514
rect 7250 26462 7252 26514
rect 7196 26450 7252 26462
rect 7084 24108 7252 24164
rect 6972 23996 7140 24052
rect 6860 23938 6916 23950
rect 6860 23886 6862 23938
rect 6914 23886 6916 23938
rect 6860 23828 6916 23886
rect 6972 23828 7028 23838
rect 6860 23772 6972 23828
rect 6972 23762 7028 23772
rect 7084 23826 7140 23996
rect 7084 23774 7086 23826
rect 7138 23774 7140 23826
rect 6748 22866 6804 22876
rect 7084 22484 7140 23774
rect 6300 22318 6302 22370
rect 6354 22318 6356 22370
rect 6300 22306 6356 22318
rect 6972 22428 7140 22484
rect 7196 22484 7252 24108
rect 7308 23828 7364 27916
rect 7420 26516 7476 28030
rect 7980 27970 8036 28476
rect 7980 27918 7982 27970
rect 8034 27918 8036 27970
rect 7980 27906 8036 27918
rect 8092 27860 8148 27870
rect 8092 26908 8148 27804
rect 7420 23940 7476 26460
rect 7980 26852 8148 26908
rect 7532 26404 7588 26414
rect 7532 26290 7588 26348
rect 7532 26238 7534 26290
rect 7586 26238 7588 26290
rect 7532 26226 7588 26238
rect 7980 26290 8036 26852
rect 7980 26238 7982 26290
rect 8034 26238 8036 26290
rect 7644 25394 7700 25406
rect 7644 25342 7646 25394
rect 7698 25342 7700 25394
rect 7644 24612 7700 25342
rect 7644 24546 7700 24556
rect 7980 25394 8036 26238
rect 8204 26180 8260 28700
rect 8428 27860 8484 27870
rect 8428 27766 8484 27804
rect 8365 27468 8629 27478
rect 8421 27412 8469 27468
rect 8525 27412 8573 27468
rect 8365 27402 8629 27412
rect 8876 27300 8932 31500
rect 8988 30882 9044 31612
rect 8988 30830 8990 30882
rect 9042 30830 9044 30882
rect 8988 30818 9044 30830
rect 9212 31666 9268 32284
rect 9212 31614 9214 31666
rect 9266 31614 9268 31666
rect 9212 31444 9268 31614
rect 9324 32452 9380 33404
rect 9996 33460 10052 34636
rect 10220 34132 10276 34142
rect 10220 34038 10276 34076
rect 9996 33394 10052 33404
rect 10668 34018 10724 34030
rect 10668 33966 10670 34018
rect 10722 33966 10724 34018
rect 10332 33234 10388 33246
rect 10332 33182 10334 33234
rect 10386 33182 10388 33234
rect 9660 32788 9716 32798
rect 9660 32694 9716 32732
rect 10332 32788 10388 33182
rect 10668 32900 10724 33966
rect 11116 34020 11172 34030
rect 11116 33926 11172 33964
rect 10668 32834 10724 32844
rect 11116 33346 11172 33358
rect 11116 33294 11118 33346
rect 11170 33294 11172 33346
rect 10332 32722 10388 32732
rect 10780 32674 10836 32686
rect 10780 32622 10782 32674
rect 10834 32622 10836 32674
rect 9436 32564 9492 32574
rect 9436 32470 9492 32508
rect 9772 32562 9828 32574
rect 9772 32510 9774 32562
rect 9826 32510 9828 32562
rect 9324 31666 9380 32396
rect 9772 31948 9828 32510
rect 9548 31892 9828 31948
rect 10108 32562 10164 32574
rect 10108 32510 10110 32562
rect 10162 32510 10164 32562
rect 9548 31778 9604 31892
rect 9548 31726 9550 31778
rect 9602 31726 9604 31778
rect 9548 31714 9604 31726
rect 9324 31614 9326 31666
rect 9378 31614 9380 31666
rect 9324 31602 9380 31614
rect 9884 31554 9940 31566
rect 9884 31502 9886 31554
rect 9938 31502 9940 31554
rect 9884 31444 9940 31502
rect 10108 31556 10164 32510
rect 10668 32564 10724 32574
rect 10668 32470 10724 32508
rect 10668 31780 10724 31790
rect 10668 31686 10724 31724
rect 10332 31556 10388 31566
rect 10108 31500 10332 31556
rect 10332 31462 10388 31500
rect 10780 31556 10836 32622
rect 11004 31556 11060 31566
rect 10780 31462 10836 31500
rect 10892 31554 11060 31556
rect 10892 31502 11006 31554
rect 11058 31502 11060 31554
rect 10892 31500 11060 31502
rect 9212 31388 9940 31444
rect 9212 28196 9268 31388
rect 10892 31108 10948 31500
rect 11004 31490 11060 31500
rect 10556 31052 10948 31108
rect 10108 30996 10164 31006
rect 10108 30902 10164 30940
rect 9660 30882 9716 30894
rect 9660 30830 9662 30882
rect 9714 30830 9716 30882
rect 9660 29876 9716 30830
rect 10332 30436 10388 30446
rect 9996 30212 10052 30222
rect 9660 29810 9716 29820
rect 9772 30156 9996 30212
rect 9436 29540 9492 29550
rect 9436 28644 9492 29484
rect 9436 28550 9492 28588
rect 9548 29092 9604 29102
rect 9324 28196 9380 28206
rect 9212 28140 9324 28196
rect 8988 27746 9044 27758
rect 8988 27694 8990 27746
rect 9042 27694 9044 27746
rect 8988 27412 9044 27694
rect 8988 27356 9268 27412
rect 8876 27244 9156 27300
rect 8540 27186 8596 27198
rect 8540 27134 8542 27186
rect 8594 27134 8596 27186
rect 8540 26908 8596 27134
rect 8316 26852 8932 26908
rect 8316 26402 8372 26852
rect 8876 26514 8932 26852
rect 8876 26462 8878 26514
rect 8930 26462 8932 26514
rect 8876 26450 8932 26462
rect 8988 26516 9044 26526
rect 8316 26350 8318 26402
rect 8370 26350 8372 26402
rect 8316 26338 8372 26350
rect 8988 26402 9044 26460
rect 8988 26350 8990 26402
rect 9042 26350 9044 26402
rect 8988 26338 9044 26350
rect 8652 26292 8708 26302
rect 8652 26198 8708 26236
rect 8204 26114 8260 26124
rect 8365 25900 8629 25910
rect 8421 25844 8469 25900
rect 8525 25844 8573 25900
rect 8365 25834 8629 25844
rect 8540 25732 8596 25742
rect 8540 25638 8596 25676
rect 8204 25620 8260 25630
rect 8204 25526 8260 25564
rect 7980 25342 7982 25394
rect 8034 25342 8036 25394
rect 7532 24164 7588 24174
rect 7532 24070 7588 24108
rect 7644 23940 7700 23950
rect 7420 23884 7644 23940
rect 7644 23846 7700 23884
rect 7868 23828 7924 23838
rect 7308 23772 7476 23828
rect 6524 22258 6580 22270
rect 6524 22206 6526 22258
rect 6578 22206 6580 22258
rect 6524 22148 6580 22206
rect 6972 22148 7028 22428
rect 7196 22418 7252 22428
rect 7308 22820 7364 22830
rect 6188 22092 6356 22148
rect 6524 22092 7028 22148
rect 7084 22258 7140 22270
rect 7084 22206 7086 22258
rect 7138 22206 7140 22258
rect 7084 22148 7140 22206
rect 7308 22148 7364 22764
rect 7420 22484 7476 23772
rect 7868 23734 7924 23772
rect 7532 23714 7588 23726
rect 7532 23662 7534 23714
rect 7586 23662 7588 23714
rect 7532 22820 7588 23662
rect 7532 22754 7588 22764
rect 7756 22596 7812 22606
rect 7756 22502 7812 22540
rect 7420 22428 7588 22484
rect 7084 22092 7364 22148
rect 7420 22258 7476 22270
rect 7420 22206 7422 22258
rect 7474 22206 7476 22258
rect 5628 20130 5908 20132
rect 5628 20078 5630 20130
rect 5682 20078 5908 20130
rect 5628 20076 5908 20078
rect 5628 20066 5684 20076
rect 6188 19908 6244 19918
rect 5964 19906 6244 19908
rect 5964 19854 6190 19906
rect 6242 19854 6244 19906
rect 5964 19852 6244 19854
rect 5740 19236 5796 19246
rect 5740 19142 5796 19180
rect 5852 18562 5908 18574
rect 5852 18510 5854 18562
rect 5906 18510 5908 18562
rect 5516 18452 5572 18462
rect 5852 18452 5908 18510
rect 5572 18396 5908 18452
rect 5516 18358 5572 18396
rect 5852 17666 5908 18396
rect 5852 17614 5854 17666
rect 5906 17614 5908 17666
rect 5852 17602 5908 17614
rect 5628 17444 5684 17454
rect 5628 17350 5684 17388
rect 5964 17220 6020 19852
rect 6188 19842 6244 19852
rect 6300 19684 6356 22092
rect 6188 19628 6356 19684
rect 6412 20690 6468 20702
rect 6412 20638 6414 20690
rect 6466 20638 6468 20690
rect 6076 19122 6132 19134
rect 6076 19070 6078 19122
rect 6130 19070 6132 19122
rect 6076 19012 6132 19070
rect 6076 18946 6132 18956
rect 6188 18676 6244 19628
rect 6300 19124 6356 19134
rect 6300 19030 6356 19068
rect 6412 19010 6468 20638
rect 6636 19906 6692 19918
rect 6636 19854 6638 19906
rect 6690 19854 6692 19906
rect 6636 19460 6692 19854
rect 6748 19796 6804 22092
rect 7420 20132 7476 22206
rect 7196 19906 7252 19918
rect 7196 19854 7198 19906
rect 7250 19854 7252 19906
rect 6748 19730 6804 19740
rect 6860 19794 6916 19806
rect 6860 19742 6862 19794
rect 6914 19742 6916 19794
rect 6636 19404 6804 19460
rect 6524 19236 6580 19246
rect 6524 19142 6580 19180
rect 6748 19012 6804 19404
rect 6412 18958 6414 19010
rect 6466 18958 6468 19010
rect 6412 18946 6468 18958
rect 6636 18956 6804 19012
rect 6860 19234 6916 19742
rect 7196 19794 7252 19854
rect 7196 19742 7198 19794
rect 7250 19742 7252 19794
rect 7196 19730 7252 19742
rect 7420 19572 7476 20076
rect 6860 19182 6862 19234
rect 6914 19182 6916 19234
rect 5628 17164 6020 17220
rect 6076 18620 6244 18676
rect 5516 15428 5572 15438
rect 5516 15334 5572 15372
rect 5628 15092 5684 17164
rect 5964 16772 6020 16782
rect 5628 15026 5684 15036
rect 5740 16770 6020 16772
rect 5740 16718 5966 16770
rect 6018 16718 6020 16770
rect 5740 16716 6020 16718
rect 5740 15538 5796 16716
rect 5964 16706 6020 16716
rect 6076 16660 6132 18620
rect 6188 18450 6244 18462
rect 6188 18398 6190 18450
rect 6242 18398 6244 18450
rect 6188 18228 6244 18398
rect 6524 18452 6580 18462
rect 6524 18358 6580 18396
rect 6412 18340 6468 18350
rect 6188 18162 6244 18172
rect 6300 18284 6412 18340
rect 6300 17108 6356 18284
rect 6412 18274 6468 18284
rect 6412 17668 6468 17678
rect 6412 17574 6468 17612
rect 6412 17108 6468 17118
rect 6300 17106 6468 17108
rect 6300 17054 6414 17106
rect 6466 17054 6468 17106
rect 6300 17052 6468 17054
rect 6300 16884 6356 17052
rect 6412 17042 6468 17052
rect 6300 16818 6356 16828
rect 6076 16604 6468 16660
rect 6300 16324 6356 16334
rect 6300 16098 6356 16268
rect 6300 16046 6302 16098
rect 6354 16046 6356 16098
rect 6300 16034 6356 16046
rect 5740 15486 5742 15538
rect 5794 15486 5796 15538
rect 5740 14532 5796 15486
rect 6076 15876 6132 15886
rect 5964 15316 6020 15326
rect 5964 15222 6020 15260
rect 5740 14466 5796 14476
rect 5852 15090 5908 15102
rect 5852 15038 5854 15090
rect 5906 15038 5908 15090
rect 5852 13748 5908 15038
rect 6076 14308 6132 15820
rect 6412 15148 6468 16604
rect 6524 15428 6580 15438
rect 6524 15334 6580 15372
rect 6076 14214 6132 14252
rect 6188 15092 6468 15148
rect 5852 13682 5908 13692
rect 5852 13524 5908 13534
rect 5740 12852 5796 12862
rect 5628 12738 5684 12750
rect 5628 12686 5630 12738
rect 5682 12686 5684 12738
rect 5516 12628 5572 12638
rect 5516 12402 5572 12572
rect 5516 12350 5518 12402
rect 5570 12350 5572 12402
rect 5516 11844 5572 12350
rect 5516 11778 5572 11788
rect 5628 11396 5684 12686
rect 5740 12068 5796 12796
rect 5740 12002 5796 12012
rect 5628 11330 5684 11340
rect 5852 11394 5908 13468
rect 6076 12066 6132 12078
rect 6076 12014 6078 12066
rect 6130 12014 6132 12066
rect 5852 11342 5854 11394
rect 5906 11342 5908 11394
rect 5404 10994 5460 11004
rect 5740 11284 5796 11294
rect 5740 10834 5796 11228
rect 5852 11172 5908 11342
rect 5964 11396 6020 11406
rect 6076 11396 6132 12014
rect 6020 11340 6132 11396
rect 5964 11282 6020 11340
rect 5964 11230 5966 11282
rect 6018 11230 6020 11282
rect 5964 11218 6020 11230
rect 5852 11106 5908 11116
rect 5740 10782 5742 10834
rect 5794 10782 5796 10834
rect 5740 10770 5796 10782
rect 5404 10500 5460 10510
rect 5852 10500 5908 10510
rect 5404 10498 5908 10500
rect 5404 10446 5406 10498
rect 5458 10446 5854 10498
rect 5906 10446 5908 10498
rect 5404 10444 5908 10446
rect 5404 10434 5460 10444
rect 5180 9938 5348 9940
rect 5180 9886 5182 9938
rect 5234 9886 5348 9938
rect 5180 9884 5348 9886
rect 5180 9874 5236 9884
rect 5292 9716 5348 9726
rect 5068 9202 5124 9212
rect 5180 9604 5236 9614
rect 4956 8988 5124 9044
rect 4620 8370 4676 8988
rect 4956 8820 5012 8830
rect 4620 8318 4622 8370
rect 4674 8318 4676 8370
rect 4620 8306 4676 8318
rect 4844 8764 4956 8820
rect 4508 7646 4510 7698
rect 4562 7646 4564 7698
rect 4508 7634 4564 7646
rect 3500 7476 3556 7486
rect 3500 7474 3668 7476
rect 3500 7422 3502 7474
rect 3554 7422 3668 7474
rect 3500 7420 3668 7422
rect 3500 7410 3556 7420
rect 3388 7196 3556 7252
rect 3276 5966 3278 6018
rect 3330 5966 3332 6018
rect 3276 5954 3332 5966
rect 3500 5234 3556 7196
rect 3612 6916 3668 7420
rect 3612 6850 3668 6860
rect 3948 7362 4004 7374
rect 4732 7364 4788 7374
rect 3948 7310 3950 7362
rect 4002 7310 4004 7362
rect 3948 6132 4004 7310
rect 3948 6066 4004 6076
rect 4620 7308 4732 7364
rect 4620 6356 4676 7308
rect 4732 7298 4788 7308
rect 4732 6804 4788 6814
rect 4844 6804 4900 8764
rect 4956 8754 5012 8764
rect 5068 8596 5124 8988
rect 4956 8540 5124 8596
rect 4956 7698 5012 8540
rect 5180 8370 5236 9548
rect 5180 8318 5182 8370
rect 5234 8318 5236 8370
rect 5180 8306 5236 8318
rect 4956 7646 4958 7698
rect 5010 7646 5012 7698
rect 4956 7634 5012 7646
rect 5292 7028 5348 9660
rect 5404 9044 5460 9054
rect 5404 8950 5460 8988
rect 5628 7700 5684 10444
rect 5852 10434 5908 10444
rect 5852 10276 5908 10286
rect 5852 9938 5908 10220
rect 5852 9886 5854 9938
rect 5906 9886 5908 9938
rect 5852 9874 5908 9886
rect 6188 9604 6244 15092
rect 6636 14980 6692 18956
rect 6860 18564 6916 19182
rect 7196 19346 7252 19358
rect 7196 19294 7198 19346
rect 7250 19294 7252 19346
rect 7196 19236 7252 19294
rect 7196 19170 7252 19180
rect 7308 19012 7364 19022
rect 7420 19012 7476 19516
rect 7532 19348 7588 22428
rect 7980 21588 8036 25342
rect 8316 24836 8372 24846
rect 8204 24780 8316 24836
rect 8092 24612 8148 24622
rect 8092 23826 8148 24556
rect 8204 24164 8260 24780
rect 8316 24770 8372 24780
rect 8652 24612 8708 24622
rect 8652 24518 8708 24556
rect 8365 24332 8629 24342
rect 8421 24276 8469 24332
rect 8525 24276 8573 24332
rect 8365 24266 8629 24276
rect 8204 24108 8372 24164
rect 8204 23940 8260 23950
rect 8204 23846 8260 23884
rect 8092 23774 8094 23826
rect 8146 23774 8148 23826
rect 8092 23762 8148 23774
rect 8092 23042 8148 23054
rect 8092 22990 8094 23042
rect 8146 22990 8148 23042
rect 8092 22820 8148 22990
rect 8316 22932 8372 24108
rect 9100 23492 9156 27244
rect 8428 23436 9156 23492
rect 8428 23378 8484 23436
rect 8428 23326 8430 23378
rect 8482 23326 8484 23378
rect 8428 23314 8484 23326
rect 8092 22754 8148 22764
rect 8204 22876 8372 22932
rect 8764 23154 8820 23166
rect 8764 23102 8766 23154
rect 8818 23102 8820 23154
rect 8092 22596 8148 22606
rect 8204 22596 8260 22876
rect 8365 22764 8629 22774
rect 8421 22708 8469 22764
rect 8525 22708 8573 22764
rect 8365 22698 8629 22708
rect 8092 22594 8260 22596
rect 8092 22542 8094 22594
rect 8146 22542 8260 22594
rect 8092 22540 8260 22542
rect 8092 22530 8148 22540
rect 8764 22372 8820 23102
rect 8764 22260 8820 22316
rect 8988 22260 9044 22270
rect 8764 22258 9044 22260
rect 8764 22206 8990 22258
rect 9042 22206 9044 22258
rect 8764 22204 9044 22206
rect 8988 21924 9044 22204
rect 8988 21858 9044 21868
rect 9100 21812 9156 23436
rect 9212 26964 9268 27356
rect 9212 23268 9268 26908
rect 9324 23548 9380 28140
rect 9548 28082 9604 29036
rect 9772 28868 9828 30156
rect 9996 30118 10052 30156
rect 10220 30100 10276 30110
rect 10108 30098 10276 30100
rect 10108 30046 10222 30098
rect 10274 30046 10276 30098
rect 10108 30044 10276 30046
rect 10108 29092 10164 30044
rect 10220 30034 10276 30044
rect 10220 29876 10276 29886
rect 10220 29426 10276 29820
rect 10220 29374 10222 29426
rect 10274 29374 10276 29426
rect 10220 29362 10276 29374
rect 10108 29026 10164 29036
rect 9548 28030 9550 28082
rect 9602 28030 9604 28082
rect 9548 28018 9604 28030
rect 9660 28812 9828 28868
rect 9884 28868 9940 28878
rect 9884 28866 10164 28868
rect 9884 28814 9886 28866
rect 9938 28814 10164 28866
rect 9884 28812 10164 28814
rect 9660 26908 9716 28812
rect 9884 28802 9940 28812
rect 9436 26852 9716 26908
rect 9772 28644 9828 28654
rect 10108 28644 10164 28812
rect 10220 28644 10276 28654
rect 10108 28642 10276 28644
rect 10108 28590 10222 28642
rect 10274 28590 10276 28642
rect 10108 28588 10276 28590
rect 9772 28420 9828 28588
rect 10220 28578 10276 28588
rect 9996 28530 10052 28542
rect 9996 28478 9998 28530
rect 10050 28478 10052 28530
rect 9884 28420 9940 28430
rect 9772 28418 9940 28420
rect 9772 28366 9886 28418
rect 9938 28366 9940 28418
rect 9772 28364 9940 28366
rect 9436 24052 9492 26852
rect 9772 26404 9828 28364
rect 9884 28354 9940 28364
rect 9884 27858 9940 27870
rect 9884 27806 9886 27858
rect 9938 27806 9940 27858
rect 9884 26964 9940 27806
rect 9996 27188 10052 28478
rect 10332 28084 10388 30380
rect 10556 30210 10612 31052
rect 10780 30882 10836 30894
rect 10780 30830 10782 30882
rect 10834 30830 10836 30882
rect 10668 30324 10724 30334
rect 10780 30324 10836 30830
rect 10668 30322 10836 30324
rect 10668 30270 10670 30322
rect 10722 30270 10836 30322
rect 10668 30268 10836 30270
rect 10668 30258 10724 30268
rect 10556 30158 10558 30210
rect 10610 30158 10612 30210
rect 10556 30146 10612 30158
rect 10780 30100 10836 30110
rect 10780 30006 10836 30044
rect 11116 30098 11172 33294
rect 11116 30046 11118 30098
rect 11170 30046 11172 30098
rect 11116 29876 11172 30046
rect 11116 29810 11172 29820
rect 10892 29316 10948 29326
rect 10444 29314 10948 29316
rect 10444 29262 10894 29314
rect 10946 29262 10948 29314
rect 10444 29260 10948 29262
rect 10444 28754 10500 29260
rect 10892 29250 10948 29260
rect 10444 28702 10446 28754
rect 10498 28702 10500 28754
rect 10444 28690 10500 28702
rect 10668 28756 10724 28766
rect 10668 28642 10724 28700
rect 11116 28644 11172 28654
rect 10668 28590 10670 28642
rect 10722 28590 10724 28642
rect 10668 28578 10724 28590
rect 11004 28642 11172 28644
rect 11004 28590 11118 28642
rect 11170 28590 11172 28642
rect 11004 28588 11172 28590
rect 10892 28530 10948 28542
rect 10892 28478 10894 28530
rect 10946 28478 10948 28530
rect 10780 28084 10836 28094
rect 10332 28082 10780 28084
rect 10332 28030 10334 28082
rect 10386 28030 10780 28082
rect 10332 28028 10780 28030
rect 10332 28018 10388 28028
rect 10780 27990 10836 28028
rect 10668 27858 10724 27870
rect 10668 27806 10670 27858
rect 10722 27806 10724 27858
rect 10668 27188 10724 27806
rect 10892 27300 10948 28478
rect 11004 28082 11060 28588
rect 11116 28578 11172 28588
rect 11228 28420 11284 36764
rect 11676 35700 11732 35710
rect 11676 35698 11844 35700
rect 11676 35646 11678 35698
rect 11730 35646 11844 35698
rect 11676 35644 11844 35646
rect 11676 35634 11732 35644
rect 11788 35026 11844 35644
rect 11900 35588 11956 39200
rect 14140 39060 14196 39200
rect 14476 39060 14532 39228
rect 14140 39004 14532 39060
rect 13804 37380 13860 37390
rect 12236 37044 12292 37054
rect 12124 35588 12180 35598
rect 11900 35586 12180 35588
rect 11900 35534 12126 35586
rect 12178 35534 12180 35586
rect 11900 35532 12180 35534
rect 12124 35522 12180 35532
rect 11788 34974 11790 35026
rect 11842 34974 11844 35026
rect 11788 34962 11844 34974
rect 12124 35364 12180 35374
rect 12124 34802 12180 35308
rect 12124 34750 12126 34802
rect 12178 34750 12180 34802
rect 12124 34738 12180 34750
rect 11564 34468 11620 34478
rect 11564 33458 11620 34412
rect 11676 34356 11732 34366
rect 11900 34356 11956 34366
rect 11732 34300 11844 34356
rect 11676 34290 11732 34300
rect 11788 33684 11844 34300
rect 11900 34262 11956 34300
rect 11788 33618 11844 33628
rect 11564 33406 11566 33458
rect 11618 33406 11620 33458
rect 11564 33394 11620 33406
rect 12012 33460 12068 33470
rect 12012 33366 12068 33404
rect 11788 32788 11844 32798
rect 11788 32694 11844 32732
rect 11452 32452 11508 32462
rect 11452 32358 11508 32396
rect 11340 30212 11396 30222
rect 11340 30118 11396 30156
rect 12236 28868 12292 36988
rect 12572 36596 12628 36606
rect 12572 36502 12628 36540
rect 13244 36260 13300 36270
rect 13132 36204 13244 36260
rect 13132 35700 13188 36204
rect 13244 36166 13300 36204
rect 13692 36260 13748 36270
rect 13692 36166 13748 36204
rect 13804 35812 13860 37324
rect 14364 36596 14420 36606
rect 14364 36482 14420 36540
rect 14812 36594 14868 39228
rect 16352 39200 16464 40000
rect 18592 39200 18704 40000
rect 18956 39228 19348 39284
rect 16380 36932 16436 39200
rect 18620 39060 18676 39200
rect 18956 39060 19012 39228
rect 18620 39004 19012 39060
rect 16380 36866 16436 36876
rect 17388 36932 17444 36942
rect 14812 36542 14814 36594
rect 14866 36542 14868 36594
rect 14812 36530 14868 36542
rect 17388 36594 17444 36876
rect 17388 36542 17390 36594
rect 17442 36542 17444 36594
rect 17388 36530 17444 36542
rect 18060 36596 18116 36606
rect 14364 36430 14366 36482
rect 14418 36430 14420 36482
rect 14364 36418 14420 36430
rect 12796 35698 13188 35700
rect 12796 35646 13134 35698
rect 13186 35646 13188 35698
rect 12796 35644 13188 35646
rect 12796 35588 12852 35644
rect 13132 35634 13188 35644
rect 13692 35756 13860 35812
rect 14028 36372 14084 36382
rect 12348 34914 12404 34926
rect 12348 34862 12350 34914
rect 12402 34862 12404 34914
rect 12348 34018 12404 34862
rect 12796 34356 12852 35532
rect 13132 35476 13188 35486
rect 13020 34804 13076 34814
rect 13020 34710 13076 34748
rect 12796 34130 12852 34300
rect 12796 34078 12798 34130
rect 12850 34078 12852 34130
rect 12796 34066 12852 34078
rect 12348 33966 12350 34018
rect 12402 33966 12404 34018
rect 12348 31948 12404 33966
rect 12908 34020 12964 34030
rect 12572 33684 12628 33694
rect 12572 33458 12628 33628
rect 12572 33406 12574 33458
rect 12626 33406 12628 33458
rect 12572 33394 12628 33406
rect 12908 33458 12964 33964
rect 12908 33406 12910 33458
rect 12962 33406 12964 33458
rect 12908 33394 12964 33406
rect 13020 33236 13076 33246
rect 13020 32338 13076 33180
rect 13020 32286 13022 32338
rect 13074 32286 13076 32338
rect 13020 32274 13076 32286
rect 12348 31892 12852 31948
rect 12796 29092 12852 31892
rect 12908 31556 12964 31566
rect 12908 30882 12964 31500
rect 12908 30830 12910 30882
rect 12962 30830 12964 30882
rect 12908 30818 12964 30830
rect 13132 29988 13188 35420
rect 13468 34020 13524 34030
rect 13468 34018 13636 34020
rect 13468 33966 13470 34018
rect 13522 33966 13636 34018
rect 13468 33964 13636 33966
rect 13468 33954 13524 33964
rect 13580 33234 13636 33964
rect 13580 33182 13582 33234
rect 13634 33182 13636 33234
rect 13580 33170 13636 33182
rect 13244 32562 13300 32574
rect 13244 32510 13246 32562
rect 13298 32510 13300 32562
rect 13244 31780 13300 32510
rect 13692 31948 13748 35756
rect 13804 35586 13860 35598
rect 13804 35534 13806 35586
rect 13858 35534 13860 35586
rect 13804 34802 13860 35534
rect 13804 34750 13806 34802
rect 13858 34750 13860 34802
rect 13804 34738 13860 34750
rect 13916 33236 13972 33246
rect 13916 33142 13972 33180
rect 14028 31948 14084 36316
rect 15820 36372 15876 36382
rect 15820 36278 15876 36316
rect 16492 36372 16548 36382
rect 15148 36260 15204 36270
rect 14924 35028 14980 35038
rect 15148 35028 15204 36204
rect 16156 36260 16212 36270
rect 16156 36166 16212 36204
rect 15518 36092 15782 36102
rect 15574 36036 15622 36092
rect 15678 36036 15726 36092
rect 15518 36026 15782 36036
rect 16268 35812 16324 35822
rect 16044 35810 16324 35812
rect 16044 35758 16270 35810
rect 16322 35758 16324 35810
rect 16044 35756 16324 35758
rect 15932 35588 15988 35598
rect 15932 35494 15988 35532
rect 14364 35026 15204 35028
rect 14364 34974 14926 35026
rect 14978 34974 15204 35026
rect 14364 34972 15204 34974
rect 14140 34804 14196 34814
rect 14140 34710 14196 34748
rect 14364 33458 14420 34972
rect 14924 34962 14980 34972
rect 15148 34916 15204 34972
rect 15932 35140 15988 35150
rect 15260 34916 15316 34926
rect 15148 34914 15316 34916
rect 15148 34862 15262 34914
rect 15314 34862 15316 34914
rect 15148 34860 15316 34862
rect 15260 34850 15316 34860
rect 15518 34524 15782 34534
rect 15574 34468 15622 34524
rect 15678 34468 15726 34524
rect 15518 34458 15782 34468
rect 15932 34356 15988 35084
rect 16044 35026 16100 35756
rect 16268 35746 16324 35756
rect 16492 35698 16548 36316
rect 16492 35646 16494 35698
rect 16546 35646 16548 35698
rect 16492 35634 16548 35646
rect 16940 36258 16996 36270
rect 16940 36206 16942 36258
rect 16994 36206 16996 36258
rect 16940 35588 16996 36206
rect 16940 35522 16996 35532
rect 17836 35586 17892 35598
rect 17836 35534 17838 35586
rect 17890 35534 17892 35586
rect 16044 34974 16046 35026
rect 16098 34974 16100 35026
rect 16044 34962 16100 34974
rect 15596 34300 15988 34356
rect 17724 34804 17780 34814
rect 15596 34018 15652 34300
rect 16604 34244 16660 34254
rect 16604 34242 16772 34244
rect 16604 34190 16606 34242
rect 16658 34190 16772 34242
rect 16604 34188 16772 34190
rect 16604 34178 16660 34188
rect 16268 34132 16324 34142
rect 15596 33966 15598 34018
rect 15650 33966 15652 34018
rect 15596 33954 15652 33966
rect 15708 34130 16324 34132
rect 15708 34078 16270 34130
rect 16322 34078 16324 34130
rect 15708 34076 16324 34078
rect 14364 33406 14366 33458
rect 14418 33406 14420 33458
rect 14364 33394 14420 33406
rect 14924 33458 14980 33470
rect 14924 33406 14926 33458
rect 14978 33406 14980 33458
rect 14588 32564 14644 32574
rect 14588 32470 14644 32508
rect 14700 32450 14756 32462
rect 14700 32398 14702 32450
rect 14754 32398 14756 32450
rect 14700 32340 14756 32398
rect 14700 32274 14756 32284
rect 13244 31714 13300 31724
rect 13468 31892 13748 31948
rect 13916 31892 14084 31948
rect 13132 29932 13412 29988
rect 12796 29026 12852 29036
rect 12908 29652 12964 29662
rect 13356 29652 13412 29932
rect 11900 28812 12292 28868
rect 12796 28866 12852 28878
rect 12796 28814 12798 28866
rect 12850 28814 12852 28866
rect 11452 28644 11508 28654
rect 11452 28550 11508 28588
rect 11676 28642 11732 28654
rect 11676 28590 11678 28642
rect 11730 28590 11732 28642
rect 11228 28354 11284 28364
rect 11452 28420 11508 28430
rect 11452 28326 11508 28364
rect 11004 28030 11006 28082
rect 11058 28030 11060 28082
rect 11004 28018 11060 28030
rect 11452 27860 11508 27870
rect 11452 27766 11508 27804
rect 10892 27244 11060 27300
rect 9996 27132 10724 27188
rect 9996 26964 10052 26974
rect 9884 26908 9996 26964
rect 9996 26870 10052 26908
rect 9772 26348 9940 26404
rect 9772 26180 9828 26190
rect 9772 24164 9828 26124
rect 9884 25060 9940 26348
rect 10108 26290 10164 27132
rect 10892 27076 10948 27086
rect 10444 27074 10948 27076
rect 10444 27022 10894 27074
rect 10946 27022 10948 27074
rect 10444 27020 10948 27022
rect 10332 26964 10388 26974
rect 10332 26870 10388 26908
rect 10444 26514 10500 27020
rect 10892 27010 10948 27020
rect 10668 26852 10724 26862
rect 11004 26852 11060 27244
rect 11228 27076 11284 27114
rect 11228 27010 11284 27020
rect 11564 26964 11620 26974
rect 11676 26964 11732 28590
rect 11788 27076 11844 27086
rect 11788 26982 11844 27020
rect 11564 26962 11732 26964
rect 11564 26910 11566 26962
rect 11618 26910 11732 26962
rect 11564 26908 11732 26910
rect 10668 26850 11060 26852
rect 10668 26798 10670 26850
rect 10722 26798 11060 26850
rect 10668 26796 11060 26798
rect 10668 26786 10724 26796
rect 10444 26462 10446 26514
rect 10498 26462 10500 26514
rect 10444 26450 10500 26462
rect 10108 26238 10110 26290
rect 10162 26238 10164 26290
rect 10108 25396 10164 26238
rect 10220 26402 10276 26414
rect 10220 26350 10222 26402
rect 10274 26350 10276 26402
rect 10220 26180 10276 26350
rect 10220 26114 10276 26124
rect 10780 26290 10836 26302
rect 10780 26238 10782 26290
rect 10834 26238 10836 26290
rect 10780 25620 10836 26238
rect 11004 26180 11060 26796
rect 11228 26850 11284 26862
rect 11228 26798 11230 26850
rect 11282 26798 11284 26850
rect 11228 26404 11284 26798
rect 11452 26404 11508 26414
rect 11228 26402 11508 26404
rect 11228 26350 11454 26402
rect 11506 26350 11508 26402
rect 11228 26348 11508 26350
rect 11452 26338 11508 26348
rect 11564 26180 11620 26908
rect 11004 26124 11620 26180
rect 10780 25564 11060 25620
rect 10332 25396 10388 25406
rect 10108 25394 10388 25396
rect 10108 25342 10334 25394
rect 10386 25342 10388 25394
rect 10108 25340 10388 25342
rect 9996 25284 10052 25294
rect 9996 25190 10052 25228
rect 10332 25060 10388 25340
rect 10668 25396 10724 25406
rect 10892 25396 10948 25406
rect 10668 25394 10948 25396
rect 10668 25342 10670 25394
rect 10722 25342 10894 25394
rect 10946 25342 10948 25394
rect 10668 25340 10948 25342
rect 10668 25330 10724 25340
rect 10892 25330 10948 25340
rect 10444 25284 10500 25294
rect 10444 25190 10500 25228
rect 9884 25004 10276 25060
rect 10332 25004 10500 25060
rect 10220 24164 10276 25004
rect 9772 24108 9940 24164
rect 9436 24050 9828 24052
rect 9436 23998 9438 24050
rect 9490 23998 9828 24050
rect 9436 23996 9828 23998
rect 9436 23986 9492 23996
rect 9324 23492 9716 23548
rect 9212 23202 9268 23212
rect 9100 21746 9156 21756
rect 9212 22932 9268 22942
rect 8652 21700 8708 21710
rect 8652 21698 8820 21700
rect 8652 21646 8654 21698
rect 8706 21646 8820 21698
rect 8652 21644 8820 21646
rect 8652 21634 8708 21644
rect 8204 21588 8260 21598
rect 7980 21586 8260 21588
rect 7980 21534 8206 21586
rect 8258 21534 8260 21586
rect 7980 21532 8260 21534
rect 7756 21474 7812 21486
rect 7756 21422 7758 21474
rect 7810 21422 7812 21474
rect 7756 19572 7812 21422
rect 8204 20916 8260 21532
rect 8540 21364 8596 21402
rect 8540 21298 8596 21308
rect 8365 21196 8629 21206
rect 8421 21140 8469 21196
rect 8525 21140 8573 21196
rect 8365 21130 8629 21140
rect 8540 20916 8596 20926
rect 8204 20914 8596 20916
rect 8204 20862 8542 20914
rect 8594 20862 8596 20914
rect 8204 20860 8596 20862
rect 8764 20916 8820 21644
rect 8876 21364 8932 21374
rect 8876 21362 9156 21364
rect 8876 21310 8878 21362
rect 8930 21310 9156 21362
rect 8876 21308 9156 21310
rect 8876 21298 8932 21308
rect 9100 21026 9156 21308
rect 9100 20974 9102 21026
rect 9154 20974 9156 21026
rect 8876 20916 8932 20926
rect 8764 20914 9044 20916
rect 8764 20862 8878 20914
rect 8930 20862 9044 20914
rect 8764 20860 9044 20862
rect 8540 20850 8596 20860
rect 8876 20850 8932 20860
rect 8652 20130 8708 20142
rect 8652 20078 8654 20130
rect 8706 20078 8708 20130
rect 8092 20020 8148 20030
rect 8316 20020 8372 20030
rect 8092 20018 8372 20020
rect 8092 19966 8094 20018
rect 8146 19966 8318 20018
rect 8370 19966 8372 20018
rect 8092 19964 8372 19966
rect 8092 19954 8148 19964
rect 7756 19506 7812 19516
rect 8092 19460 8148 19470
rect 7532 19292 7924 19348
rect 7308 19010 7476 19012
rect 7308 18958 7310 19010
rect 7362 18958 7476 19010
rect 7308 18956 7476 18958
rect 7308 18946 7364 18956
rect 6748 18562 6916 18564
rect 6748 18510 6862 18562
rect 6914 18510 6916 18562
rect 6748 18508 6916 18510
rect 6748 16324 6804 18508
rect 6860 18498 6916 18508
rect 7308 18340 7364 18350
rect 7308 18246 7364 18284
rect 7196 17780 7252 17790
rect 7084 17724 7196 17780
rect 7084 17666 7140 17724
rect 7196 17714 7252 17724
rect 7084 17614 7086 17666
rect 7138 17614 7140 17666
rect 7084 17602 7140 17614
rect 6972 16996 7028 17006
rect 6972 16770 7028 16940
rect 6972 16718 6974 16770
rect 7026 16718 7028 16770
rect 6972 16706 7028 16718
rect 7196 16660 7252 16670
rect 6748 16268 6916 16324
rect 6748 16100 6804 16110
rect 6748 15314 6804 16044
rect 6748 15262 6750 15314
rect 6802 15262 6804 15314
rect 6748 15250 6804 15262
rect 6860 15148 6916 16268
rect 6636 14914 6692 14924
rect 6748 15092 6916 15148
rect 6972 16210 7028 16222
rect 6972 16158 6974 16210
rect 7026 16158 7028 16210
rect 6748 14532 6804 15092
rect 6636 14476 6804 14532
rect 6860 14754 6916 14766
rect 6860 14702 6862 14754
rect 6914 14702 6916 14754
rect 6860 14642 6916 14702
rect 6860 14590 6862 14642
rect 6914 14590 6916 14642
rect 6412 14306 6468 14318
rect 6412 14254 6414 14306
rect 6466 14254 6468 14306
rect 6412 14084 6468 14254
rect 6300 13748 6356 13758
rect 6412 13748 6468 14028
rect 6300 13746 6468 13748
rect 6300 13694 6302 13746
rect 6354 13694 6468 13746
rect 6300 13692 6468 13694
rect 6300 13636 6356 13692
rect 6300 13570 6356 13580
rect 6524 13522 6580 13534
rect 6524 13470 6526 13522
rect 6578 13470 6580 13522
rect 6524 13076 6580 13470
rect 6636 13524 6692 14476
rect 6748 13748 6804 13758
rect 6860 13748 6916 14590
rect 6972 14644 7028 16158
rect 7196 16098 7252 16604
rect 7196 16046 7198 16098
rect 7250 16046 7252 16098
rect 7196 16034 7252 16046
rect 7420 15876 7476 18956
rect 7532 19122 7588 19134
rect 7532 19070 7534 19122
rect 7586 19070 7588 19122
rect 7532 19012 7588 19070
rect 7532 18676 7588 18956
rect 7532 18610 7588 18620
rect 7644 18450 7700 18462
rect 7644 18398 7646 18450
rect 7698 18398 7700 18450
rect 7644 18228 7700 18398
rect 6972 14578 7028 14588
rect 7196 15820 7476 15876
rect 7532 17668 7588 17678
rect 7644 17668 7700 18172
rect 7532 17666 7700 17668
rect 7532 17614 7534 17666
rect 7586 17614 7700 17666
rect 7532 17612 7700 17614
rect 6748 13746 6916 13748
rect 6748 13694 6750 13746
rect 6802 13694 6916 13746
rect 6748 13692 6916 13694
rect 6748 13682 6804 13692
rect 7084 13636 7140 13646
rect 6636 13468 6804 13524
rect 6300 13074 6580 13076
rect 6300 13022 6526 13074
rect 6578 13022 6580 13074
rect 6300 13020 6580 13022
rect 6300 12178 6356 13020
rect 6524 13010 6580 13020
rect 6636 12852 6692 12862
rect 6636 12758 6692 12796
rect 6748 12740 6804 13468
rect 6748 12674 6804 12684
rect 7084 12292 7140 13580
rect 7196 12404 7252 15820
rect 7420 15426 7476 15438
rect 7420 15374 7422 15426
rect 7474 15374 7476 15426
rect 7308 15092 7364 15102
rect 7308 14754 7364 15036
rect 7308 14702 7310 14754
rect 7362 14702 7364 14754
rect 7308 14642 7364 14702
rect 7308 14590 7310 14642
rect 7362 14590 7364 14642
rect 7308 14420 7364 14590
rect 7308 14354 7364 14364
rect 7308 13860 7364 13870
rect 7308 13766 7364 13804
rect 7196 12348 7364 12404
rect 7084 12236 7252 12292
rect 6300 12126 6302 12178
rect 6354 12126 6356 12178
rect 6300 11732 6356 12126
rect 6636 12180 6692 12190
rect 6972 12180 7028 12190
rect 6636 12178 7028 12180
rect 6636 12126 6638 12178
rect 6690 12126 6974 12178
rect 7026 12126 7028 12178
rect 6636 12124 7028 12126
rect 6636 12114 6692 12124
rect 6972 12114 7028 12124
rect 7196 12178 7252 12236
rect 7196 12126 7198 12178
rect 7250 12126 7252 12178
rect 7196 12114 7252 12126
rect 7084 12066 7140 12078
rect 7084 12014 7086 12066
rect 7138 12014 7140 12066
rect 7084 11956 7140 12014
rect 6300 11666 6356 11676
rect 6972 11900 7140 11956
rect 6636 11396 6692 11406
rect 6300 11170 6356 11182
rect 6300 11118 6302 11170
rect 6354 11118 6356 11170
rect 6300 9826 6356 11118
rect 6412 11172 6468 11182
rect 6412 10498 6468 11116
rect 6636 10610 6692 11340
rect 6748 11394 6804 11406
rect 6748 11342 6750 11394
rect 6802 11342 6804 11394
rect 6748 11284 6804 11342
rect 6748 11218 6804 11228
rect 6636 10558 6638 10610
rect 6690 10558 6692 10610
rect 6636 10546 6692 10558
rect 6412 10446 6414 10498
rect 6466 10446 6468 10498
rect 6412 10434 6468 10446
rect 6300 9774 6302 9826
rect 6354 9774 6356 9826
rect 6300 9762 6356 9774
rect 6748 10386 6804 10398
rect 6748 10334 6750 10386
rect 6802 10334 6804 10386
rect 6748 9714 6804 10334
rect 6748 9662 6750 9714
rect 6802 9662 6804 9714
rect 6748 9650 6804 9662
rect 6188 9538 6244 9548
rect 6748 9380 6804 9390
rect 6300 9268 6356 9278
rect 6188 9212 6300 9268
rect 5852 9154 5908 9166
rect 5852 9102 5854 9154
rect 5906 9102 5908 9154
rect 5852 9044 5908 9102
rect 5852 8978 5908 8988
rect 6188 8258 6244 9212
rect 6300 9202 6356 9212
rect 6748 9266 6804 9324
rect 6748 9214 6750 9266
rect 6802 9214 6804 9266
rect 6748 9202 6804 9214
rect 6972 9268 7028 11900
rect 7084 11732 7140 11742
rect 7084 11282 7140 11676
rect 7084 11230 7086 11282
rect 7138 11230 7140 11282
rect 7084 11218 7140 11230
rect 7308 10388 7364 12348
rect 7420 10610 7476 15374
rect 7532 13300 7588 17612
rect 7756 17442 7812 17454
rect 7756 17390 7758 17442
rect 7810 17390 7812 17442
rect 7756 17220 7812 17390
rect 7756 17154 7812 17164
rect 7756 16882 7812 16894
rect 7756 16830 7758 16882
rect 7810 16830 7812 16882
rect 7644 16772 7700 16782
rect 7644 16678 7700 16716
rect 7756 15988 7812 16830
rect 7756 15922 7812 15932
rect 7868 15314 7924 19292
rect 8092 19234 8148 19404
rect 8092 19182 8094 19234
rect 8146 19182 8148 19234
rect 8092 19170 8148 19182
rect 8204 19348 8260 19964
rect 8316 19954 8372 19964
rect 8652 19796 8708 20078
rect 8876 19796 8932 19806
rect 8652 19730 8708 19740
rect 8764 19794 8932 19796
rect 8764 19742 8878 19794
rect 8930 19742 8932 19794
rect 8764 19740 8932 19742
rect 8365 19628 8629 19638
rect 8421 19572 8469 19628
rect 8525 19572 8573 19628
rect 8365 19562 8629 19572
rect 8540 19460 8596 19470
rect 8764 19460 8820 19740
rect 8876 19730 8932 19740
rect 8540 19458 8820 19460
rect 8540 19406 8542 19458
rect 8594 19406 8820 19458
rect 8540 19404 8820 19406
rect 8988 19458 9044 20860
rect 9100 20020 9156 20974
rect 9100 19954 9156 19964
rect 9100 19796 9156 19806
rect 9212 19796 9268 22876
rect 9324 22708 9380 22718
rect 9324 22258 9380 22652
rect 9660 22484 9716 23492
rect 9772 23492 9828 23996
rect 9772 23154 9828 23436
rect 9772 23102 9774 23154
rect 9826 23102 9828 23154
rect 9772 23090 9828 23102
rect 9324 22206 9326 22258
rect 9378 22206 9380 22258
rect 9324 22194 9380 22206
rect 9436 22428 9716 22484
rect 9100 19794 9268 19796
rect 9100 19742 9102 19794
rect 9154 19742 9268 19794
rect 9100 19740 9268 19742
rect 9324 21924 9380 21934
rect 9100 19730 9156 19740
rect 9324 19572 9380 21868
rect 9436 21026 9492 22428
rect 9884 22372 9940 24108
rect 9436 20974 9438 21026
rect 9490 20974 9492 21026
rect 9436 20962 9492 20974
rect 9660 22316 9940 22372
rect 10220 24050 10276 24108
rect 10220 23998 10222 24050
rect 10274 23998 10276 24050
rect 9660 20580 9716 22316
rect 10108 22260 10164 22270
rect 9772 22146 9828 22158
rect 9772 22094 9774 22146
rect 9826 22094 9828 22146
rect 9772 22036 9828 22094
rect 9828 21980 10052 22036
rect 9772 21970 9828 21980
rect 9996 21810 10052 21980
rect 9996 21758 9998 21810
rect 10050 21758 10052 21810
rect 9996 21746 10052 21758
rect 10108 21698 10164 22204
rect 10108 21646 10110 21698
rect 10162 21646 10164 21698
rect 10108 21634 10164 21646
rect 9996 21364 10052 21374
rect 9996 21270 10052 21308
rect 9772 20580 9828 20590
rect 9660 20524 9772 20580
rect 8988 19406 8990 19458
rect 9042 19406 9044 19458
rect 8540 19394 8596 19404
rect 8204 18450 8260 19292
rect 8316 19124 8372 19134
rect 8988 19124 9044 19406
rect 8372 19068 8484 19124
rect 8316 19030 8372 19068
rect 8428 18564 8484 19068
rect 8988 19058 9044 19068
rect 9100 19516 9380 19572
rect 9100 18900 9156 19516
rect 8988 18844 9156 18900
rect 9212 19234 9268 19246
rect 9212 19182 9214 19234
rect 9266 19182 9268 19234
rect 8652 18676 8708 18686
rect 8652 18582 8708 18620
rect 8540 18564 8596 18574
rect 8428 18562 8596 18564
rect 8428 18510 8542 18562
rect 8594 18510 8596 18562
rect 8428 18508 8596 18510
rect 8540 18498 8596 18508
rect 8204 18398 8206 18450
rect 8258 18398 8260 18450
rect 8204 18386 8260 18398
rect 8876 18450 8932 18462
rect 8876 18398 8878 18450
rect 8930 18398 8932 18450
rect 8365 18060 8629 18070
rect 8421 18004 8469 18060
rect 8525 18004 8573 18060
rect 8365 17994 8629 18004
rect 7868 15262 7870 15314
rect 7922 15262 7924 15314
rect 7644 14532 7700 14542
rect 7644 14438 7700 14476
rect 7868 14532 7924 15262
rect 7980 17780 8036 17790
rect 7980 15202 8036 17724
rect 8540 17668 8596 17678
rect 8540 17574 8596 17612
rect 8316 16996 8372 17006
rect 8092 16994 8372 16996
rect 8092 16942 8318 16994
rect 8370 16942 8372 16994
rect 8092 16940 8372 16942
rect 8092 16436 8148 16940
rect 8316 16930 8372 16940
rect 8876 16996 8932 18398
rect 8988 17220 9044 18844
rect 9212 18452 9268 19182
rect 9436 19236 9492 19246
rect 9436 19234 9604 19236
rect 9436 19182 9438 19234
rect 9490 19182 9604 19234
rect 9436 19180 9604 19182
rect 9436 19170 9492 19180
rect 9212 18386 9268 18396
rect 9436 18452 9492 18462
rect 9436 17554 9492 18396
rect 9548 17780 9604 19180
rect 9772 18900 9828 20524
rect 10220 20244 10276 23998
rect 10332 24722 10388 24734
rect 10332 24670 10334 24722
rect 10386 24670 10388 24722
rect 10332 22820 10388 24670
rect 10444 23828 10500 25004
rect 11004 24276 11060 25564
rect 11452 25508 11508 25518
rect 11564 25508 11620 26124
rect 11452 25506 11620 25508
rect 11452 25454 11454 25506
rect 11506 25454 11620 25506
rect 11452 25452 11620 25454
rect 11900 25620 11956 28812
rect 12796 28756 12852 28814
rect 12796 28690 12852 28700
rect 12012 28644 12068 28654
rect 12012 28550 12068 28588
rect 12236 28644 12292 28654
rect 12236 28530 12292 28588
rect 12236 28478 12238 28530
rect 12290 28478 12292 28530
rect 12236 28466 12292 28478
rect 12348 28532 12404 28542
rect 12684 28532 12740 28542
rect 12348 28530 12740 28532
rect 12348 28478 12350 28530
rect 12402 28478 12686 28530
rect 12738 28478 12740 28530
rect 12348 28476 12740 28478
rect 12124 28420 12180 28430
rect 12124 27970 12180 28364
rect 12124 27918 12126 27970
rect 12178 27918 12180 27970
rect 12124 27906 12180 27918
rect 12012 26964 12068 26974
rect 12012 26870 12068 26908
rect 12124 26964 12180 26974
rect 12348 26964 12404 28476
rect 12684 28466 12740 28476
rect 12796 28532 12852 28542
rect 12908 28532 12964 29596
rect 13132 29596 13412 29652
rect 13020 29314 13076 29326
rect 13020 29262 13022 29314
rect 13074 29262 13076 29314
rect 13020 29204 13076 29262
rect 13020 29138 13076 29148
rect 12796 28530 12964 28532
rect 12796 28478 12798 28530
rect 12850 28478 12964 28530
rect 12796 28476 12964 28478
rect 12796 28466 12852 28476
rect 13132 27972 13188 29596
rect 13356 29428 13412 29438
rect 13132 27906 13188 27916
rect 13244 29092 13300 29102
rect 12124 26962 12404 26964
rect 12124 26910 12126 26962
rect 12178 26910 12404 26962
rect 12124 26908 12404 26910
rect 12684 26964 12740 26974
rect 12012 26516 12068 26526
rect 12124 26516 12180 26908
rect 12684 26870 12740 26908
rect 12068 26460 12180 26516
rect 12012 26450 12068 26460
rect 11452 25442 11508 25452
rect 11228 25396 11284 25406
rect 11228 25302 11284 25340
rect 11676 25396 11732 25406
rect 11676 25302 11732 25340
rect 11900 25394 11956 25564
rect 12460 25620 12516 25630
rect 12460 25526 12516 25564
rect 12012 25508 12068 25518
rect 12012 25414 12068 25452
rect 11900 25342 11902 25394
rect 11954 25342 11956 25394
rect 11900 25330 11956 25342
rect 11116 25282 11172 25294
rect 11116 25230 11118 25282
rect 11170 25230 11172 25282
rect 11116 24834 11172 25230
rect 11116 24782 11118 24834
rect 11170 24782 11172 24834
rect 11116 24770 11172 24782
rect 12796 25284 12852 25294
rect 11004 24210 11060 24220
rect 11116 24164 11172 24174
rect 11172 24108 11396 24164
rect 11116 24098 11172 24108
rect 10892 23940 10948 23950
rect 10892 23938 11284 23940
rect 10892 23886 10894 23938
rect 10946 23886 11284 23938
rect 10892 23884 11284 23886
rect 10892 23874 10948 23884
rect 10556 23828 10612 23838
rect 10444 23826 10612 23828
rect 10444 23774 10558 23826
rect 10610 23774 10612 23826
rect 10444 23772 10612 23774
rect 10556 23762 10612 23772
rect 11116 23714 11172 23726
rect 11116 23662 11118 23714
rect 11170 23662 11172 23714
rect 10556 23044 10612 23054
rect 10556 23042 11060 23044
rect 10556 22990 10558 23042
rect 10610 22990 11060 23042
rect 10556 22988 11060 22990
rect 10556 22978 10612 22988
rect 10332 22764 10500 22820
rect 10332 22146 10388 22158
rect 10332 22094 10334 22146
rect 10386 22094 10388 22146
rect 10332 21364 10388 22094
rect 10444 21588 10500 22764
rect 10892 22708 10948 22718
rect 10892 22370 10948 22652
rect 11004 22482 11060 22988
rect 11004 22430 11006 22482
rect 11058 22430 11060 22482
rect 11004 22418 11060 22430
rect 10892 22318 10894 22370
rect 10946 22318 10948 22370
rect 10892 22306 10948 22318
rect 11116 22370 11172 23662
rect 11116 22318 11118 22370
rect 11170 22318 11172 22370
rect 11116 22306 11172 22318
rect 10444 21494 10500 21532
rect 10556 22258 10612 22270
rect 10556 22206 10558 22258
rect 10610 22206 10612 22258
rect 10556 21364 10612 22206
rect 10332 21308 10612 21364
rect 10668 21812 10724 21822
rect 10332 20468 10388 21308
rect 10668 20916 10724 21756
rect 11228 21700 11284 23884
rect 11340 23826 11396 24108
rect 11340 23774 11342 23826
rect 11394 23774 11396 23826
rect 11340 23762 11396 23774
rect 11452 23828 11508 23838
rect 11900 23828 11956 23838
rect 11452 23826 11956 23828
rect 11452 23774 11454 23826
rect 11506 23774 11902 23826
rect 11954 23774 11956 23826
rect 11452 23772 11956 23774
rect 11452 22372 11508 23772
rect 11900 23762 11956 23772
rect 12012 23828 12068 23838
rect 12012 23734 12068 23772
rect 12572 23828 12628 23838
rect 12124 23716 12180 23726
rect 11676 22372 11732 22382
rect 11452 22370 11732 22372
rect 11452 22318 11678 22370
rect 11730 22318 11732 22370
rect 11452 22316 11732 22318
rect 11340 22260 11396 22270
rect 11396 22204 11508 22260
rect 11340 22194 11396 22204
rect 11452 22146 11508 22204
rect 11452 22094 11454 22146
rect 11506 22094 11508 22146
rect 11452 22082 11508 22094
rect 11116 21644 11284 21700
rect 10668 20822 10724 20860
rect 10892 21364 10948 21374
rect 10892 20802 10948 21308
rect 10892 20750 10894 20802
rect 10946 20750 10948 20802
rect 10892 20738 10948 20750
rect 10332 20402 10388 20412
rect 10220 20188 10948 20244
rect 10780 20020 10836 20030
rect 10668 19964 10780 20020
rect 9884 19906 9940 19918
rect 9884 19854 9886 19906
rect 9938 19854 9940 19906
rect 9884 19124 9940 19854
rect 10332 19906 10388 19918
rect 10332 19854 10334 19906
rect 10386 19854 10388 19906
rect 10332 19572 10388 19854
rect 10332 19506 10388 19516
rect 10556 19906 10612 19918
rect 10556 19854 10558 19906
rect 10610 19854 10612 19906
rect 9996 19348 10052 19358
rect 9996 19346 10500 19348
rect 9996 19294 9998 19346
rect 10050 19294 10500 19346
rect 9996 19292 10500 19294
rect 9996 19282 10052 19292
rect 9884 19122 10052 19124
rect 9884 19070 9886 19122
rect 9938 19070 10052 19122
rect 9884 19068 10052 19070
rect 9884 19058 9940 19068
rect 9772 18844 9940 18900
rect 9548 17714 9604 17724
rect 9772 18226 9828 18238
rect 9772 18174 9774 18226
rect 9826 18174 9828 18226
rect 9436 17502 9438 17554
rect 9490 17502 9492 17554
rect 9436 17490 9492 17502
rect 9660 17666 9716 17678
rect 9660 17614 9662 17666
rect 9714 17614 9716 17666
rect 8988 17154 9044 17164
rect 9100 17442 9156 17454
rect 9100 17390 9102 17442
rect 9154 17390 9156 17442
rect 9100 17108 9156 17390
rect 9100 17042 9156 17052
rect 9436 17220 9492 17230
rect 8876 16930 8932 16940
rect 8540 16882 8596 16894
rect 8540 16830 8542 16882
rect 8594 16830 8596 16882
rect 8204 16660 8260 16670
rect 8540 16660 8596 16830
rect 8764 16882 8820 16894
rect 8764 16830 8766 16882
rect 8818 16830 8820 16882
rect 8764 16772 8820 16830
rect 8988 16772 9044 16782
rect 8764 16716 8932 16772
rect 8540 16604 8820 16660
rect 8204 16566 8260 16604
rect 8365 16492 8629 16502
rect 8421 16436 8469 16492
rect 8525 16436 8573 16492
rect 8092 16380 8260 16436
rect 8365 16426 8629 16436
rect 7980 15150 7982 15202
rect 8034 15150 8036 15202
rect 7980 15092 8036 15150
rect 7980 15026 8036 15036
rect 8092 15986 8148 15998
rect 8092 15934 8094 15986
rect 8146 15934 8148 15986
rect 8092 14644 8148 15934
rect 8204 15988 8260 16380
rect 8764 16324 8820 16604
rect 8540 16268 8820 16324
rect 8540 16100 8596 16268
rect 8876 16212 8932 16716
rect 8876 16146 8932 16156
rect 8540 16006 8596 16044
rect 8988 16098 9044 16716
rect 9324 16212 9380 16222
rect 8988 16046 8990 16098
rect 9042 16046 9044 16098
rect 8988 16034 9044 16046
rect 9212 16100 9268 16110
rect 8204 15922 8260 15932
rect 8764 15988 8820 15998
rect 8764 15894 8820 15932
rect 9212 15986 9268 16044
rect 9212 15934 9214 15986
rect 9266 15934 9268 15986
rect 9212 15922 9268 15934
rect 9324 15986 9380 16156
rect 9324 15934 9326 15986
rect 9378 15934 9380 15986
rect 8316 15876 8372 15886
rect 8316 15782 8372 15820
rect 8876 15874 8932 15886
rect 8876 15822 8878 15874
rect 8930 15822 8932 15874
rect 8876 15540 8932 15822
rect 8876 15484 9156 15540
rect 8092 14578 8148 14588
rect 8204 15316 8260 15326
rect 7644 14084 7700 14094
rect 7868 14084 7924 14476
rect 7700 14028 7924 14084
rect 7980 14308 8036 14318
rect 7644 13970 7700 14028
rect 7644 13918 7646 13970
rect 7698 13918 7700 13970
rect 7644 13906 7700 13918
rect 7980 13746 8036 14252
rect 7980 13694 7982 13746
rect 8034 13694 8036 13746
rect 7980 13412 8036 13694
rect 8204 13860 8260 15260
rect 8652 15204 8708 15214
rect 8988 15202 9044 15214
rect 8988 15150 8990 15202
rect 9042 15150 9044 15202
rect 8652 15092 8932 15148
rect 8365 14924 8629 14934
rect 8421 14868 8469 14924
rect 8525 14868 8573 14924
rect 8365 14858 8629 14868
rect 8428 14642 8484 14654
rect 8428 14590 8430 14642
rect 8482 14590 8484 14642
rect 8316 13860 8372 13870
rect 8204 13858 8372 13860
rect 8204 13806 8318 13858
rect 8370 13806 8372 13858
rect 8204 13804 8372 13806
rect 7980 13346 8036 13356
rect 8092 13636 8148 13646
rect 7532 13244 7924 13300
rect 7868 13188 7924 13244
rect 7868 13132 8036 13188
rect 7868 12852 7924 12862
rect 7868 12402 7924 12796
rect 7868 12350 7870 12402
rect 7922 12350 7924 12402
rect 7868 12338 7924 12350
rect 7756 12292 7812 12302
rect 7532 12290 7812 12292
rect 7532 12238 7758 12290
rect 7810 12238 7812 12290
rect 7532 12236 7812 12238
rect 7532 12178 7588 12236
rect 7756 12226 7812 12236
rect 7532 12126 7534 12178
rect 7586 12126 7588 12178
rect 7532 12114 7588 12126
rect 7980 12180 8036 13132
rect 8092 12962 8148 13580
rect 8092 12910 8094 12962
rect 8146 12910 8148 12962
rect 8092 12898 8148 12910
rect 8092 12404 8148 12414
rect 8092 12310 8148 12348
rect 8204 12292 8260 13804
rect 8316 13794 8372 13804
rect 8428 13524 8484 14590
rect 8764 14530 8820 14542
rect 8764 14478 8766 14530
rect 8818 14478 8820 14530
rect 8764 14420 8820 14478
rect 8764 14354 8820 14364
rect 8764 13972 8820 13982
rect 8876 13972 8932 15092
rect 8988 14980 9044 15150
rect 8988 14914 9044 14924
rect 8764 13970 8932 13972
rect 8764 13918 8766 13970
rect 8818 13918 8932 13970
rect 8764 13916 8932 13918
rect 8988 14756 9044 14766
rect 8764 13906 8820 13916
rect 8988 13858 9044 14700
rect 8988 13806 8990 13858
rect 9042 13806 9044 13858
rect 8988 13794 9044 13806
rect 8428 13458 8484 13468
rect 8876 13634 8932 13646
rect 8876 13582 8878 13634
rect 8930 13582 8932 13634
rect 8365 13356 8629 13366
rect 8421 13300 8469 13356
rect 8525 13300 8573 13356
rect 8365 13290 8629 13300
rect 8316 13188 8372 13198
rect 8316 12516 8372 13132
rect 8876 13076 8932 13582
rect 9100 13524 9156 15484
rect 9324 15316 9380 15934
rect 9324 15250 9380 15260
rect 9100 13458 9156 13468
rect 8876 13020 9156 13076
rect 8540 12852 8596 12862
rect 8876 12852 8932 12862
rect 8540 12850 8932 12852
rect 8540 12798 8542 12850
rect 8594 12798 8878 12850
rect 8930 12798 8932 12850
rect 8540 12796 8932 12798
rect 8540 12786 8596 12796
rect 8876 12786 8932 12796
rect 8988 12740 9044 12750
rect 8316 12460 8484 12516
rect 8316 12292 8372 12302
rect 8204 12290 8372 12292
rect 8204 12238 8318 12290
rect 8370 12238 8372 12290
rect 8204 12236 8372 12238
rect 8316 12226 8372 12236
rect 7980 12124 8148 12180
rect 7644 11732 7700 11742
rect 7644 11618 7700 11676
rect 7644 11566 7646 11618
rect 7698 11566 7700 11618
rect 7644 11554 7700 11566
rect 7980 11506 8036 11518
rect 7980 11454 7982 11506
rect 8034 11454 8036 11506
rect 7868 11284 7924 11294
rect 7868 11190 7924 11228
rect 7756 11060 7812 11070
rect 7420 10558 7422 10610
rect 7474 10558 7476 10610
rect 7420 10546 7476 10558
rect 7644 10724 7700 10734
rect 7308 10332 7588 10388
rect 6972 9202 7028 9212
rect 7532 9154 7588 10332
rect 7532 9102 7534 9154
rect 7586 9102 7588 9154
rect 7532 9090 7588 9102
rect 7644 9044 7700 10668
rect 7644 8950 7700 8988
rect 7756 8820 7812 11004
rect 7868 10836 7924 10846
rect 7868 10722 7924 10780
rect 7868 10670 7870 10722
rect 7922 10670 7924 10722
rect 7868 10658 7924 10670
rect 7980 9826 8036 11454
rect 7980 9774 7982 9826
rect 8034 9774 8036 9826
rect 7980 9762 8036 9774
rect 8092 9604 8148 12124
rect 8428 12068 8484 12460
rect 8204 12012 8484 12068
rect 8204 10836 8260 12012
rect 8365 11788 8629 11798
rect 8421 11732 8469 11788
rect 8525 11732 8573 11788
rect 8365 11722 8629 11732
rect 8988 11620 9044 12684
rect 9100 12404 9156 13020
rect 9212 12852 9268 12862
rect 9212 12758 9268 12796
rect 9100 12348 9268 12404
rect 9100 12066 9156 12078
rect 9100 12014 9102 12066
rect 9154 12014 9156 12066
rect 9100 11956 9156 12014
rect 9100 11890 9156 11900
rect 8988 11564 9156 11620
rect 8316 11394 8372 11406
rect 8316 11342 8318 11394
rect 8370 11342 8372 11394
rect 8316 11060 8372 11342
rect 8652 11282 8708 11294
rect 8652 11230 8654 11282
rect 8706 11230 8708 11282
rect 8316 10994 8372 11004
rect 8540 11170 8596 11182
rect 8540 11118 8542 11170
rect 8594 11118 8596 11170
rect 8204 10770 8260 10780
rect 8316 10724 8372 10734
rect 8316 10610 8372 10668
rect 8316 10558 8318 10610
rect 8370 10558 8372 10610
rect 8316 10546 8372 10558
rect 8540 10388 8596 11118
rect 8652 10612 8708 11230
rect 8988 11172 9044 11182
rect 8652 10546 8708 10556
rect 8876 11170 9044 11172
rect 8876 11118 8990 11170
rect 9042 11118 9044 11170
rect 8876 11116 9044 11118
rect 8540 10332 8820 10388
rect 8365 10220 8629 10230
rect 8421 10164 8469 10220
rect 8525 10164 8573 10220
rect 8365 10154 8629 10164
rect 8764 10052 8820 10332
rect 8764 9986 8820 9996
rect 6188 8206 6190 8258
rect 6242 8206 6244 8258
rect 5740 8036 5796 8046
rect 5740 7942 5796 7980
rect 5404 7474 5460 7486
rect 5404 7422 5406 7474
rect 5458 7422 5460 7474
rect 5404 7252 5460 7422
rect 5628 7474 5684 7644
rect 5628 7422 5630 7474
rect 5682 7422 5684 7474
rect 5628 7410 5684 7422
rect 5964 7476 6020 7486
rect 5964 7382 6020 7420
rect 6188 7474 6244 8206
rect 7532 8764 7812 8820
rect 7980 9548 8148 9604
rect 8764 9602 8820 9614
rect 8764 9550 8766 9602
rect 8818 9550 8820 9602
rect 7196 8146 7252 8158
rect 7196 8094 7198 8146
rect 7250 8094 7252 8146
rect 6636 7700 6692 7710
rect 6636 7606 6692 7644
rect 7196 7700 7252 8094
rect 7196 7634 7252 7644
rect 6188 7422 6190 7474
rect 6242 7422 6244 7474
rect 6188 7410 6244 7422
rect 6860 7474 6916 7486
rect 6860 7422 6862 7474
rect 6914 7422 6916 7474
rect 5516 7364 5572 7374
rect 5516 7270 5572 7308
rect 6748 7364 6804 7374
rect 6748 7270 6804 7308
rect 5404 7186 5460 7196
rect 6860 7252 6916 7422
rect 7196 7476 7252 7486
rect 7196 7382 7252 7420
rect 7308 7364 7364 7374
rect 7308 7270 7364 7308
rect 6860 7186 6916 7196
rect 5292 6972 5572 7028
rect 4732 6802 4900 6804
rect 4732 6750 4734 6802
rect 4786 6750 4900 6802
rect 4732 6748 4900 6750
rect 4732 6738 4788 6748
rect 4956 6692 5012 6702
rect 4620 6300 4900 6356
rect 4620 6018 4676 6300
rect 4620 5966 4622 6018
rect 4674 5966 4676 6018
rect 4620 5954 4676 5966
rect 4732 6130 4788 6142
rect 4732 6078 4734 6130
rect 4786 6078 4788 6130
rect 3612 5908 3668 5918
rect 3612 5814 3668 5852
rect 3500 5182 3502 5234
rect 3554 5182 3556 5234
rect 3500 5170 3556 5182
rect 3948 5236 4004 5246
rect 3948 4900 4004 5180
rect 4396 4900 4452 4910
rect 3948 4898 4452 4900
rect 3948 4846 3950 4898
rect 4002 4846 4398 4898
rect 4450 4846 4452 4898
rect 3948 4844 4452 4846
rect 3948 4834 4004 4844
rect 4396 4338 4452 4844
rect 4396 4286 4398 4338
rect 4450 4286 4452 4338
rect 4396 3668 4452 4286
rect 4396 3602 4452 3612
rect 2940 3390 2942 3442
rect 2994 3390 2996 3442
rect 2940 3378 2996 3390
rect 3164 3554 3220 3566
rect 3164 3502 3166 3554
rect 3218 3502 3220 3554
rect 3164 3220 3220 3502
rect 4732 3554 4788 6078
rect 4844 5010 4900 6300
rect 4956 5234 5012 6636
rect 5292 6132 5348 6142
rect 5292 6038 5348 6076
rect 5516 5906 5572 6972
rect 6412 6802 6468 6814
rect 6412 6750 6414 6802
rect 6466 6750 6468 6802
rect 5740 6692 5796 6702
rect 5740 6598 5796 6636
rect 6300 6690 6356 6702
rect 6300 6638 6302 6690
rect 6354 6638 6356 6690
rect 6188 6580 6244 6590
rect 6076 6524 6188 6580
rect 5516 5854 5518 5906
rect 5570 5854 5572 5906
rect 5516 5842 5572 5854
rect 5964 6132 6020 6142
rect 5964 5906 6020 6076
rect 5964 5854 5966 5906
rect 6018 5854 6020 5906
rect 5964 5842 6020 5854
rect 5964 5684 6020 5694
rect 5068 5682 6020 5684
rect 5068 5630 5966 5682
rect 6018 5630 6020 5682
rect 5068 5628 6020 5630
rect 5068 5346 5124 5628
rect 5964 5618 6020 5628
rect 6076 5460 6132 6524
rect 6188 6514 6244 6524
rect 6300 5908 6356 6638
rect 6300 5814 6356 5852
rect 5068 5294 5070 5346
rect 5122 5294 5124 5346
rect 5068 5282 5124 5294
rect 5852 5404 6132 5460
rect 4956 5182 4958 5234
rect 5010 5182 5012 5234
rect 4956 5170 5012 5182
rect 5852 5234 5908 5404
rect 6412 5348 6468 6750
rect 7532 6690 7588 8764
rect 7532 6638 7534 6690
rect 7586 6638 7588 6690
rect 7532 6626 7588 6638
rect 7756 8370 7812 8382
rect 7756 8318 7758 8370
rect 7810 8318 7812 8370
rect 7756 7362 7812 8318
rect 7756 7310 7758 7362
rect 7810 7310 7812 7362
rect 7756 7252 7812 7310
rect 6524 6578 6580 6590
rect 6524 6526 6526 6578
rect 6578 6526 6580 6578
rect 6524 6132 6580 6526
rect 6580 6076 6692 6132
rect 6524 6066 6580 6076
rect 6636 6018 6692 6076
rect 6636 5966 6638 6018
rect 6690 5966 6692 6018
rect 6636 5954 6692 5966
rect 6748 6020 6804 6030
rect 6636 5348 6692 5358
rect 6412 5292 6636 5348
rect 5852 5182 5854 5234
rect 5906 5182 5908 5234
rect 5852 5170 5908 5182
rect 6636 5122 6692 5292
rect 6636 5070 6638 5122
rect 6690 5070 6692 5122
rect 6636 5058 6692 5070
rect 4844 4958 4846 5010
rect 4898 4958 4900 5010
rect 4844 4946 4900 4958
rect 6412 4900 6468 4910
rect 6412 4806 6468 4844
rect 5068 4228 5124 4238
rect 4732 3502 4734 3554
rect 4786 3502 4788 3554
rect 4732 3490 4788 3502
rect 4956 4226 5124 4228
rect 4956 4174 5070 4226
rect 5122 4174 5124 4226
rect 4956 4172 5124 4174
rect 4956 3442 5012 4172
rect 5068 4162 5124 4172
rect 6300 3668 6356 3678
rect 6300 3574 6356 3612
rect 6748 3666 6804 5964
rect 7756 5906 7812 7196
rect 7868 6690 7924 6702
rect 7868 6638 7870 6690
rect 7922 6638 7924 6690
rect 7868 6132 7924 6638
rect 7868 6066 7924 6076
rect 7756 5854 7758 5906
rect 7810 5854 7812 5906
rect 7756 5842 7812 5854
rect 7868 5236 7924 5246
rect 7868 5010 7924 5180
rect 7868 4958 7870 5010
rect 7922 4958 7924 5010
rect 7868 4946 7924 4958
rect 7644 4340 7700 4350
rect 7196 4338 7700 4340
rect 7196 4286 7646 4338
rect 7698 4286 7700 4338
rect 7196 4284 7700 4286
rect 7196 4226 7252 4284
rect 7644 4274 7700 4284
rect 7196 4174 7198 4226
rect 7250 4174 7252 4226
rect 7196 4162 7252 4174
rect 7756 4114 7812 4126
rect 7756 4062 7758 4114
rect 7810 4062 7812 4114
rect 7644 3780 7700 3790
rect 6748 3614 6750 3666
rect 6802 3614 6804 3666
rect 6748 3602 6804 3614
rect 7196 3668 7252 3678
rect 7196 3574 7252 3612
rect 7644 3666 7700 3724
rect 7644 3614 7646 3666
rect 7698 3614 7700 3666
rect 7644 3602 7700 3614
rect 4956 3390 4958 3442
rect 5010 3390 5012 3442
rect 4956 3378 5012 3390
rect 5852 3444 5908 3482
rect 5852 3378 5908 3388
rect 7756 3332 7812 4062
rect 7868 3444 7924 3454
rect 7980 3444 8036 9548
rect 8204 9380 8260 9390
rect 8092 9324 8204 9380
rect 8092 7476 8148 9324
rect 8204 9314 8260 9324
rect 8204 8820 8260 8830
rect 8204 8726 8260 8764
rect 8540 8820 8596 8858
rect 8540 8754 8596 8764
rect 8365 8652 8629 8662
rect 8421 8596 8469 8652
rect 8525 8596 8573 8652
rect 8365 8586 8629 8596
rect 8764 8260 8820 9550
rect 8652 8204 8820 8260
rect 8204 7476 8260 7486
rect 8092 7474 8260 7476
rect 8092 7422 8206 7474
rect 8258 7422 8260 7474
rect 8092 7420 8260 7422
rect 8204 7410 8260 7420
rect 8652 7364 8708 8204
rect 8764 8036 8820 8046
rect 8764 7942 8820 7980
rect 8652 7298 8708 7308
rect 8316 7252 8372 7262
rect 8204 7196 8316 7252
rect 8204 6130 8260 7196
rect 8316 7186 8372 7196
rect 8365 7084 8629 7094
rect 8421 7028 8469 7084
rect 8525 7028 8573 7084
rect 8365 7018 8629 7028
rect 8540 6692 8596 6702
rect 8876 6692 8932 11116
rect 8988 11106 9044 11116
rect 9100 11060 9156 11564
rect 9212 11618 9268 12348
rect 9436 12292 9492 17164
rect 9548 16996 9604 17006
rect 9548 16902 9604 16940
rect 9548 16660 9604 16670
rect 9548 15204 9604 16604
rect 9660 16212 9716 17614
rect 9772 17556 9828 18174
rect 9772 17490 9828 17500
rect 9772 16772 9828 16782
rect 9772 16678 9828 16716
rect 9884 16660 9940 18844
rect 9996 17668 10052 19068
rect 10332 19122 10388 19134
rect 10332 19070 10334 19122
rect 10386 19070 10388 19122
rect 10220 18450 10276 18462
rect 10220 18398 10222 18450
rect 10274 18398 10276 18450
rect 10220 17780 10276 18398
rect 10332 18452 10388 19070
rect 10444 19124 10500 19292
rect 10444 19030 10500 19068
rect 10332 17890 10388 18396
rect 10556 18452 10612 19854
rect 10668 19234 10724 19964
rect 10780 19926 10836 19964
rect 10668 19182 10670 19234
rect 10722 19182 10724 19234
rect 10668 19170 10724 19182
rect 10780 19572 10836 19582
rect 10332 17838 10334 17890
rect 10386 17838 10388 17890
rect 10332 17826 10388 17838
rect 10444 18116 10500 18126
rect 10220 17714 10276 17724
rect 10108 17668 10164 17678
rect 9996 17666 10164 17668
rect 9996 17614 10110 17666
rect 10162 17614 10164 17666
rect 9996 17612 10164 17614
rect 10108 17108 10164 17612
rect 10108 17042 10164 17052
rect 9884 16594 9940 16604
rect 10108 16658 10164 16670
rect 10108 16606 10110 16658
rect 10162 16606 10164 16658
rect 9772 16212 9828 16222
rect 9660 16210 10052 16212
rect 9660 16158 9774 16210
rect 9826 16158 10052 16210
rect 9660 16156 10052 16158
rect 9772 16146 9828 16156
rect 9884 15426 9940 15438
rect 9884 15374 9886 15426
rect 9938 15374 9940 15426
rect 9548 15138 9604 15148
rect 9772 15316 9828 15326
rect 9772 15092 9828 15260
rect 9772 15026 9828 15036
rect 9884 14756 9940 15374
rect 9996 15148 10052 16156
rect 10108 15428 10164 16606
rect 10220 15874 10276 15886
rect 10220 15822 10222 15874
rect 10274 15822 10276 15874
rect 10220 15652 10276 15822
rect 10220 15586 10276 15596
rect 10108 15314 10164 15372
rect 10108 15262 10110 15314
rect 10162 15262 10164 15314
rect 10108 15250 10164 15262
rect 9996 15092 10164 15148
rect 9884 14690 9940 14700
rect 9884 14532 9940 14542
rect 9884 14438 9940 14476
rect 10108 14308 10164 15092
rect 10108 14242 10164 14252
rect 10220 14532 10276 14542
rect 9548 13748 9604 13758
rect 9548 13654 9604 13692
rect 10108 13636 10164 13646
rect 10108 13542 10164 13580
rect 9772 13524 9828 13534
rect 9772 13430 9828 13468
rect 9548 13074 9604 13086
rect 9548 13022 9550 13074
rect 9602 13022 9604 13074
rect 9548 12516 9604 13022
rect 9548 12450 9604 12460
rect 9548 12292 9604 12302
rect 9436 12290 9604 12292
rect 9436 12238 9550 12290
rect 9602 12238 9604 12290
rect 9436 12236 9604 12238
rect 9548 12226 9604 12236
rect 9884 12290 9940 12302
rect 9884 12238 9886 12290
rect 9938 12238 9940 12290
rect 9212 11566 9214 11618
rect 9266 11566 9268 11618
rect 9212 11554 9268 11566
rect 9212 11396 9268 11406
rect 9436 11396 9492 11406
rect 9212 11302 9268 11340
rect 9324 11394 9492 11396
rect 9324 11342 9438 11394
rect 9490 11342 9492 11394
rect 9324 11340 9492 11342
rect 9100 11004 9268 11060
rect 8988 10612 9044 10622
rect 9044 10556 9156 10612
rect 8988 10518 9044 10556
rect 8988 9156 9044 9166
rect 8988 8258 9044 9100
rect 8988 8206 8990 8258
rect 9042 8206 9044 8258
rect 8988 8194 9044 8206
rect 9100 7588 9156 10556
rect 8540 6690 8932 6692
rect 8540 6638 8542 6690
rect 8594 6638 8932 6690
rect 8540 6636 8932 6638
rect 8988 7532 9156 7588
rect 8540 6626 8596 6636
rect 8988 6580 9044 7532
rect 9100 7364 9156 7374
rect 9212 7364 9268 11004
rect 9100 7362 9268 7364
rect 9100 7310 9102 7362
rect 9154 7310 9268 7362
rect 9100 7308 9268 7310
rect 9100 7298 9156 7308
rect 9324 7028 9380 11340
rect 9436 11330 9492 11340
rect 9884 11396 9940 12238
rect 10220 11396 10276 14476
rect 10444 13860 10500 18060
rect 10556 17890 10612 18396
rect 10556 17838 10558 17890
rect 10610 17838 10612 17890
rect 10556 16772 10612 17838
rect 10556 15986 10612 16716
rect 10668 18340 10724 18350
rect 10780 18340 10836 19516
rect 10668 18338 10836 18340
rect 10668 18286 10670 18338
rect 10722 18286 10836 18338
rect 10668 18284 10836 18286
rect 10668 17668 10724 18284
rect 10892 18116 10948 20188
rect 11116 20132 11172 21644
rect 11228 21474 11284 21486
rect 11228 21422 11230 21474
rect 11282 21422 11284 21474
rect 11228 20578 11284 21422
rect 11452 20916 11508 20926
rect 11340 20804 11396 20814
rect 11340 20710 11396 20748
rect 11452 20802 11508 20860
rect 11452 20750 11454 20802
rect 11506 20750 11508 20802
rect 11452 20738 11508 20750
rect 11228 20526 11230 20578
rect 11282 20526 11284 20578
rect 11228 20514 11284 20526
rect 11676 20468 11732 22316
rect 12124 20692 12180 23660
rect 12236 23714 12292 23726
rect 12236 23662 12238 23714
rect 12290 23662 12292 23714
rect 12236 23268 12292 23662
rect 12572 23548 12628 23772
rect 12236 23202 12292 23212
rect 12348 23492 12628 23548
rect 12348 22372 12404 23492
rect 12796 23156 12852 25228
rect 12796 23090 12852 23100
rect 12684 23044 12740 23054
rect 12684 22950 12740 22988
rect 12236 22316 12404 22372
rect 13020 22372 13076 22382
rect 12236 20916 12292 22316
rect 13020 22278 13076 22316
rect 12684 22260 12740 22270
rect 12684 22166 12740 22204
rect 12348 22146 12404 22158
rect 12348 22094 12350 22146
rect 12402 22094 12404 22146
rect 12348 22036 12404 22094
rect 12796 22146 12852 22158
rect 12796 22094 12798 22146
rect 12850 22094 12852 22146
rect 12796 22036 12852 22094
rect 12348 21980 12852 22036
rect 12236 20860 12404 20916
rect 12236 20692 12292 20702
rect 12124 20690 12292 20692
rect 12124 20638 12238 20690
rect 12290 20638 12292 20690
rect 12124 20636 12292 20638
rect 12236 20626 12292 20636
rect 11116 20066 11172 20076
rect 11564 20412 11732 20468
rect 11900 20578 11956 20590
rect 11900 20526 11902 20578
rect 11954 20526 11956 20578
rect 11452 20020 11508 20030
rect 11452 19926 11508 19964
rect 11116 19908 11172 19918
rect 11116 19814 11172 19852
rect 11452 19460 11508 19470
rect 11564 19460 11620 20412
rect 11452 19458 11620 19460
rect 11452 19406 11454 19458
rect 11506 19406 11620 19458
rect 11452 19404 11620 19406
rect 11676 20130 11732 20142
rect 11676 20078 11678 20130
rect 11730 20078 11732 20130
rect 11452 19394 11508 19404
rect 11676 19348 11732 20078
rect 11788 20132 11844 20142
rect 11788 19906 11844 20076
rect 11788 19854 11790 19906
rect 11842 19854 11844 19906
rect 11788 19842 11844 19854
rect 11900 19908 11956 20526
rect 11900 19842 11956 19852
rect 12124 20356 12180 20366
rect 11676 19346 11956 19348
rect 11676 19294 11678 19346
rect 11730 19294 11956 19346
rect 11676 19292 11956 19294
rect 11676 19282 11732 19292
rect 11116 19234 11172 19246
rect 11116 19182 11118 19234
rect 11170 19182 11172 19234
rect 11116 18228 11172 19182
rect 11564 19234 11620 19246
rect 11564 19182 11566 19234
rect 11618 19182 11620 19234
rect 11452 19124 11508 19134
rect 11564 19124 11620 19182
rect 11340 19068 11452 19124
rect 11508 19068 11620 19124
rect 11228 18452 11284 18462
rect 11340 18452 11396 19068
rect 11452 19058 11508 19068
rect 11228 18450 11396 18452
rect 11228 18398 11230 18450
rect 11282 18398 11396 18450
rect 11228 18396 11396 18398
rect 11452 18452 11508 18462
rect 11676 18452 11732 18462
rect 11508 18450 11732 18452
rect 11508 18398 11678 18450
rect 11730 18398 11732 18450
rect 11508 18396 11732 18398
rect 11228 18386 11284 18396
rect 11452 18386 11508 18396
rect 11676 18386 11732 18396
rect 11452 18228 11508 18238
rect 11116 18226 11508 18228
rect 11116 18174 11454 18226
rect 11506 18174 11508 18226
rect 11116 18172 11508 18174
rect 10892 18050 10948 18060
rect 10668 16324 10724 17612
rect 11452 17668 11508 18172
rect 11900 18004 11956 19292
rect 12124 18674 12180 20300
rect 12124 18622 12126 18674
rect 12178 18622 12180 18674
rect 12124 18610 12180 18622
rect 11452 17602 11508 17612
rect 11564 17948 11956 18004
rect 12348 18004 12404 20860
rect 12684 20578 12740 20590
rect 12684 20526 12686 20578
rect 12738 20526 12740 20578
rect 12572 20132 12628 20142
rect 12460 20018 12516 20030
rect 12460 19966 12462 20018
rect 12514 19966 12516 20018
rect 12460 19908 12516 19966
rect 12460 19842 12516 19852
rect 12572 19234 12628 20076
rect 12572 19182 12574 19234
rect 12626 19182 12628 19234
rect 12572 19170 12628 19182
rect 12684 19236 12740 20526
rect 12796 19348 12852 21980
rect 12796 19282 12852 19292
rect 12908 19906 12964 19918
rect 12908 19854 12910 19906
rect 12962 19854 12964 19906
rect 12684 18450 12740 19180
rect 12796 19124 12852 19134
rect 12796 19030 12852 19068
rect 12908 18564 12964 19854
rect 12908 18498 12964 18508
rect 13020 18562 13076 18574
rect 13020 18510 13022 18562
rect 13074 18510 13076 18562
rect 12684 18398 12686 18450
rect 12738 18398 12740 18450
rect 12684 18228 12740 18398
rect 12684 18162 12740 18172
rect 12908 18116 12964 18126
rect 12348 17948 12852 18004
rect 11004 17444 11060 17454
rect 11004 17350 11060 17388
rect 10668 16258 10724 16268
rect 10780 17164 11508 17220
rect 10780 16100 10836 17164
rect 11452 17106 11508 17164
rect 11452 17054 11454 17106
rect 11506 17054 11508 17106
rect 11452 17042 11508 17054
rect 10892 16996 10948 17006
rect 10892 16902 10948 16940
rect 11564 16884 11620 17948
rect 11788 17780 11844 17790
rect 11788 17666 11844 17724
rect 11900 17780 11956 17948
rect 12572 17780 12628 17790
rect 11900 17778 12068 17780
rect 11900 17726 11902 17778
rect 11954 17726 12068 17778
rect 11900 17724 12068 17726
rect 11900 17714 11956 17724
rect 11788 17614 11790 17666
rect 11842 17614 11844 17666
rect 11788 17556 11844 17614
rect 11788 17500 11956 17556
rect 11116 16828 11620 16884
rect 11004 16770 11060 16782
rect 11004 16718 11006 16770
rect 11058 16718 11060 16770
rect 11004 16212 11060 16718
rect 11116 16770 11172 16828
rect 11116 16718 11118 16770
rect 11170 16718 11172 16770
rect 11116 16706 11172 16718
rect 11004 16156 11396 16212
rect 11340 16100 11396 16156
rect 10780 16098 10948 16100
rect 10780 16046 10782 16098
rect 10834 16046 10948 16098
rect 10780 16044 10948 16046
rect 10780 16034 10836 16044
rect 10556 15934 10558 15986
rect 10610 15934 10612 15986
rect 10556 15922 10612 15934
rect 10668 15988 10724 15998
rect 10556 15426 10612 15438
rect 10556 15374 10558 15426
rect 10610 15374 10612 15426
rect 10556 14868 10612 15374
rect 10668 15204 10724 15932
rect 10780 15428 10836 15438
rect 10780 15314 10836 15372
rect 10780 15262 10782 15314
rect 10834 15262 10836 15314
rect 10780 15250 10836 15262
rect 10668 15092 10836 15148
rect 10556 14802 10612 14812
rect 10668 14532 10724 14542
rect 10668 14438 10724 14476
rect 10780 14418 10836 15092
rect 10780 14366 10782 14418
rect 10834 14366 10836 14418
rect 10780 14354 10836 14366
rect 10556 13860 10612 13870
rect 10444 13804 10556 13860
rect 10556 13746 10612 13804
rect 10556 13694 10558 13746
rect 10610 13694 10612 13746
rect 10556 13682 10612 13694
rect 10892 13748 10948 16044
rect 11340 16006 11396 16044
rect 11452 15876 11508 15886
rect 11340 15820 11452 15876
rect 11228 14756 11284 14766
rect 11228 14530 11284 14700
rect 11340 14644 11396 15820
rect 11452 15782 11508 15820
rect 11676 15874 11732 15886
rect 11676 15822 11678 15874
rect 11730 15822 11732 15874
rect 11452 15540 11508 15550
rect 11452 15446 11508 15484
rect 11676 15316 11732 15822
rect 11676 15260 11844 15316
rect 11564 15204 11620 15214
rect 11676 15148 11732 15158
rect 11564 15146 11732 15148
rect 11564 15094 11678 15146
rect 11730 15094 11732 15146
rect 11564 15092 11732 15094
rect 11676 15082 11732 15092
rect 11340 14588 11508 14644
rect 11228 14478 11230 14530
rect 11282 14478 11284 14530
rect 11004 14420 11060 14430
rect 11004 14326 11060 14364
rect 10892 13692 11060 13748
rect 10668 13634 10724 13646
rect 10668 13582 10670 13634
rect 10722 13582 10724 13634
rect 10444 12290 10500 12302
rect 10444 12238 10446 12290
rect 10498 12238 10500 12290
rect 10444 11620 10500 12238
rect 10444 11554 10500 11564
rect 10668 11618 10724 13582
rect 10892 13524 10948 13534
rect 10780 13468 10892 13524
rect 10780 12402 10836 13468
rect 10892 13430 10948 13468
rect 10780 12350 10782 12402
rect 10834 12350 10836 12402
rect 10780 12338 10836 12350
rect 10892 12740 10948 12750
rect 10668 11566 10670 11618
rect 10722 11566 10724 11618
rect 10668 11554 10724 11566
rect 9884 11330 9940 11340
rect 9996 11394 10276 11396
rect 9996 11342 10222 11394
rect 10274 11342 10276 11394
rect 9996 11340 10276 11342
rect 9772 11282 9828 11294
rect 9772 11230 9774 11282
rect 9826 11230 9828 11282
rect 9772 11172 9828 11230
rect 9996 11172 10052 11340
rect 10220 11330 10276 11340
rect 10556 11396 10612 11406
rect 10556 11394 10836 11396
rect 10556 11342 10558 11394
rect 10610 11342 10836 11394
rect 10556 11340 10836 11342
rect 10556 11330 10612 11340
rect 9772 11116 10052 11172
rect 10332 11170 10388 11182
rect 10332 11118 10334 11170
rect 10386 11118 10388 11170
rect 9884 10612 9940 10622
rect 9772 10610 9940 10612
rect 9772 10558 9886 10610
rect 9938 10558 9940 10610
rect 9772 10556 9940 10558
rect 9772 9940 9828 10556
rect 9884 10546 9940 10556
rect 9996 10500 10052 10510
rect 9996 10164 10052 10444
rect 9772 9874 9828 9884
rect 9884 10108 10052 10164
rect 10108 10386 10164 10398
rect 10108 10334 10110 10386
rect 10162 10334 10164 10386
rect 9660 9826 9716 9838
rect 9660 9774 9662 9826
rect 9714 9774 9716 9826
rect 9436 9716 9492 9726
rect 9436 9622 9492 9660
rect 9548 9604 9604 9614
rect 9548 9042 9604 9548
rect 9660 9380 9716 9774
rect 9660 9314 9716 9324
rect 9772 9604 9828 9614
rect 9548 8990 9550 9042
rect 9602 8990 9604 9042
rect 9548 8978 9604 8990
rect 9660 8932 9716 8942
rect 9660 8838 9716 8876
rect 9772 8370 9828 9548
rect 9884 9154 9940 10108
rect 10108 9828 10164 10334
rect 9884 9102 9886 9154
rect 9938 9102 9940 9154
rect 9884 9090 9940 9102
rect 9996 9772 10164 9828
rect 10220 9828 10276 9838
rect 9996 8932 10052 9772
rect 10220 9268 10276 9772
rect 10220 9202 10276 9212
rect 10220 9044 10276 9054
rect 9996 8866 10052 8876
rect 10108 9042 10276 9044
rect 10108 8990 10222 9042
rect 10274 8990 10276 9042
rect 10108 8988 10276 8990
rect 10108 8484 10164 8988
rect 10220 8978 10276 8988
rect 9772 8318 9774 8370
rect 9826 8318 9828 8370
rect 9772 8306 9828 8318
rect 9884 8428 10164 8484
rect 10220 8820 10276 8830
rect 8988 6514 9044 6524
rect 9100 6972 9380 7028
rect 9660 7476 9716 7486
rect 9884 7476 9940 8428
rect 9660 7474 9940 7476
rect 9660 7422 9662 7474
rect 9714 7422 9940 7474
rect 9660 7420 9940 7422
rect 8204 6078 8206 6130
rect 8258 6078 8260 6130
rect 8204 6066 8260 6078
rect 8988 6132 9044 6142
rect 8988 6038 9044 6076
rect 8652 6020 8708 6030
rect 8652 5926 8708 5964
rect 8876 5572 8932 5582
rect 8365 5516 8629 5526
rect 8421 5460 8469 5516
rect 8525 5460 8573 5516
rect 8365 5450 8629 5460
rect 8204 5234 8260 5246
rect 8204 5182 8206 5234
rect 8258 5182 8260 5234
rect 8204 5124 8260 5182
rect 8876 5234 8932 5516
rect 9100 5348 9156 6972
rect 9660 6132 9716 7420
rect 9660 6066 9716 6076
rect 9772 6132 9828 6142
rect 10220 6132 10276 8764
rect 10332 7586 10388 11118
rect 10444 10610 10500 10622
rect 10444 10558 10446 10610
rect 10498 10558 10500 10610
rect 10444 9940 10500 10558
rect 10668 10610 10724 10622
rect 10668 10558 10670 10610
rect 10722 10558 10724 10610
rect 10444 9874 10500 9884
rect 10556 10498 10612 10510
rect 10556 10446 10558 10498
rect 10610 10446 10612 10498
rect 10556 9716 10612 10446
rect 10668 10500 10724 10558
rect 10668 10434 10724 10444
rect 10668 9828 10724 9866
rect 10668 9762 10724 9772
rect 10556 9650 10612 9660
rect 10668 9604 10724 9614
rect 10668 9510 10724 9548
rect 10332 7534 10334 7586
rect 10386 7534 10388 7586
rect 10332 7522 10388 7534
rect 10780 8036 10836 11340
rect 10892 11394 10948 12684
rect 10892 11342 10894 11394
rect 10946 11342 10948 11394
rect 10892 11330 10948 11342
rect 11004 10724 11060 13692
rect 11228 13524 11284 14478
rect 11228 13458 11284 13468
rect 11340 14308 11396 14318
rect 11228 13188 11284 13198
rect 11228 12740 11284 13132
rect 11228 12402 11284 12684
rect 11228 12350 11230 12402
rect 11282 12350 11284 12402
rect 11228 12338 11284 12350
rect 11340 11396 11396 14252
rect 11452 13636 11508 14588
rect 11564 14532 11620 14542
rect 11564 14306 11620 14476
rect 11788 14532 11844 15260
rect 11788 14466 11844 14476
rect 11564 14254 11566 14306
rect 11618 14254 11620 14306
rect 11564 13860 11620 14254
rect 11564 13794 11620 13804
rect 11788 13858 11844 13870
rect 11788 13806 11790 13858
rect 11842 13806 11844 13858
rect 11564 13636 11620 13646
rect 11452 13580 11564 13636
rect 11564 13542 11620 13580
rect 11676 12852 11732 12862
rect 11676 12758 11732 12796
rect 11564 12180 11620 12190
rect 11788 12180 11844 13806
rect 11900 12404 11956 17500
rect 12012 16882 12068 17724
rect 12012 16830 12014 16882
rect 12066 16830 12068 16882
rect 12012 16818 12068 16830
rect 12124 17668 12180 17678
rect 12012 16098 12068 16110
rect 12012 16046 12014 16098
rect 12066 16046 12068 16098
rect 12012 15148 12068 16046
rect 12124 15652 12180 17612
rect 12572 17666 12628 17724
rect 12572 17614 12574 17666
rect 12626 17614 12628 17666
rect 12572 16996 12628 17614
rect 12796 17106 12852 17948
rect 12908 17778 12964 18060
rect 13020 17892 13076 18510
rect 13244 18452 13300 29036
rect 13356 25732 13412 29372
rect 13468 26628 13524 31892
rect 13692 29986 13748 29998
rect 13692 29934 13694 29986
rect 13746 29934 13748 29986
rect 13580 29428 13636 29438
rect 13692 29428 13748 29934
rect 13804 29652 13860 29662
rect 13804 29558 13860 29596
rect 13580 29426 13748 29428
rect 13580 29374 13582 29426
rect 13634 29374 13748 29426
rect 13580 29372 13748 29374
rect 13580 29204 13636 29372
rect 13580 29138 13636 29148
rect 13916 28644 13972 31892
rect 14252 31780 14308 31790
rect 14252 31686 14308 31724
rect 14812 31778 14868 31790
rect 14812 31726 14814 31778
rect 14866 31726 14868 31778
rect 14812 31220 14868 31726
rect 14812 31154 14868 31164
rect 14924 31108 14980 33406
rect 15708 33458 15764 34076
rect 16268 34066 16324 34076
rect 15708 33406 15710 33458
rect 15762 33406 15764 33458
rect 15708 33394 15764 33406
rect 16716 33460 16772 34188
rect 16828 33460 16884 33470
rect 16716 33458 16884 33460
rect 16716 33406 16830 33458
rect 16882 33406 16884 33458
rect 16716 33404 16884 33406
rect 16828 33394 16884 33404
rect 15260 33346 15316 33358
rect 15260 33294 15262 33346
rect 15314 33294 15316 33346
rect 15260 32786 15316 33294
rect 16156 33346 16212 33358
rect 16156 33294 16158 33346
rect 16210 33294 16212 33346
rect 15518 32956 15782 32966
rect 15574 32900 15622 32956
rect 15678 32900 15726 32956
rect 15518 32890 15782 32900
rect 16156 32900 16212 33294
rect 16156 32834 16212 32844
rect 16828 32900 16884 32910
rect 15260 32734 15262 32786
rect 15314 32734 15316 32786
rect 15260 32722 15316 32734
rect 16156 32676 16212 32686
rect 16212 32620 16324 32676
rect 16156 32582 16212 32620
rect 15148 32562 15204 32574
rect 15148 32510 15150 32562
rect 15202 32510 15204 32562
rect 15148 32452 15204 32510
rect 15148 32386 15204 32396
rect 15372 32564 15428 32574
rect 15372 32340 15428 32508
rect 15820 32564 15876 32574
rect 15820 32562 15988 32564
rect 15820 32510 15822 32562
rect 15874 32510 15988 32562
rect 15820 32508 15988 32510
rect 15820 32498 15876 32508
rect 15372 32274 15428 32284
rect 15820 32340 15876 32350
rect 15596 32116 15652 32126
rect 15148 31780 15204 31790
rect 15148 31778 15428 31780
rect 15148 31726 15150 31778
rect 15202 31726 15428 31778
rect 15148 31724 15428 31726
rect 15148 31714 15204 31724
rect 14924 31042 14980 31052
rect 15372 31220 15428 31724
rect 15596 31666 15652 32060
rect 15820 31780 15876 32284
rect 15932 31892 15988 32508
rect 16044 32452 16100 32462
rect 16044 32358 16100 32396
rect 16268 32116 16324 32620
rect 16828 32452 16884 32844
rect 17724 32786 17780 34748
rect 17836 34692 17892 35534
rect 17836 34354 17892 34636
rect 17836 34302 17838 34354
rect 17890 34302 17892 34354
rect 17836 34290 17892 34302
rect 17724 32734 17726 32786
rect 17778 32734 17780 32786
rect 17724 32722 17780 32734
rect 18060 32788 18116 36540
rect 19292 36594 19348 39228
rect 20832 39200 20944 40000
rect 21196 39228 21588 39284
rect 20860 39060 20916 39200
rect 21196 39060 21252 39228
rect 20860 39004 21252 39060
rect 19292 36542 19294 36594
rect 19346 36542 19348 36594
rect 19292 36530 19348 36542
rect 21532 36594 21588 39228
rect 23072 39200 23184 40000
rect 25312 39200 25424 40000
rect 27552 39200 27664 40000
rect 29792 39200 29904 40000
rect 32032 39200 32144 40000
rect 34272 39200 34384 40000
rect 36512 39200 36624 40000
rect 38752 39200 38864 40000
rect 40992 39200 41104 40000
rect 43232 39200 43344 40000
rect 45472 39200 45584 40000
rect 47712 39200 47824 40000
rect 49952 39200 50064 40000
rect 52192 39200 52304 40000
rect 54432 39200 54544 40000
rect 56672 39200 56784 40000
rect 22672 36876 22936 36886
rect 22728 36820 22776 36876
rect 22832 36820 22880 36876
rect 22672 36810 22936 36820
rect 21532 36542 21534 36594
rect 21586 36542 21588 36594
rect 21532 36530 21588 36542
rect 23100 36596 23156 39200
rect 23212 36596 23268 36606
rect 23100 36594 23268 36596
rect 23100 36542 23214 36594
rect 23266 36542 23268 36594
rect 23100 36540 23268 36542
rect 25340 36596 25396 39200
rect 25676 36596 25732 36606
rect 25340 36594 25732 36596
rect 25340 36542 25678 36594
rect 25730 36542 25732 36594
rect 25340 36540 25732 36542
rect 23212 36530 23268 36540
rect 25676 36530 25732 36540
rect 27356 36596 27412 36606
rect 27580 36596 27636 39200
rect 27356 36594 27636 36596
rect 27356 36542 27358 36594
rect 27410 36542 27636 36594
rect 27356 36540 27636 36542
rect 27692 37268 27748 37278
rect 27356 36530 27412 36540
rect 21196 36484 21252 36494
rect 18508 36260 18564 36270
rect 18284 36204 18508 36260
rect 18284 35698 18340 36204
rect 18508 36166 18564 36204
rect 18844 36258 18900 36270
rect 18844 36206 18846 36258
rect 18898 36206 18900 36258
rect 18284 35646 18286 35698
rect 18338 35646 18340 35698
rect 18284 35634 18340 35646
rect 18172 35588 18228 35598
rect 18172 35026 18228 35532
rect 18844 35588 18900 36206
rect 20300 36258 20356 36270
rect 21084 36260 21140 36270
rect 20300 36206 20302 36258
rect 20354 36206 20356 36258
rect 20300 36036 20356 36206
rect 20300 35970 20356 35980
rect 20972 36258 21140 36260
rect 20972 36206 21086 36258
rect 21138 36206 21140 36258
rect 20972 36204 21140 36206
rect 18844 35522 18900 35532
rect 18956 35588 19012 35598
rect 18956 35586 19124 35588
rect 18956 35534 18958 35586
rect 19010 35534 19124 35586
rect 18956 35532 19124 35534
rect 18956 35522 19012 35532
rect 18172 34974 18174 35026
rect 18226 34974 18228 35026
rect 18172 34962 18228 34974
rect 18732 34804 18788 34814
rect 18732 34710 18788 34748
rect 19068 34802 19124 35532
rect 20300 34914 20356 34926
rect 20300 34862 20302 34914
rect 20354 34862 20356 34914
rect 19068 34750 19070 34802
rect 19122 34750 19124 34802
rect 19068 34738 19124 34750
rect 19628 34802 19684 34814
rect 19628 34750 19630 34802
rect 19682 34750 19684 34802
rect 18060 32722 18116 32732
rect 18172 34580 18228 34590
rect 18060 32562 18116 32574
rect 18060 32510 18062 32562
rect 18114 32510 18116 32562
rect 16828 32450 16996 32452
rect 16828 32398 16830 32450
rect 16882 32398 16996 32450
rect 16828 32396 16996 32398
rect 16828 32386 16884 32396
rect 16380 32340 16436 32350
rect 16380 32338 16548 32340
rect 16380 32286 16382 32338
rect 16434 32286 16548 32338
rect 16380 32284 16548 32286
rect 16380 32274 16436 32284
rect 15932 31836 16212 31892
rect 15820 31778 16100 31780
rect 15820 31726 15822 31778
rect 15874 31726 16100 31778
rect 15820 31724 16100 31726
rect 15820 31714 15876 31724
rect 15596 31614 15598 31666
rect 15650 31614 15652 31666
rect 15596 31602 15652 31614
rect 15518 31388 15782 31398
rect 15574 31332 15622 31388
rect 15678 31332 15726 31388
rect 15518 31322 15782 31332
rect 16044 31332 16100 31724
rect 16156 31778 16212 31836
rect 16156 31726 16158 31778
rect 16210 31726 16212 31778
rect 16156 31714 16212 31726
rect 16268 31668 16324 32060
rect 16492 31780 16548 32284
rect 16492 31686 16548 31724
rect 16716 32116 16772 32126
rect 16380 31668 16436 31678
rect 16268 31666 16436 31668
rect 16268 31614 16382 31666
rect 16434 31614 16436 31666
rect 16268 31612 16436 31614
rect 16380 31602 16436 31612
rect 16044 31276 16324 31332
rect 15820 31220 15876 31230
rect 15372 31164 15764 31220
rect 14812 30994 14868 31006
rect 14812 30942 14814 30994
rect 14866 30942 14868 30994
rect 14700 29876 14756 29886
rect 14700 29426 14756 29820
rect 14700 29374 14702 29426
rect 14754 29374 14756 29426
rect 14700 29362 14756 29374
rect 14812 29316 14868 30942
rect 15036 30994 15092 31006
rect 15036 30942 15038 30994
rect 15090 30942 15092 30994
rect 14924 30882 14980 30894
rect 14924 30830 14926 30882
rect 14978 30830 14980 30882
rect 14924 30548 14980 30830
rect 15036 30660 15092 30942
rect 15036 30604 15204 30660
rect 14924 30492 15092 30548
rect 14924 30212 14980 30222
rect 14924 30098 14980 30156
rect 15036 30210 15092 30492
rect 15036 30158 15038 30210
rect 15090 30158 15092 30210
rect 15036 30146 15092 30158
rect 14924 30046 14926 30098
rect 14978 30046 14980 30098
rect 14924 30034 14980 30046
rect 15036 29988 15092 29998
rect 15148 29988 15204 30604
rect 15092 29932 15204 29988
rect 15036 29922 15092 29932
rect 15372 29538 15428 31164
rect 15708 31106 15764 31164
rect 16268 31220 16324 31276
rect 16380 31220 16436 31230
rect 16268 31218 16436 31220
rect 16268 31166 16382 31218
rect 16434 31166 16436 31218
rect 16268 31164 16436 31166
rect 15820 31126 15876 31164
rect 16380 31154 16436 31164
rect 15708 31054 15710 31106
rect 15762 31054 15764 31106
rect 15708 31042 15764 31054
rect 16604 31108 16660 31118
rect 15484 30994 15540 31006
rect 15484 30942 15486 30994
rect 15538 30942 15540 30994
rect 15484 30772 15540 30942
rect 15820 30772 15876 30782
rect 15484 30770 15876 30772
rect 15484 30718 15822 30770
rect 15874 30718 15876 30770
rect 15484 30716 15876 30718
rect 15820 30706 15876 30716
rect 16604 30322 16660 31052
rect 16604 30270 16606 30322
rect 16658 30270 16660 30322
rect 16604 30258 16660 30270
rect 16380 30098 16436 30110
rect 16380 30046 16382 30098
rect 16434 30046 16436 30098
rect 15518 29820 15782 29830
rect 15574 29764 15622 29820
rect 15678 29764 15726 29820
rect 15518 29754 15782 29764
rect 15372 29486 15374 29538
rect 15426 29486 15428 29538
rect 15372 29474 15428 29486
rect 14924 29316 14980 29326
rect 14812 29314 14980 29316
rect 14812 29262 14926 29314
rect 14978 29262 14980 29314
rect 14812 29260 14980 29262
rect 14924 28866 14980 29260
rect 14924 28814 14926 28866
rect 14978 28814 14980 28866
rect 14924 28802 14980 28814
rect 14476 28756 14532 28766
rect 13468 26562 13524 26572
rect 13804 28588 13972 28644
rect 14252 28642 14308 28654
rect 14252 28590 14254 28642
rect 14306 28590 14308 28642
rect 13580 26180 13636 26190
rect 13580 26178 13748 26180
rect 13580 26126 13582 26178
rect 13634 26126 13748 26178
rect 13580 26124 13748 26126
rect 13580 26114 13636 26124
rect 13356 25666 13412 25676
rect 13692 25732 13748 26124
rect 13692 25618 13748 25676
rect 13692 25566 13694 25618
rect 13746 25566 13748 25618
rect 13692 25554 13748 25566
rect 13356 24610 13412 24622
rect 13356 24558 13358 24610
rect 13410 24558 13412 24610
rect 13356 24164 13412 24558
rect 13356 24098 13412 24108
rect 13468 24276 13524 24286
rect 13468 23938 13524 24220
rect 13468 23886 13470 23938
rect 13522 23886 13524 23938
rect 13356 23156 13412 23166
rect 13356 23042 13412 23100
rect 13356 22990 13358 23042
rect 13410 22990 13412 23042
rect 13356 22148 13412 22990
rect 13356 22082 13412 22092
rect 13468 21812 13524 23886
rect 13692 23268 13748 23278
rect 13692 23154 13748 23212
rect 13692 23102 13694 23154
rect 13746 23102 13748 23154
rect 13692 23090 13748 23102
rect 13804 22932 13860 28588
rect 13916 28420 13972 28430
rect 14252 28420 14308 28590
rect 14476 28530 14532 28700
rect 14476 28478 14478 28530
rect 14530 28478 14532 28530
rect 14476 28466 14532 28478
rect 15148 28754 15204 28766
rect 15148 28702 15150 28754
rect 15202 28702 15204 28754
rect 13916 28418 14308 28420
rect 13916 28366 13918 28418
rect 13970 28366 14308 28418
rect 13916 28364 14308 28366
rect 13916 28354 13972 28364
rect 13916 27860 13972 27870
rect 13916 23268 13972 27804
rect 14252 27746 14308 28364
rect 14252 27694 14254 27746
rect 14306 27694 14308 27746
rect 14252 27636 14308 27694
rect 14812 27748 14868 27758
rect 14812 27654 14868 27692
rect 14252 27570 14308 27580
rect 15148 27188 15204 28702
rect 15372 28642 15428 28654
rect 15372 28590 15374 28642
rect 15426 28590 15428 28642
rect 15372 28084 15428 28590
rect 15518 28252 15782 28262
rect 15574 28196 15622 28252
rect 15678 28196 15726 28252
rect 15518 28186 15782 28196
rect 16380 28084 16436 30046
rect 16492 28084 16548 28094
rect 15372 28028 15764 28084
rect 16380 28082 16548 28084
rect 16380 28030 16494 28082
rect 16546 28030 16548 28082
rect 16380 28028 16548 28030
rect 15260 27972 15316 27982
rect 15260 27970 15652 27972
rect 15260 27918 15262 27970
rect 15314 27918 15652 27970
rect 15260 27916 15652 27918
rect 15260 27906 15316 27916
rect 14812 27132 15540 27188
rect 14028 26964 14084 26974
rect 14028 25284 14084 26908
rect 14812 26066 14868 27132
rect 15484 27074 15540 27132
rect 15596 27186 15652 27916
rect 15596 27134 15598 27186
rect 15650 27134 15652 27186
rect 15596 27122 15652 27134
rect 15708 27300 15764 28028
rect 16492 28018 16548 28028
rect 16604 27970 16660 27982
rect 16604 27918 16606 27970
rect 16658 27918 16660 27970
rect 16492 27300 16548 27310
rect 15484 27022 15486 27074
rect 15538 27022 15540 27074
rect 15484 27010 15540 27022
rect 15708 27074 15764 27244
rect 16156 27298 16548 27300
rect 16156 27246 16494 27298
rect 16546 27246 16548 27298
rect 16156 27244 16548 27246
rect 15708 27022 15710 27074
rect 15762 27022 15764 27074
rect 15708 27010 15764 27022
rect 15932 27188 15988 27198
rect 15518 26684 15782 26694
rect 15574 26628 15622 26684
rect 15678 26628 15726 26684
rect 15518 26618 15782 26628
rect 15932 26404 15988 27132
rect 16156 27074 16212 27244
rect 16492 27234 16548 27244
rect 16156 27022 16158 27074
rect 16210 27022 16212 27074
rect 16156 27010 16212 27022
rect 16380 26962 16436 26974
rect 16380 26910 16382 26962
rect 16434 26910 16436 26962
rect 16380 26908 16436 26910
rect 15820 26348 15988 26404
rect 16044 26852 16436 26908
rect 14812 26014 14814 26066
rect 14866 26014 14868 26066
rect 14812 26002 14868 26014
rect 15036 26290 15092 26302
rect 15036 26238 15038 26290
rect 15090 26238 15092 26290
rect 14364 25732 14420 25742
rect 14364 25506 14420 25676
rect 14364 25454 14366 25506
rect 14418 25454 14420 25506
rect 14364 25442 14420 25454
rect 15036 25508 15092 26238
rect 15036 25442 15092 25452
rect 15596 26180 15652 26190
rect 15596 25506 15652 26124
rect 15820 25732 15876 26348
rect 15820 25676 15988 25732
rect 15596 25454 15598 25506
rect 15650 25454 15652 25506
rect 15596 25442 15652 25454
rect 15820 25508 15876 25518
rect 15820 25414 15876 25452
rect 14028 25190 14084 25228
rect 15518 25116 15782 25126
rect 15574 25060 15622 25116
rect 15678 25060 15726 25116
rect 15518 25050 15782 25060
rect 15484 24948 15540 24958
rect 15484 24724 15540 24892
rect 15484 24630 15540 24668
rect 15932 24724 15988 25676
rect 16044 25618 16100 26852
rect 16492 26850 16548 26862
rect 16492 26798 16494 26850
rect 16546 26798 16548 26850
rect 16380 26516 16436 26526
rect 16492 26516 16548 26798
rect 16436 26460 16548 26516
rect 16380 26290 16436 26460
rect 16380 26238 16382 26290
rect 16434 26238 16436 26290
rect 16380 26226 16436 26238
rect 16492 26180 16548 26190
rect 16492 26086 16548 26124
rect 16604 25844 16660 27918
rect 16044 25566 16046 25618
rect 16098 25566 16100 25618
rect 16044 25554 16100 25566
rect 16268 25788 16660 25844
rect 16268 25172 16324 25788
rect 16716 25732 16772 32060
rect 16492 25676 16772 25732
rect 16268 25106 16324 25116
rect 16380 25620 16436 25630
rect 16380 25506 16436 25564
rect 16380 25454 16382 25506
rect 16434 25454 16436 25506
rect 15932 24722 16324 24724
rect 15932 24670 15934 24722
rect 15986 24670 16324 24722
rect 15932 24668 16324 24670
rect 15932 24658 15988 24668
rect 15036 24612 15092 24622
rect 14252 23828 14308 23838
rect 14028 23826 14308 23828
rect 14028 23774 14254 23826
rect 14306 23774 14308 23826
rect 14028 23772 14308 23774
rect 14028 23378 14084 23772
rect 14252 23762 14308 23772
rect 14028 23326 14030 23378
rect 14082 23326 14084 23378
rect 14028 23314 14084 23326
rect 13916 23202 13972 23212
rect 14140 23156 14196 23166
rect 14140 23062 14196 23100
rect 14252 23154 14308 23166
rect 14252 23102 14254 23154
rect 14306 23102 14308 23154
rect 13804 22866 13860 22876
rect 14252 22820 14308 23102
rect 14924 23154 14980 23166
rect 14924 23102 14926 23154
rect 14978 23102 14980 23154
rect 14252 22754 14308 22764
rect 14700 22820 14756 22830
rect 14756 22764 14868 22820
rect 14700 22754 14756 22764
rect 13916 22596 13972 22606
rect 13916 22372 13972 22540
rect 14476 22428 14756 22484
rect 13692 22316 13972 22372
rect 14028 22372 14084 22382
rect 14476 22372 14532 22428
rect 14028 22370 14532 22372
rect 14028 22318 14030 22370
rect 14082 22318 14532 22370
rect 14028 22316 14532 22318
rect 14700 22370 14756 22428
rect 14700 22318 14702 22370
rect 14754 22318 14756 22370
rect 13692 22260 13748 22316
rect 14028 22306 14084 22316
rect 14700 22306 14756 22318
rect 14588 22260 14644 22270
rect 13692 22166 13748 22204
rect 14252 22202 14308 22214
rect 13804 22148 13860 22158
rect 13804 22054 13860 22092
rect 14252 22150 14254 22202
rect 14306 22150 14308 22202
rect 14588 22166 14644 22204
rect 14028 22036 14084 22046
rect 13468 21746 13524 21756
rect 13916 21812 13972 21822
rect 13356 21476 13412 21486
rect 13356 21382 13412 21420
rect 13692 20580 13748 20590
rect 13692 20486 13748 20524
rect 13916 20580 13972 21756
rect 14028 21698 14084 21980
rect 14252 21924 14308 22150
rect 14364 22148 14420 22158
rect 14364 22054 14420 22092
rect 14252 21868 14756 21924
rect 14700 21812 14756 21868
rect 14700 21718 14756 21756
rect 14028 21646 14030 21698
rect 14082 21646 14084 21698
rect 14028 20580 14084 21646
rect 14140 21700 14196 21710
rect 14140 20802 14196 21644
rect 14364 21700 14420 21710
rect 14364 21606 14420 21644
rect 14140 20750 14142 20802
rect 14194 20750 14196 20802
rect 14140 20738 14196 20750
rect 14812 20802 14868 22764
rect 14924 22708 14980 23102
rect 15036 23044 15092 24556
rect 16268 23716 16324 24668
rect 16380 24050 16436 25454
rect 16380 23998 16382 24050
rect 16434 23998 16436 24050
rect 16380 23986 16436 23998
rect 15148 23660 16324 23716
rect 15148 23378 15204 23660
rect 15518 23548 15782 23558
rect 15574 23492 15622 23548
rect 15678 23492 15726 23548
rect 15518 23482 15782 23492
rect 15148 23326 15150 23378
rect 15202 23326 15204 23378
rect 15148 23314 15204 23326
rect 15708 23380 15764 23390
rect 16268 23380 16324 23660
rect 16380 23380 16436 23390
rect 16268 23378 16436 23380
rect 16268 23326 16382 23378
rect 16434 23326 16436 23378
rect 16268 23324 16436 23326
rect 15708 23286 15764 23324
rect 16380 23314 16436 23324
rect 15036 22978 15092 22988
rect 15260 23156 15316 23166
rect 15596 23156 15652 23166
rect 15260 23154 15652 23156
rect 15260 23102 15262 23154
rect 15314 23102 15598 23154
rect 15650 23102 15652 23154
rect 15260 23100 15652 23102
rect 15260 22932 15316 23100
rect 15596 23090 15652 23100
rect 15932 23156 15988 23166
rect 15932 23062 15988 23100
rect 14924 22642 14980 22652
rect 15148 22876 15316 22932
rect 15036 22372 15092 22382
rect 14924 22370 15092 22372
rect 14924 22318 15038 22370
rect 15090 22318 15092 22370
rect 14924 22316 15092 22318
rect 14924 21812 14980 22316
rect 15036 22306 15092 22316
rect 15036 22148 15092 22158
rect 15148 22148 15204 22876
rect 15260 22708 15316 22718
rect 15260 22372 15316 22652
rect 15932 22596 15988 22606
rect 15988 22540 16100 22596
rect 15932 22530 15988 22540
rect 15708 22372 15764 22382
rect 15260 22370 15764 22372
rect 15260 22318 15262 22370
rect 15314 22318 15710 22370
rect 15762 22318 15764 22370
rect 15260 22316 15764 22318
rect 15260 22306 15316 22316
rect 15708 22306 15764 22316
rect 15932 22260 15988 22270
rect 15932 22166 15988 22204
rect 15148 22092 15428 22148
rect 15036 22054 15092 22092
rect 15260 21812 15316 21822
rect 14924 21810 15316 21812
rect 14924 21758 15262 21810
rect 15314 21758 15316 21810
rect 14924 21756 15316 21758
rect 15260 21746 15316 21756
rect 15372 21700 15428 22092
rect 16044 22036 16100 22540
rect 16268 22484 16324 22494
rect 16268 22370 16324 22428
rect 16268 22318 16270 22370
rect 16322 22318 16324 22370
rect 16268 22306 16324 22318
rect 15518 21980 15782 21990
rect 15574 21924 15622 21980
rect 15678 21924 15726 21980
rect 15518 21914 15782 21924
rect 15932 21980 16100 22036
rect 16156 22146 16212 22158
rect 16156 22094 16158 22146
rect 16210 22094 16212 22146
rect 15372 21634 15428 21644
rect 15484 21698 15540 21710
rect 15484 21646 15486 21698
rect 15538 21646 15540 21698
rect 14812 20750 14814 20802
rect 14866 20750 14868 20802
rect 14812 20738 14868 20750
rect 14924 21586 14980 21598
rect 14924 21534 14926 21586
rect 14978 21534 14980 21586
rect 14924 20692 14980 21534
rect 15484 21588 15540 21646
rect 15596 21700 15652 21710
rect 15596 21606 15652 21644
rect 15932 21698 15988 21980
rect 15932 21646 15934 21698
rect 15986 21646 15988 21698
rect 15932 21634 15988 21646
rect 16044 21700 16100 21710
rect 16044 21606 16100 21644
rect 15484 21522 15540 21532
rect 15036 21364 15092 21374
rect 16044 21364 16100 21374
rect 15036 20802 15092 21308
rect 15596 21362 16100 21364
rect 15596 21310 16046 21362
rect 16098 21310 16100 21362
rect 15596 21308 16100 21310
rect 15484 21252 15540 21262
rect 15036 20750 15038 20802
rect 15090 20750 15092 20802
rect 15036 20738 15092 20750
rect 15148 21196 15484 21252
rect 14364 20580 14420 20590
rect 14028 20578 14420 20580
rect 14028 20526 14366 20578
rect 14418 20526 14420 20578
rect 14028 20524 14420 20526
rect 13916 20018 13972 20524
rect 14364 20514 14420 20524
rect 14924 20356 14980 20636
rect 14924 20290 14980 20300
rect 15036 20578 15092 20590
rect 15036 20526 15038 20578
rect 15090 20526 15092 20578
rect 14700 20132 14756 20142
rect 15036 20132 15092 20526
rect 14700 20130 15092 20132
rect 14700 20078 14702 20130
rect 14754 20078 15092 20130
rect 14700 20076 15092 20078
rect 14700 20066 14756 20076
rect 13916 19966 13918 20018
rect 13970 19966 13972 20018
rect 13916 19954 13972 19966
rect 13692 19908 13748 19918
rect 13692 19814 13748 19852
rect 14588 19908 14644 19918
rect 13468 19796 13524 19806
rect 13468 19234 13524 19740
rect 13468 19182 13470 19234
rect 13522 19182 13524 19234
rect 13468 19170 13524 19182
rect 13692 19404 13972 19460
rect 13692 18674 13748 19404
rect 13804 19234 13860 19246
rect 13804 19182 13806 19234
rect 13858 19182 13860 19234
rect 13804 19012 13860 19182
rect 13916 19236 13972 19404
rect 14028 19236 14084 19246
rect 13916 19234 14084 19236
rect 13916 19182 14030 19234
rect 14082 19182 14084 19234
rect 13916 19180 14084 19182
rect 14028 19170 14084 19180
rect 14588 19122 14644 19852
rect 14588 19070 14590 19122
rect 14642 19070 14644 19122
rect 14588 19058 14644 19070
rect 14700 19124 14756 19134
rect 14700 19122 14868 19124
rect 14700 19070 14702 19122
rect 14754 19070 14868 19122
rect 14700 19068 14868 19070
rect 14700 19058 14756 19068
rect 13804 18946 13860 18956
rect 13916 19012 13972 19022
rect 14364 19012 14420 19022
rect 13916 19010 14308 19012
rect 13916 18958 13918 19010
rect 13970 18958 14308 19010
rect 13916 18956 14308 18958
rect 13916 18946 13972 18956
rect 13692 18622 13694 18674
rect 13746 18622 13748 18674
rect 13692 18610 13748 18622
rect 14252 18676 14308 18956
rect 14364 18918 14420 18956
rect 14252 18620 14756 18676
rect 13468 18562 13524 18574
rect 13468 18510 13470 18562
rect 13522 18510 13524 18562
rect 13244 18386 13300 18396
rect 13356 18450 13412 18462
rect 13356 18398 13358 18450
rect 13410 18398 13412 18450
rect 13020 17836 13188 17892
rect 12908 17726 12910 17778
rect 12962 17726 12964 17778
rect 12908 17714 12964 17726
rect 12796 17054 12798 17106
rect 12850 17054 12852 17106
rect 12684 16996 12740 17006
rect 12572 16994 12740 16996
rect 12572 16942 12686 16994
rect 12738 16942 12740 16994
rect 12572 16940 12740 16942
rect 12684 16930 12740 16940
rect 12684 16324 12740 16334
rect 12460 16322 12740 16324
rect 12460 16270 12686 16322
rect 12738 16270 12740 16322
rect 12460 16268 12740 16270
rect 12236 15988 12292 15998
rect 12236 15894 12292 15932
rect 12124 15596 12292 15652
rect 12124 15148 12180 15158
rect 12012 15092 12124 15148
rect 12124 15082 12180 15092
rect 12124 14532 12180 14542
rect 12124 14438 12180 14476
rect 12124 13746 12180 13758
rect 12124 13694 12126 13746
rect 12178 13694 12180 13746
rect 12124 13300 12180 13694
rect 12124 13234 12180 13244
rect 11900 12338 11956 12348
rect 12236 12180 12292 15596
rect 12348 15204 12404 15214
rect 12348 14642 12404 15148
rect 12348 14590 12350 14642
rect 12402 14590 12404 14642
rect 12348 14578 12404 14590
rect 12460 13858 12516 16268
rect 12684 16258 12740 16268
rect 12572 16100 12628 16110
rect 12572 16006 12628 16044
rect 12684 15988 12740 15998
rect 12796 15988 12852 17054
rect 13020 17668 13076 17678
rect 13020 17106 13076 17612
rect 13020 17054 13022 17106
rect 13074 17054 13076 17106
rect 13020 17042 13076 17054
rect 12684 15986 12852 15988
rect 12684 15934 12686 15986
rect 12738 15934 12852 15986
rect 12684 15932 12852 15934
rect 13132 16884 13188 17836
rect 13356 17780 13412 18398
rect 13468 18116 13524 18510
rect 14700 18562 14756 18620
rect 14700 18510 14702 18562
rect 14754 18510 14756 18562
rect 14700 18498 14756 18510
rect 13468 18050 13524 18060
rect 13916 18450 13972 18462
rect 13916 18398 13918 18450
rect 13970 18398 13972 18450
rect 13356 17668 13412 17724
rect 13468 17668 13524 17678
rect 13356 17666 13524 17668
rect 13356 17614 13470 17666
rect 13522 17614 13524 17666
rect 13356 17612 13524 17614
rect 13468 17602 13524 17612
rect 13580 17556 13636 17566
rect 13580 17462 13636 17500
rect 13804 17442 13860 17454
rect 13804 17390 13806 17442
rect 13858 17390 13860 17442
rect 13356 17108 13412 17118
rect 13412 17052 13636 17108
rect 13356 17014 13412 17052
rect 12684 15540 12740 15932
rect 12684 15474 12740 15484
rect 13132 15148 13188 16828
rect 13244 16996 13300 17006
rect 13244 16660 13300 16940
rect 13468 16882 13524 16894
rect 13468 16830 13470 16882
rect 13522 16830 13524 16882
rect 13356 16660 13412 16670
rect 13244 16658 13412 16660
rect 13244 16606 13358 16658
rect 13410 16606 13412 16658
rect 13244 16604 13412 16606
rect 13356 16594 13412 16604
rect 12684 15092 12740 15102
rect 12572 14420 12628 14430
rect 12572 14326 12628 14364
rect 12460 13806 12462 13858
rect 12514 13806 12516 13858
rect 12460 13794 12516 13806
rect 12572 13636 12628 13646
rect 12348 13634 12628 13636
rect 12348 13582 12574 13634
rect 12626 13582 12628 13634
rect 12348 13580 12628 13582
rect 12348 12290 12404 13580
rect 12572 13570 12628 13580
rect 12460 13412 12516 13422
rect 12460 12964 12516 13356
rect 12572 13300 12628 13310
rect 12684 13300 12740 15036
rect 12796 15092 13188 15148
rect 12796 14532 12852 15092
rect 12796 14530 12964 14532
rect 12796 14478 12798 14530
rect 12850 14478 12964 14530
rect 12796 14476 12964 14478
rect 12796 14466 12852 14476
rect 12796 13748 12852 13758
rect 12796 13654 12852 13692
rect 12908 13746 12964 14476
rect 13468 14308 13524 16830
rect 13580 16100 13636 17052
rect 13804 16996 13860 17390
rect 13804 16930 13860 16940
rect 13916 16212 13972 18398
rect 14812 18004 14868 19068
rect 14812 17938 14868 17948
rect 15036 17892 15092 17902
rect 14588 17724 14980 17780
rect 14028 17668 14084 17678
rect 14028 17574 14084 17612
rect 14476 17668 14532 17678
rect 14588 17668 14644 17724
rect 14476 17666 14644 17668
rect 14476 17614 14478 17666
rect 14530 17614 14644 17666
rect 14476 17612 14644 17614
rect 14924 17666 14980 17724
rect 14924 17614 14926 17666
rect 14978 17614 14980 17666
rect 14476 17602 14532 17612
rect 14924 17602 14980 17614
rect 14252 17556 14308 17566
rect 14028 17444 14084 17454
rect 14028 17106 14084 17388
rect 14028 17054 14030 17106
rect 14082 17054 14084 17106
rect 14028 16772 14084 17054
rect 14252 17108 14308 17500
rect 14700 17554 14756 17566
rect 14700 17502 14702 17554
rect 14754 17502 14756 17554
rect 14364 17444 14420 17454
rect 14364 17442 14532 17444
rect 14364 17390 14366 17442
rect 14418 17390 14532 17442
rect 14364 17388 14532 17390
rect 14364 17378 14420 17388
rect 14364 17108 14420 17118
rect 14252 17106 14420 17108
rect 14252 17054 14366 17106
rect 14418 17054 14420 17106
rect 14252 17052 14420 17054
rect 14364 17042 14420 17052
rect 14476 17108 14532 17388
rect 14476 17042 14532 17052
rect 14700 16884 14756 17502
rect 14700 16790 14756 16828
rect 15036 16882 15092 17836
rect 15148 17554 15204 21196
rect 15484 21186 15540 21196
rect 15372 20804 15428 20814
rect 15596 20804 15652 21308
rect 16044 21298 16100 21308
rect 16156 20916 16212 22094
rect 16492 22036 16548 25676
rect 16716 25396 16772 25406
rect 16716 25282 16772 25340
rect 16716 25230 16718 25282
rect 16770 25230 16772 25282
rect 16604 23380 16660 23390
rect 16716 23380 16772 25230
rect 16660 23324 16772 23380
rect 16604 23314 16660 23324
rect 16380 21980 16548 22036
rect 16716 22146 16772 22158
rect 16716 22094 16718 22146
rect 16770 22094 16772 22146
rect 16716 22036 16772 22094
rect 16380 21252 16436 21980
rect 16380 21186 16436 21196
rect 16492 21700 16548 21710
rect 16268 21140 16324 21150
rect 16268 21026 16324 21084
rect 16268 20974 16270 21026
rect 16322 20974 16324 21026
rect 16268 20962 16324 20974
rect 16156 20850 16212 20860
rect 15372 20802 15652 20804
rect 15372 20750 15374 20802
rect 15426 20750 15652 20802
rect 15372 20748 15652 20750
rect 16268 20804 16324 20814
rect 15372 20738 15428 20748
rect 15932 20692 15988 20702
rect 15518 20412 15782 20422
rect 15574 20356 15622 20412
rect 15678 20356 15726 20412
rect 15518 20346 15782 20356
rect 15932 20244 15988 20636
rect 15932 20178 15988 20188
rect 16268 19236 16324 20748
rect 16044 19180 16324 19236
rect 15820 19124 15876 19134
rect 15484 19012 15540 19050
rect 15820 19030 15876 19068
rect 15484 18946 15540 18956
rect 15932 19012 15988 19022
rect 15932 18918 15988 18956
rect 15518 18844 15782 18854
rect 15574 18788 15622 18844
rect 15678 18788 15726 18844
rect 15518 18778 15782 18788
rect 15148 17502 15150 17554
rect 15202 17502 15204 17554
rect 15148 17490 15204 17502
rect 15260 18004 15316 18014
rect 15260 17556 15316 17948
rect 15820 17556 15876 17566
rect 15260 17462 15316 17500
rect 15372 17554 15876 17556
rect 15372 17502 15822 17554
rect 15874 17502 15876 17554
rect 15372 17500 15876 17502
rect 15260 16996 15316 17006
rect 15260 16902 15316 16940
rect 15036 16830 15038 16882
rect 15090 16830 15092 16882
rect 15036 16818 15092 16830
rect 15372 16884 15428 17500
rect 15820 17490 15876 17500
rect 16044 17554 16100 19180
rect 16156 19012 16212 19022
rect 16492 19012 16548 21644
rect 16604 21588 16660 21598
rect 16604 21494 16660 21532
rect 16604 20804 16660 20814
rect 16604 20710 16660 20748
rect 16716 20020 16772 21980
rect 16716 19954 16772 19964
rect 16828 19906 16884 19918
rect 16828 19854 16830 19906
rect 16882 19854 16884 19906
rect 16828 19684 16884 19854
rect 16716 19628 16884 19684
rect 16716 19124 16772 19628
rect 16828 19458 16884 19470
rect 16828 19406 16830 19458
rect 16882 19406 16884 19458
rect 16828 19346 16884 19406
rect 16828 19294 16830 19346
rect 16882 19294 16884 19346
rect 16828 19282 16884 19294
rect 16716 19068 16884 19124
rect 16156 19010 16436 19012
rect 16156 18958 16158 19010
rect 16210 18958 16436 19010
rect 16156 18956 16436 18958
rect 16156 18946 16212 18956
rect 16044 17502 16046 17554
rect 16098 17502 16100 17554
rect 16044 17332 16100 17502
rect 15518 17276 15782 17286
rect 15574 17220 15622 17276
rect 15678 17220 15726 17276
rect 16044 17266 16100 17276
rect 16156 17778 16212 17790
rect 16156 17726 16158 17778
rect 16210 17726 16212 17778
rect 15518 17210 15782 17220
rect 15372 16818 15428 16828
rect 15708 16996 15764 17006
rect 16156 16996 16212 17726
rect 14028 16706 14084 16716
rect 14812 16772 14868 16782
rect 14364 16212 14420 16222
rect 13916 16156 14084 16212
rect 13580 16044 13972 16100
rect 13916 15874 13972 16044
rect 14028 15988 14084 16156
rect 14364 16118 14420 16156
rect 14028 15922 14084 15932
rect 13916 15822 13918 15874
rect 13970 15822 13972 15874
rect 13804 15204 13860 15242
rect 13804 15138 13860 15148
rect 13692 14308 13748 14318
rect 13468 14252 13692 14308
rect 13692 14214 13748 14252
rect 13356 13860 13412 13870
rect 13356 13766 13412 13804
rect 13468 13860 13524 13870
rect 13468 13858 13636 13860
rect 13468 13806 13470 13858
rect 13522 13806 13636 13858
rect 13468 13804 13636 13806
rect 13468 13794 13524 13804
rect 12908 13694 12910 13746
rect 12962 13694 12964 13746
rect 12908 13682 12964 13694
rect 12628 13244 12740 13300
rect 12572 13234 12628 13244
rect 12460 12962 12852 12964
rect 12460 12910 12462 12962
rect 12514 12910 12852 12962
rect 12460 12908 12852 12910
rect 12460 12898 12516 12908
rect 12572 12404 12628 12414
rect 12628 12348 12740 12404
rect 12572 12338 12628 12348
rect 12348 12238 12350 12290
rect 12402 12238 12404 12290
rect 12348 12226 12404 12238
rect 11564 12178 11844 12180
rect 11564 12126 11566 12178
rect 11618 12126 11844 12178
rect 11564 12124 11844 12126
rect 11900 12124 12292 12180
rect 11564 11844 11620 12124
rect 11564 11778 11620 11788
rect 11900 11506 11956 12124
rect 12236 12068 12292 12124
rect 12236 12012 12628 12068
rect 11900 11454 11902 11506
rect 11954 11454 11956 11506
rect 11900 11442 11956 11454
rect 12348 11844 12404 11854
rect 11452 11396 11508 11406
rect 11340 11394 11508 11396
rect 11340 11342 11454 11394
rect 11506 11342 11508 11394
rect 11340 11340 11508 11342
rect 10892 10668 11060 10724
rect 10892 9828 10948 10668
rect 11004 10500 11060 10510
rect 11452 10500 11508 11340
rect 12348 11396 12404 11788
rect 12348 11302 12404 11340
rect 12572 10610 12628 12012
rect 12684 11506 12740 12348
rect 12684 11454 12686 11506
rect 12738 11454 12740 11506
rect 12684 10722 12740 11454
rect 12684 10670 12686 10722
rect 12738 10670 12740 10722
rect 12684 10658 12740 10670
rect 12572 10558 12574 10610
rect 12626 10558 12628 10610
rect 12572 10546 12628 10558
rect 12796 10500 12852 12908
rect 13468 12850 13524 12862
rect 13468 12798 13470 12850
rect 13522 12798 13524 12850
rect 13020 12740 13076 12750
rect 13020 12646 13076 12684
rect 13468 12628 13524 12798
rect 13468 12562 13524 12572
rect 11452 10444 11620 10500
rect 11004 10276 11060 10444
rect 11004 10220 11508 10276
rect 11004 10052 11060 10062
rect 11004 9958 11060 9996
rect 10892 9772 11172 9828
rect 11004 9604 11060 9614
rect 11004 9154 11060 9548
rect 11004 9102 11006 9154
rect 11058 9102 11060 9154
rect 11004 9090 11060 9102
rect 11116 8932 11172 9772
rect 11452 9826 11508 10220
rect 11452 9774 11454 9826
rect 11506 9774 11508 9826
rect 11452 9762 11508 9774
rect 10780 6692 10836 7980
rect 10780 6626 10836 6636
rect 11004 8876 11172 8932
rect 11228 9714 11284 9726
rect 11228 9662 11230 9714
rect 11282 9662 11284 9714
rect 11228 8932 11284 9662
rect 9772 6130 10276 6132
rect 9772 6078 9774 6130
rect 9826 6078 10222 6130
rect 10274 6078 10276 6130
rect 9772 6076 10276 6078
rect 9772 6066 9828 6076
rect 10220 6066 10276 6076
rect 10780 6466 10836 6478
rect 10780 6414 10782 6466
rect 10834 6414 10836 6466
rect 10780 6356 10836 6414
rect 10444 6020 10500 6030
rect 8876 5182 8878 5234
rect 8930 5182 8932 5234
rect 8876 5170 8932 5182
rect 8988 5346 9156 5348
rect 8988 5294 9102 5346
rect 9154 5294 9156 5346
rect 8988 5292 9156 5294
rect 8988 5236 9044 5292
rect 9100 5282 9156 5292
rect 10108 5348 10164 5358
rect 8988 5170 9044 5180
rect 9212 5236 9268 5246
rect 9212 5142 9268 5180
rect 9772 5236 9828 5246
rect 8204 5058 8260 5068
rect 9548 5124 9604 5134
rect 9548 5030 9604 5068
rect 9772 5010 9828 5180
rect 9772 4958 9774 5010
rect 9826 4958 9828 5010
rect 9772 4946 9828 4958
rect 9884 5234 9940 5246
rect 9884 5182 9886 5234
rect 9938 5182 9940 5234
rect 8092 4900 8148 4910
rect 8092 4450 8148 4844
rect 8988 4564 9044 4574
rect 8988 4470 9044 4508
rect 8092 4398 8094 4450
rect 8146 4398 8148 4450
rect 8092 4386 8148 4398
rect 8428 4450 8484 4462
rect 8428 4398 8430 4450
rect 8482 4398 8484 4450
rect 8428 4116 8484 4398
rect 9884 4450 9940 5182
rect 10108 4562 10164 5292
rect 10444 5236 10500 5964
rect 10780 6018 10836 6300
rect 10780 5966 10782 6018
rect 10834 5966 10836 6018
rect 10780 5954 10836 5966
rect 10444 5122 10500 5180
rect 10444 5070 10446 5122
rect 10498 5070 10500 5122
rect 10444 5058 10500 5070
rect 10668 5122 10724 5134
rect 10668 5070 10670 5122
rect 10722 5070 10724 5122
rect 10108 4510 10110 4562
rect 10162 4510 10164 4562
rect 10108 4498 10164 4510
rect 10220 5010 10276 5022
rect 10220 4958 10222 5010
rect 10274 4958 10276 5010
rect 9884 4398 9886 4450
rect 9938 4398 9940 4450
rect 9884 4386 9940 4398
rect 8428 4050 8484 4060
rect 8876 4226 8932 4238
rect 8876 4174 8878 4226
rect 8930 4174 8932 4226
rect 8365 3948 8629 3958
rect 8421 3892 8469 3948
rect 8525 3892 8573 3948
rect 8365 3882 8629 3892
rect 8876 3892 8932 4174
rect 10220 4226 10276 4958
rect 10668 4452 10724 5070
rect 10780 5124 10836 5134
rect 10780 5030 10836 5068
rect 11004 5122 11060 8876
rect 11228 8866 11284 8876
rect 11228 6580 11284 6590
rect 11228 6244 11284 6524
rect 11340 6466 11396 6478
rect 11340 6414 11342 6466
rect 11394 6414 11396 6466
rect 11340 6356 11396 6414
rect 11564 6356 11620 10444
rect 12684 10444 12852 10500
rect 13468 11284 13524 11294
rect 13580 11284 13636 13804
rect 13692 13748 13748 13758
rect 13692 13654 13748 13692
rect 13804 13300 13860 13310
rect 13804 12850 13860 13244
rect 13804 12798 13806 12850
rect 13858 12798 13860 12850
rect 13804 12786 13860 12798
rect 13916 11788 13972 15822
rect 14588 15314 14644 15326
rect 14588 15262 14590 15314
rect 14642 15262 14644 15314
rect 14588 15204 14644 15262
rect 14812 15148 14868 16716
rect 15148 16770 15204 16782
rect 15148 16718 15150 16770
rect 15202 16718 15204 16770
rect 15148 16436 15204 16718
rect 15148 16380 15652 16436
rect 15596 16210 15652 16380
rect 15596 16158 15598 16210
rect 15650 16158 15652 16210
rect 15596 16146 15652 16158
rect 14588 15138 14644 15148
rect 14028 15092 14084 15102
rect 14028 13970 14084 15036
rect 14700 15092 14868 15148
rect 14924 16098 14980 16110
rect 14924 16046 14926 16098
rect 14978 16046 14980 16098
rect 14924 15988 14980 16046
rect 15708 15988 15764 16940
rect 16044 16940 16212 16996
rect 16268 17444 16324 17454
rect 14924 15204 14980 15932
rect 15372 15932 15764 15988
rect 15932 16884 15988 16894
rect 15036 15316 15092 15326
rect 15372 15316 15428 15932
rect 15518 15708 15782 15718
rect 15574 15652 15622 15708
rect 15678 15652 15726 15708
rect 15518 15642 15782 15652
rect 15484 15540 15540 15550
rect 15484 15446 15540 15484
rect 15932 15538 15988 16828
rect 16044 16660 16100 16940
rect 16268 16884 16324 17388
rect 16268 16818 16324 16828
rect 16268 16660 16324 16670
rect 16044 16658 16324 16660
rect 16044 16606 16270 16658
rect 16322 16606 16324 16658
rect 16044 16604 16324 16606
rect 16380 16660 16436 18956
rect 16492 18946 16548 18956
rect 16828 18788 16884 19068
rect 16828 18722 16884 18732
rect 16828 18338 16884 18350
rect 16828 18286 16830 18338
rect 16882 18286 16884 18338
rect 16604 17892 16660 17902
rect 16604 17798 16660 17836
rect 16716 17780 16772 17790
rect 16492 17556 16548 17566
rect 16492 17220 16548 17500
rect 16604 17556 16660 17566
rect 16716 17556 16772 17724
rect 16604 17554 16772 17556
rect 16604 17502 16606 17554
rect 16658 17502 16772 17554
rect 16604 17500 16772 17502
rect 16604 17490 16660 17500
rect 16828 17220 16884 18286
rect 16940 18340 16996 32396
rect 17052 31780 17108 31790
rect 17052 31686 17108 31724
rect 17388 31666 17444 31678
rect 17388 31614 17390 31666
rect 17442 31614 17444 31666
rect 17276 31554 17332 31566
rect 17276 31502 17278 31554
rect 17330 31502 17332 31554
rect 17276 30772 17332 31502
rect 17388 31444 17444 31614
rect 17388 31378 17444 31388
rect 17948 31556 18004 31566
rect 17612 30884 17668 30894
rect 17948 30884 18004 31500
rect 18060 31444 18116 32510
rect 18060 31378 18116 31388
rect 17612 30882 18004 30884
rect 17612 30830 17614 30882
rect 17666 30830 18004 30882
rect 17612 30828 18004 30830
rect 17612 30772 17668 30828
rect 17164 30716 17668 30772
rect 17052 30212 17108 30222
rect 17052 29988 17108 30156
rect 17052 29894 17108 29932
rect 17164 26908 17220 30716
rect 17612 29988 17668 29998
rect 17276 27188 17332 27198
rect 17276 27094 17332 27132
rect 16940 18274 16996 18284
rect 17052 26852 17220 26908
rect 16492 17164 16772 17220
rect 16828 17164 16996 17220
rect 16716 16996 16772 17164
rect 16828 16996 16884 17006
rect 16716 16994 16884 16996
rect 16716 16942 16830 16994
rect 16882 16942 16884 16994
rect 16716 16940 16884 16942
rect 16828 16930 16884 16940
rect 16604 16884 16660 16894
rect 16604 16790 16660 16828
rect 16716 16770 16772 16782
rect 16716 16718 16718 16770
rect 16770 16718 16772 16770
rect 16380 16604 16660 16660
rect 16268 16594 16324 16604
rect 15932 15486 15934 15538
rect 15986 15486 15988 15538
rect 15092 15260 15428 15316
rect 15036 15222 15092 15260
rect 14924 15138 14980 15148
rect 14700 15026 14756 15036
rect 14812 15090 14868 15092
rect 14812 15038 14814 15090
rect 14866 15038 14868 15090
rect 14812 15026 14868 15038
rect 14588 14644 14644 14654
rect 14588 14550 14644 14588
rect 14700 14532 14756 14542
rect 14140 14420 14196 14430
rect 14140 14326 14196 14364
rect 14028 13918 14030 13970
rect 14082 13918 14084 13970
rect 14028 13906 14084 13918
rect 14364 13858 14420 13870
rect 14364 13806 14366 13858
rect 14418 13806 14420 13858
rect 14364 13524 14420 13806
rect 14700 13746 14756 14476
rect 15036 14420 15092 14430
rect 15036 14326 15092 14364
rect 15260 14420 15316 14430
rect 14700 13694 14702 13746
rect 14754 13694 14756 13746
rect 14700 13636 14756 13694
rect 15148 14306 15204 14318
rect 15148 14254 15150 14306
rect 15202 14254 15204 14306
rect 15148 13748 15204 14254
rect 15148 13682 15204 13692
rect 15260 13748 15316 14364
rect 15372 13972 15428 15260
rect 15596 15090 15652 15102
rect 15596 15038 15598 15090
rect 15650 15038 15652 15090
rect 15596 14530 15652 15038
rect 15932 14644 15988 15486
rect 16380 15540 16436 15550
rect 15988 14588 16100 14644
rect 15932 14578 15988 14588
rect 15596 14478 15598 14530
rect 15650 14478 15652 14530
rect 15596 14466 15652 14478
rect 15932 14420 15988 14430
rect 15932 14326 15988 14364
rect 15518 14140 15782 14150
rect 15574 14084 15622 14140
rect 15678 14084 15726 14140
rect 15518 14074 15782 14084
rect 15596 13972 15652 13982
rect 15372 13970 15652 13972
rect 15372 13918 15598 13970
rect 15650 13918 15652 13970
rect 15372 13916 15652 13918
rect 15596 13906 15652 13916
rect 15372 13748 15428 13758
rect 15260 13746 15428 13748
rect 15260 13694 15374 13746
rect 15426 13694 15428 13746
rect 15260 13692 15428 13694
rect 14700 13570 14756 13580
rect 14924 13634 14980 13646
rect 14924 13582 14926 13634
rect 14978 13582 14980 13634
rect 14364 13458 14420 13468
rect 14924 13300 14980 13582
rect 15036 13524 15092 13534
rect 15260 13524 15316 13692
rect 15372 13682 15428 13692
rect 16044 13746 16100 14588
rect 16380 14532 16436 15484
rect 16604 15148 16660 16604
rect 16716 15428 16772 16718
rect 16940 15988 16996 17164
rect 17052 16884 17108 26852
rect 17500 26180 17556 26190
rect 17164 25620 17220 25630
rect 17164 25526 17220 25564
rect 17500 24834 17556 26124
rect 17500 24782 17502 24834
rect 17554 24782 17556 24834
rect 17500 24770 17556 24782
rect 17388 23716 17444 23726
rect 17388 23622 17444 23660
rect 17388 23156 17444 23166
rect 17388 23062 17444 23100
rect 17500 21700 17556 21710
rect 17500 21606 17556 21644
rect 17388 20916 17444 20926
rect 17388 20822 17444 20860
rect 17500 20244 17556 20254
rect 17500 20130 17556 20188
rect 17500 20078 17502 20130
rect 17554 20078 17556 20130
rect 17500 20066 17556 20078
rect 17612 20132 17668 29932
rect 18172 29876 18228 34524
rect 19068 34580 19124 34590
rect 18956 34132 19012 34142
rect 18956 34038 19012 34076
rect 18284 34018 18340 34030
rect 18284 33966 18286 34018
rect 18338 33966 18340 34018
rect 18284 33796 18340 33966
rect 18284 33730 18340 33740
rect 18732 34018 18788 34030
rect 18732 33966 18734 34018
rect 18786 33966 18788 34018
rect 18732 33460 18788 33966
rect 18732 33394 18788 33404
rect 18844 33908 18900 33918
rect 18508 32564 18564 32574
rect 18508 31890 18564 32508
rect 18508 31838 18510 31890
rect 18562 31838 18564 31890
rect 18508 31826 18564 31838
rect 18732 32452 18788 32462
rect 18284 31780 18340 31790
rect 18284 31686 18340 31724
rect 18732 31666 18788 32396
rect 18732 31614 18734 31666
rect 18786 31614 18788 31666
rect 18732 31602 18788 31614
rect 18396 30882 18452 30894
rect 18396 30830 18398 30882
rect 18450 30830 18452 30882
rect 18396 30324 18452 30830
rect 18844 30884 18900 33852
rect 18956 33460 19012 33470
rect 19068 33460 19124 34524
rect 19628 34244 19684 34750
rect 20300 34804 20356 34862
rect 20300 34356 20356 34748
rect 20524 34914 20580 34926
rect 20524 34862 20526 34914
rect 20578 34862 20580 34914
rect 20524 34692 20580 34862
rect 20524 34626 20580 34636
rect 20972 34580 21028 36204
rect 21084 36194 21140 36204
rect 21084 35588 21140 35598
rect 21196 35588 21252 36428
rect 25004 36484 25060 36494
rect 25004 36390 25060 36428
rect 22540 36258 22596 36270
rect 22764 36260 22820 36270
rect 22540 36206 22542 36258
rect 22594 36206 22596 36258
rect 21084 35586 21252 35588
rect 21084 35534 21086 35586
rect 21138 35534 21252 35586
rect 21084 35532 21252 35534
rect 21308 36036 21364 36046
rect 22540 36036 22596 36206
rect 21084 35522 21140 35532
rect 21308 35028 21364 35980
rect 22316 35980 22596 36036
rect 22652 36258 22820 36260
rect 22652 36206 22766 36258
rect 22818 36206 22820 36258
rect 22652 36204 22820 36206
rect 21644 35924 21700 35962
rect 21644 35858 21700 35868
rect 20972 34514 21028 34524
rect 21196 34972 21364 35028
rect 21420 35698 21476 35710
rect 21420 35646 21422 35698
rect 21474 35646 21476 35698
rect 21420 35028 21476 35646
rect 20412 34356 20468 34366
rect 20300 34354 20468 34356
rect 20300 34302 20414 34354
rect 20466 34302 20468 34354
rect 20300 34300 20468 34302
rect 21196 34356 21252 34972
rect 21420 34962 21476 34972
rect 21644 35700 21700 35710
rect 21644 34916 21700 35644
rect 21756 35476 21812 35486
rect 22092 35476 22148 35486
rect 21756 35474 22148 35476
rect 21756 35422 21758 35474
rect 21810 35422 22094 35474
rect 22146 35422 22148 35474
rect 21756 35420 22148 35422
rect 21756 35410 21812 35420
rect 22092 35410 22148 35420
rect 22316 35028 22372 35980
rect 22652 35924 22708 36204
rect 22764 36194 22820 36204
rect 24108 36260 24164 36270
rect 24668 36260 24724 36270
rect 24108 36258 24276 36260
rect 24108 36206 24110 36258
rect 24162 36206 24276 36258
rect 24108 36204 24276 36206
rect 24108 36194 24164 36204
rect 22428 35868 22708 35924
rect 22764 36036 22820 36046
rect 22428 35140 22484 35868
rect 22764 35810 22820 35980
rect 22764 35758 22766 35810
rect 22818 35758 22820 35810
rect 22764 35746 22820 35758
rect 22876 35924 22932 35934
rect 22428 35074 22484 35084
rect 22540 35698 22596 35710
rect 22540 35646 22542 35698
rect 22594 35646 22596 35698
rect 21532 34914 21700 34916
rect 21532 34862 21646 34914
rect 21698 34862 21700 34914
rect 21532 34860 21700 34862
rect 21308 34802 21364 34814
rect 21308 34750 21310 34802
rect 21362 34750 21364 34802
rect 21308 34580 21364 34750
rect 21420 34804 21476 34814
rect 21420 34710 21476 34748
rect 21308 34514 21364 34524
rect 21196 34300 21476 34356
rect 20412 34290 20468 34300
rect 19628 34178 19684 34188
rect 19516 34130 19572 34142
rect 19516 34078 19518 34130
rect 19570 34078 19572 34130
rect 19516 33908 19572 34078
rect 19852 34132 19908 34142
rect 20300 34132 20356 34142
rect 19852 34130 20356 34132
rect 19852 34078 19854 34130
rect 19906 34078 20302 34130
rect 20354 34078 20356 34130
rect 19852 34076 20356 34078
rect 19852 34066 19908 34076
rect 19516 33842 19572 33852
rect 18956 33458 19124 33460
rect 18956 33406 18958 33458
rect 19010 33406 19124 33458
rect 18956 33404 19124 33406
rect 19852 33796 19908 33806
rect 18956 33394 19012 33404
rect 19852 33346 19908 33740
rect 19852 33294 19854 33346
rect 19906 33294 19908 33346
rect 19852 33124 19908 33294
rect 20188 33460 20244 33470
rect 20188 33346 20244 33404
rect 20300 33458 20356 34076
rect 20524 34130 20580 34142
rect 20524 34078 20526 34130
rect 20578 34078 20580 34130
rect 20524 33908 20580 34078
rect 20972 34132 21028 34142
rect 20972 34130 21252 34132
rect 20972 34078 20974 34130
rect 21026 34078 21252 34130
rect 20972 34076 21252 34078
rect 20972 34066 21028 34076
rect 20524 33842 20580 33852
rect 20300 33406 20302 33458
rect 20354 33406 20356 33458
rect 20300 33394 20356 33406
rect 20188 33294 20190 33346
rect 20242 33294 20244 33346
rect 20188 33282 20244 33294
rect 21196 33346 21252 34076
rect 21420 34020 21476 34300
rect 21532 34242 21588 34860
rect 21644 34850 21700 34860
rect 21756 34916 21812 34926
rect 21756 34354 21812 34860
rect 21868 34804 21924 34814
rect 21868 34802 22036 34804
rect 21868 34750 21870 34802
rect 21922 34750 22036 34802
rect 21868 34748 22036 34750
rect 21868 34738 21924 34748
rect 21756 34302 21758 34354
rect 21810 34302 21812 34354
rect 21756 34290 21812 34302
rect 21532 34190 21534 34242
rect 21586 34190 21588 34242
rect 21532 34178 21588 34190
rect 21756 34130 21812 34142
rect 21756 34078 21758 34130
rect 21810 34078 21812 34130
rect 21756 34020 21812 34078
rect 21420 33964 21812 34020
rect 21980 33684 22036 34748
rect 22092 34244 22148 34254
rect 22092 34150 22148 34188
rect 21980 33618 22036 33628
rect 21980 33460 22036 33470
rect 21196 33294 21198 33346
rect 21250 33294 21252 33346
rect 21196 33282 21252 33294
rect 21532 33404 21980 33460
rect 21532 33346 21588 33404
rect 21980 33366 22036 33404
rect 21532 33294 21534 33346
rect 21586 33294 21588 33346
rect 21532 33282 21588 33294
rect 19516 33012 19572 33022
rect 18956 32674 19012 32686
rect 18956 32622 18958 32674
rect 19010 32622 19012 32674
rect 18956 31556 19012 32622
rect 19516 32452 19572 32956
rect 19516 32358 19572 32396
rect 19404 31780 19460 31790
rect 19740 31780 19796 31790
rect 19404 31778 19796 31780
rect 19404 31726 19406 31778
rect 19458 31726 19742 31778
rect 19794 31726 19796 31778
rect 19404 31724 19796 31726
rect 19404 31714 19460 31724
rect 19740 31714 19796 31724
rect 18956 31490 19012 31500
rect 18956 31220 19012 31230
rect 19292 31220 19348 31230
rect 18956 31218 19348 31220
rect 18956 31166 18958 31218
rect 19010 31166 19294 31218
rect 19346 31166 19348 31218
rect 18956 31164 19348 31166
rect 18956 31154 19012 31164
rect 19292 31154 19348 31164
rect 19404 31220 19460 31258
rect 19404 31154 19460 31164
rect 19740 31106 19796 31118
rect 19740 31054 19742 31106
rect 19794 31054 19796 31106
rect 19516 30994 19572 31006
rect 19516 30942 19518 30994
rect 19570 30942 19572 30994
rect 18844 30828 19012 30884
rect 18620 30770 18676 30782
rect 18620 30718 18622 30770
rect 18674 30718 18676 30770
rect 18620 30436 18676 30718
rect 18396 30258 18452 30268
rect 18508 30324 18564 30334
rect 18620 30324 18676 30380
rect 18508 30322 18676 30324
rect 18508 30270 18510 30322
rect 18562 30270 18676 30322
rect 18508 30268 18676 30270
rect 18508 30258 18564 30268
rect 18844 30212 18900 30222
rect 18844 30118 18900 30156
rect 18172 29810 18228 29820
rect 18172 29538 18228 29550
rect 18172 29486 18174 29538
rect 18226 29486 18228 29538
rect 17724 29314 17780 29326
rect 17724 29262 17726 29314
rect 17778 29262 17780 29314
rect 17724 28644 17780 29262
rect 18172 28980 18228 29486
rect 18956 29204 19012 30828
rect 19292 30098 19348 30110
rect 19292 30046 19294 30098
rect 19346 30046 19348 30098
rect 19292 29426 19348 30046
rect 19292 29374 19294 29426
rect 19346 29374 19348 29426
rect 19292 29362 19348 29374
rect 19404 29876 19460 29886
rect 18956 29148 19348 29204
rect 18172 28914 18228 28924
rect 19068 28980 19124 28990
rect 17724 26180 17780 28588
rect 18844 28644 18900 28654
rect 18844 28550 18900 28588
rect 19068 28642 19124 28924
rect 19068 28590 19070 28642
rect 19122 28590 19124 28642
rect 19068 28578 19124 28590
rect 18508 28196 18564 28206
rect 18060 28084 18116 28094
rect 18508 28084 18564 28140
rect 18060 28082 18564 28084
rect 18060 28030 18062 28082
rect 18114 28030 18510 28082
rect 18562 28030 18564 28082
rect 18060 28028 18564 28030
rect 18060 28018 18116 28028
rect 18060 27524 18116 27534
rect 17836 27076 17892 27086
rect 18060 27076 18116 27468
rect 17836 27074 18116 27076
rect 17836 27022 17838 27074
rect 17890 27022 18062 27074
rect 18114 27022 18116 27074
rect 17836 27020 18116 27022
rect 17836 27010 17892 27020
rect 18060 27010 18116 27020
rect 18172 27188 18228 28028
rect 18508 28018 18564 28028
rect 18620 27972 18676 27982
rect 18620 27878 18676 27916
rect 18284 27860 18340 27870
rect 18284 27766 18340 27804
rect 18956 27748 19012 27758
rect 18956 27654 19012 27692
rect 18172 26962 18228 27132
rect 19180 27412 19236 27422
rect 18396 27076 18452 27086
rect 18620 27076 18676 27086
rect 18396 27074 18620 27076
rect 18396 27022 18398 27074
rect 18450 27022 18620 27074
rect 18396 27020 18620 27022
rect 18396 27010 18452 27020
rect 18620 26982 18676 27020
rect 18844 27074 18900 27086
rect 18844 27022 18846 27074
rect 18898 27022 18900 27074
rect 18172 26910 18174 26962
rect 18226 26910 18228 26962
rect 18172 26898 18228 26910
rect 18844 26852 18900 27022
rect 18844 26786 18900 26796
rect 19180 26850 19236 27356
rect 19180 26798 19182 26850
rect 19234 26798 19236 26850
rect 19180 26786 19236 26798
rect 17948 26628 18004 26638
rect 17948 26290 18004 26572
rect 18956 26292 19012 26302
rect 17948 26238 17950 26290
rect 18002 26238 18004 26290
rect 17948 26226 18004 26238
rect 18732 26290 19012 26292
rect 18732 26238 18958 26290
rect 19010 26238 19012 26290
rect 18732 26236 19012 26238
rect 17724 26178 17892 26180
rect 17724 26126 17726 26178
rect 17778 26126 17892 26178
rect 17724 26124 17892 26126
rect 17724 26114 17780 26124
rect 17724 24052 17780 24062
rect 17724 23958 17780 23996
rect 17836 21812 17892 26124
rect 18732 25618 18788 26236
rect 18956 26226 19012 26236
rect 18732 25566 18734 25618
rect 18786 25566 18788 25618
rect 18732 25554 18788 25566
rect 19180 26066 19236 26078
rect 19180 26014 19182 26066
rect 19234 26014 19236 26066
rect 18284 24948 18340 24958
rect 18284 24724 18340 24892
rect 19180 24948 19236 26014
rect 19180 24882 19236 24892
rect 18284 24722 18564 24724
rect 18284 24670 18286 24722
rect 18338 24670 18564 24722
rect 18284 24668 18564 24670
rect 18284 24658 18340 24668
rect 18284 24500 18340 24510
rect 17948 24052 18004 24062
rect 18284 24052 18340 24444
rect 17948 24050 18340 24052
rect 17948 23998 17950 24050
rect 18002 23998 18286 24050
rect 18338 23998 18340 24050
rect 17948 23996 18340 23998
rect 17948 23986 18004 23996
rect 18284 23986 18340 23996
rect 18508 24162 18564 24668
rect 18508 24110 18510 24162
rect 18562 24110 18564 24162
rect 18508 24052 18564 24110
rect 18508 23986 18564 23996
rect 18844 23828 18900 23838
rect 19180 23828 19236 23838
rect 18844 23826 19236 23828
rect 18844 23774 18846 23826
rect 18898 23774 19182 23826
rect 19234 23774 19236 23826
rect 18844 23772 19236 23774
rect 18844 23762 18900 23772
rect 19180 23762 19236 23772
rect 18172 23042 18228 23054
rect 18172 22990 18174 23042
rect 18226 22990 18228 23042
rect 18172 22148 18228 22990
rect 18172 22082 18228 22092
rect 18956 22260 19012 22270
rect 18396 21812 18452 21822
rect 17836 21746 17892 21756
rect 18060 21810 18452 21812
rect 18060 21758 18398 21810
rect 18450 21758 18452 21810
rect 18060 21756 18452 21758
rect 18060 21698 18116 21756
rect 18396 21746 18452 21756
rect 18956 21810 19012 22204
rect 18956 21758 18958 21810
rect 19010 21758 19012 21810
rect 18956 21746 19012 21758
rect 18060 21646 18062 21698
rect 18114 21646 18116 21698
rect 18060 20356 18116 21646
rect 18508 21700 18564 21710
rect 18396 21364 18452 21374
rect 18396 21270 18452 21308
rect 18060 20290 18116 20300
rect 18508 20468 18564 21644
rect 19068 21700 19124 21710
rect 19068 21606 19124 21644
rect 18956 21362 19012 21374
rect 18956 21310 18958 21362
rect 19010 21310 19012 21362
rect 18956 21028 19012 21310
rect 18956 20962 19012 20972
rect 19180 21252 19236 21262
rect 18172 20244 18228 20254
rect 17612 20066 17668 20076
rect 17724 20130 17780 20142
rect 17724 20078 17726 20130
rect 17778 20078 17780 20130
rect 17388 19460 17444 19470
rect 17724 19460 17780 20078
rect 18172 20130 18228 20188
rect 18508 20242 18564 20412
rect 18508 20190 18510 20242
rect 18562 20190 18564 20242
rect 18508 20178 18564 20190
rect 18172 20078 18174 20130
rect 18226 20078 18228 20130
rect 18172 20066 18228 20078
rect 18956 20018 19012 20030
rect 18956 19966 18958 20018
rect 19010 19966 19012 20018
rect 18956 19908 19012 19966
rect 19180 20020 19236 21196
rect 19292 20580 19348 29148
rect 19404 28980 19460 29820
rect 19516 29092 19572 30942
rect 19628 30436 19684 30446
rect 19740 30436 19796 31054
rect 19628 30434 19796 30436
rect 19628 30382 19630 30434
rect 19682 30382 19796 30434
rect 19628 30380 19796 30382
rect 19628 30370 19684 30380
rect 19740 29428 19796 29438
rect 19852 29428 19908 33068
rect 20860 33124 20916 33134
rect 21420 33124 21476 33134
rect 20860 33122 21476 33124
rect 20860 33070 20862 33122
rect 20914 33070 21422 33122
rect 21474 33070 21476 33122
rect 20860 33068 21476 33070
rect 22316 33124 22372 34972
rect 22428 34914 22484 34926
rect 22428 34862 22430 34914
rect 22482 34862 22484 34914
rect 22428 34692 22484 34862
rect 22428 34626 22484 34636
rect 22540 34804 22596 35646
rect 22652 35700 22708 35710
rect 22652 35606 22708 35644
rect 22876 35700 22932 35868
rect 22876 35634 22932 35644
rect 24220 35698 24276 36204
rect 24220 35646 24222 35698
rect 24274 35646 24276 35698
rect 24220 35588 24276 35646
rect 24220 35522 24276 35532
rect 24332 36036 24388 36046
rect 22672 35308 22936 35318
rect 22728 35252 22776 35308
rect 22832 35252 22880 35308
rect 22672 35242 22936 35252
rect 23996 35140 24052 35150
rect 22540 34244 22596 34748
rect 22540 34178 22596 34188
rect 22764 34914 22820 34926
rect 22764 34862 22766 34914
rect 22818 34862 22820 34914
rect 22428 34018 22484 34030
rect 22428 33966 22430 34018
rect 22482 33966 22484 34018
rect 22428 33236 22484 33966
rect 22764 33908 22820 34862
rect 23996 34914 24052 35084
rect 23996 34862 23998 34914
rect 24050 34862 24052 34914
rect 23996 34850 24052 34862
rect 23436 34804 23492 34814
rect 23436 34710 23492 34748
rect 24220 34692 24276 34702
rect 24220 34354 24276 34636
rect 24332 34468 24388 35980
rect 24668 35700 24724 36204
rect 26684 36260 26740 36270
rect 24444 35586 24500 35598
rect 24444 35534 24446 35586
rect 24498 35534 24500 35586
rect 24444 35140 24500 35534
rect 24556 35476 24612 35486
rect 24556 35382 24612 35420
rect 24444 35074 24500 35084
rect 24668 35028 24724 35644
rect 26012 35700 26068 35710
rect 26012 35606 26068 35644
rect 26684 35700 26740 36204
rect 26684 35634 26740 35644
rect 25676 35588 25732 35598
rect 25228 35028 25284 35038
rect 24668 34972 25060 35028
rect 24332 34412 24500 34468
rect 24220 34302 24222 34354
rect 24274 34302 24276 34354
rect 24220 34290 24276 34302
rect 22764 33842 22820 33852
rect 23100 34130 23156 34142
rect 23100 34078 23102 34130
rect 23154 34078 23156 34130
rect 22672 33740 22936 33750
rect 22728 33684 22776 33740
rect 22832 33684 22880 33740
rect 22672 33674 22936 33684
rect 22764 33236 22820 33246
rect 22428 33234 22820 33236
rect 22428 33182 22766 33234
rect 22818 33182 22820 33234
rect 22428 33180 22820 33182
rect 22764 33170 22820 33180
rect 22316 33068 22484 33124
rect 20860 33058 20916 33068
rect 20188 33012 20244 33022
rect 20188 32786 20244 32956
rect 20188 32734 20190 32786
rect 20242 32734 20244 32786
rect 20188 32722 20244 32734
rect 21420 32788 21476 33068
rect 21420 32722 21476 32732
rect 21532 33012 21588 33022
rect 20748 32450 20804 32462
rect 21420 32452 21476 32462
rect 20748 32398 20750 32450
rect 20802 32398 20804 32450
rect 20748 32004 20804 32398
rect 20188 31948 20804 32004
rect 21308 32450 21476 32452
rect 21308 32398 21422 32450
rect 21474 32398 21476 32450
rect 21308 32396 21476 32398
rect 20188 31890 20244 31948
rect 20188 31838 20190 31890
rect 20242 31838 20244 31890
rect 20188 31556 20244 31838
rect 20188 31220 20244 31500
rect 20300 31778 20356 31790
rect 20300 31726 20302 31778
rect 20354 31726 20356 31778
rect 20300 31444 20356 31726
rect 20300 31378 20356 31388
rect 20300 31220 20356 31230
rect 20188 31218 20356 31220
rect 20188 31166 20302 31218
rect 20354 31166 20356 31218
rect 20188 31164 20356 31166
rect 20300 31154 20356 31164
rect 20412 30994 20468 31006
rect 20412 30942 20414 30994
rect 20466 30942 20468 30994
rect 20412 30884 20468 30942
rect 20860 30884 20916 30894
rect 20412 30882 20916 30884
rect 20412 30830 20862 30882
rect 20914 30830 20916 30882
rect 20412 30828 20916 30830
rect 20860 30772 20916 30828
rect 20860 30706 20916 30716
rect 19964 30436 20020 30446
rect 19964 29650 20020 30380
rect 20188 30212 20244 30222
rect 20188 30100 20244 30156
rect 20188 30098 20356 30100
rect 20188 30046 20190 30098
rect 20242 30046 20356 30098
rect 20188 30044 20356 30046
rect 20188 30034 20244 30044
rect 19964 29598 19966 29650
rect 20018 29598 20020 29650
rect 19964 29586 20020 29598
rect 20300 29652 20356 30044
rect 20860 29764 20916 29774
rect 21308 29764 21364 32396
rect 21420 32386 21476 32396
rect 21532 32116 21588 32956
rect 21868 32900 21924 32910
rect 21756 32676 21812 32686
rect 21756 32582 21812 32620
rect 21420 32060 21588 32116
rect 21420 31218 21476 32060
rect 21532 31890 21588 31902
rect 21532 31838 21534 31890
rect 21586 31838 21588 31890
rect 21532 31780 21588 31838
rect 21532 31714 21588 31724
rect 21420 31166 21422 31218
rect 21474 31166 21476 31218
rect 21420 31154 21476 31166
rect 21644 31666 21700 31678
rect 21644 31614 21646 31666
rect 21698 31614 21700 31666
rect 21644 31220 21700 31614
rect 21644 31154 21700 31164
rect 21532 30324 21588 30334
rect 21532 30230 21588 30268
rect 21644 30098 21700 30110
rect 21644 30046 21646 30098
rect 21698 30046 21700 30098
rect 21308 29708 21476 29764
rect 20524 29652 20580 29662
rect 20300 29650 20580 29652
rect 20300 29598 20526 29650
rect 20578 29598 20580 29650
rect 20300 29596 20580 29598
rect 20524 29586 20580 29596
rect 20748 29652 20804 29662
rect 20748 29558 20804 29596
rect 20188 29538 20244 29550
rect 20188 29486 20190 29538
rect 20242 29486 20244 29538
rect 19852 29372 20020 29428
rect 19740 29334 19796 29372
rect 19516 29036 19796 29092
rect 19404 28924 19572 28980
rect 19404 27860 19460 27870
rect 19404 27766 19460 27804
rect 19516 27524 19572 28924
rect 19740 28754 19796 29036
rect 19740 28702 19742 28754
rect 19794 28702 19796 28754
rect 19740 28532 19796 28702
rect 19740 28466 19796 28476
rect 19852 27748 19908 27758
rect 19852 27654 19908 27692
rect 19516 27468 19908 27524
rect 19516 27076 19572 27086
rect 19516 26962 19572 27020
rect 19516 26910 19518 26962
rect 19570 26910 19572 26962
rect 19404 25508 19460 25518
rect 19516 25508 19572 26910
rect 19740 27074 19796 27086
rect 19740 27022 19742 27074
rect 19794 27022 19796 27074
rect 19740 26908 19796 27022
rect 19628 26852 19796 26908
rect 19628 26292 19684 26796
rect 19628 25618 19684 26236
rect 19628 25566 19630 25618
rect 19682 25566 19684 25618
rect 19628 25554 19684 25566
rect 19404 25506 19572 25508
rect 19404 25454 19406 25506
rect 19458 25454 19572 25506
rect 19404 25452 19572 25454
rect 19404 25442 19460 25452
rect 19628 24724 19684 24734
rect 19516 24668 19628 24724
rect 19516 23938 19572 24668
rect 19628 24630 19684 24668
rect 19740 24610 19796 24622
rect 19740 24558 19742 24610
rect 19794 24558 19796 24610
rect 19740 24500 19796 24558
rect 19740 24434 19796 24444
rect 19628 24052 19684 24062
rect 19628 23958 19684 23996
rect 19516 23886 19518 23938
rect 19570 23886 19572 23938
rect 19516 23874 19572 23886
rect 19740 23826 19796 23838
rect 19740 23774 19742 23826
rect 19794 23774 19796 23826
rect 19740 23716 19796 23774
rect 19740 23650 19796 23660
rect 19404 22260 19460 22270
rect 19404 22166 19460 22204
rect 19516 21588 19572 21598
rect 19516 21586 19796 21588
rect 19516 21534 19518 21586
rect 19570 21534 19796 21586
rect 19516 21532 19796 21534
rect 19516 21522 19572 21532
rect 19516 21028 19572 21038
rect 19516 20914 19572 20972
rect 19516 20862 19518 20914
rect 19570 20862 19572 20914
rect 19516 20850 19572 20862
rect 19740 20916 19796 21532
rect 19852 21028 19908 27468
rect 19964 21252 20020 29372
rect 20076 28980 20132 28990
rect 20076 28532 20132 28924
rect 20188 28756 20244 29486
rect 20860 29538 20916 29708
rect 21196 29652 21252 29662
rect 21252 29596 21364 29652
rect 21196 29586 21252 29596
rect 20860 29486 20862 29538
rect 20914 29486 20916 29538
rect 20860 29474 20916 29486
rect 21308 29538 21364 29596
rect 21308 29486 21310 29538
rect 21362 29486 21364 29538
rect 21308 29474 21364 29486
rect 20188 28690 20244 28700
rect 20300 29426 20356 29438
rect 21196 29428 21252 29438
rect 20300 29374 20302 29426
rect 20354 29374 20356 29426
rect 20300 29316 20356 29374
rect 20972 29426 21252 29428
rect 20972 29374 21198 29426
rect 21250 29374 21252 29426
rect 20972 29372 21252 29374
rect 20972 29316 21028 29372
rect 21196 29362 21252 29372
rect 20300 29260 21028 29316
rect 21308 29316 21364 29326
rect 20188 28532 20244 28542
rect 20076 28530 20244 28532
rect 20076 28478 20190 28530
rect 20242 28478 20244 28530
rect 20076 28476 20244 28478
rect 20188 28466 20244 28476
rect 20300 28084 20356 29260
rect 20636 28980 20692 28990
rect 20636 28754 20692 28924
rect 21308 28756 21364 29260
rect 20636 28702 20638 28754
rect 20690 28702 20692 28754
rect 20188 28028 20356 28084
rect 20524 28532 20580 28542
rect 20524 28082 20580 28476
rect 20524 28030 20526 28082
rect 20578 28030 20580 28082
rect 20188 27972 20244 28028
rect 20524 28018 20580 28030
rect 20076 27860 20132 27870
rect 20076 27298 20132 27804
rect 20076 27246 20078 27298
rect 20130 27246 20132 27298
rect 20076 27234 20132 27246
rect 20188 26908 20244 27916
rect 20300 27858 20356 27870
rect 20300 27806 20302 27858
rect 20354 27806 20356 27858
rect 20300 27412 20356 27806
rect 20412 27748 20468 27758
rect 20412 27654 20468 27692
rect 20300 27346 20356 27356
rect 20636 26908 20692 28702
rect 21196 28700 21364 28756
rect 21196 28642 21252 28700
rect 21420 28644 21476 29708
rect 21532 29652 21588 29662
rect 21644 29652 21700 30046
rect 21868 29988 21924 32844
rect 21868 29922 21924 29932
rect 22316 31106 22372 31118
rect 22316 31054 22318 31106
rect 22370 31054 22372 31106
rect 21868 29764 21924 29774
rect 21532 29650 21700 29652
rect 21532 29598 21534 29650
rect 21586 29598 21700 29650
rect 21532 29596 21700 29598
rect 21756 29652 21812 29662
rect 21532 29586 21588 29596
rect 21196 28590 21198 28642
rect 21250 28590 21252 28642
rect 21196 28578 21252 28590
rect 21308 28588 21476 28644
rect 21756 28644 21812 29596
rect 21868 29314 21924 29708
rect 21868 29262 21870 29314
rect 21922 29262 21924 29314
rect 21868 29092 21924 29262
rect 22316 29316 22372 31054
rect 22316 29250 22372 29260
rect 22428 30772 22484 33068
rect 23100 32900 23156 34078
rect 23996 34130 24052 34142
rect 23996 34078 23998 34130
rect 24050 34078 24052 34130
rect 23324 34020 23380 34030
rect 23324 33926 23380 33964
rect 23996 33908 24052 34078
rect 23996 33842 24052 33852
rect 24108 34018 24164 34030
rect 24108 33966 24110 34018
rect 24162 33966 24164 34018
rect 23100 32834 23156 32844
rect 23212 33346 23268 33358
rect 23212 33294 23214 33346
rect 23266 33294 23268 33346
rect 23212 32786 23268 33294
rect 24108 33346 24164 33966
rect 24108 33294 24110 33346
rect 24162 33294 24164 33346
rect 24108 33282 24164 33294
rect 24444 33796 24500 34412
rect 24556 34130 24612 34142
rect 24556 34078 24558 34130
rect 24610 34078 24612 34130
rect 24556 34018 24612 34078
rect 24556 33966 24558 34018
rect 24610 33966 24612 34018
rect 24556 33954 24612 33966
rect 24780 34020 24836 34030
rect 24780 34018 24948 34020
rect 24780 33966 24782 34018
rect 24834 33966 24948 34018
rect 24780 33964 24948 33966
rect 24780 33954 24836 33964
rect 24332 33122 24388 33134
rect 24332 33070 24334 33122
rect 24386 33070 24388 33122
rect 23212 32734 23214 32786
rect 23266 32734 23268 32786
rect 23212 32722 23268 32734
rect 23884 32900 23940 32910
rect 23884 32786 23940 32844
rect 23884 32734 23886 32786
rect 23938 32734 23940 32786
rect 23884 32722 23940 32734
rect 23100 32674 23156 32686
rect 23100 32622 23102 32674
rect 23154 32622 23156 32674
rect 22672 32172 22936 32182
rect 22728 32116 22776 32172
rect 22832 32116 22880 32172
rect 22672 32106 22936 32116
rect 23100 31556 23156 32622
rect 24332 32004 24388 33070
rect 24444 32786 24500 33740
rect 24892 33346 24948 33964
rect 24892 33294 24894 33346
rect 24946 33294 24948 33346
rect 24892 33282 24948 33294
rect 24444 32734 24446 32786
rect 24498 32734 24500 32786
rect 24444 32722 24500 32734
rect 24332 31938 24388 31948
rect 23324 31668 23380 31678
rect 23324 31666 23940 31668
rect 23324 31614 23326 31666
rect 23378 31614 23940 31666
rect 23324 31612 23940 31614
rect 23324 31602 23380 31612
rect 23212 31556 23268 31566
rect 23100 31554 23268 31556
rect 23100 31502 23214 31554
rect 23266 31502 23268 31554
rect 23100 31500 23268 31502
rect 23212 31490 23268 31500
rect 23884 31218 23940 31612
rect 23884 31166 23886 31218
rect 23938 31166 23940 31218
rect 23884 31154 23940 31166
rect 24108 31554 24164 31566
rect 24108 31502 24110 31554
rect 24162 31502 24164 31554
rect 23996 31106 24052 31118
rect 23996 31054 23998 31106
rect 24050 31054 24052 31106
rect 22876 30996 22932 31006
rect 23996 30996 24052 31054
rect 22876 30994 23156 30996
rect 22876 30942 22878 30994
rect 22930 30942 23156 30994
rect 22876 30940 23156 30942
rect 22876 30930 22932 30940
rect 21868 29036 22148 29092
rect 22092 28980 22148 29036
rect 22092 28924 22260 28980
rect 21980 28866 22036 28878
rect 21980 28814 21982 28866
rect 22034 28814 22036 28866
rect 21980 28756 22036 28814
rect 21980 28690 22036 28700
rect 21756 28588 21924 28644
rect 20860 27860 20916 27870
rect 20860 27766 20916 27804
rect 21308 27076 21364 28588
rect 21532 28530 21588 28542
rect 21532 28478 21534 28530
rect 21586 28478 21588 28530
rect 21420 28420 21476 28430
rect 21420 28326 21476 28364
rect 21532 27748 21588 28478
rect 21868 28532 21924 28588
rect 21980 28532 22036 28542
rect 21868 28530 22036 28532
rect 21868 28478 21982 28530
rect 22034 28478 22036 28530
rect 21868 28476 22036 28478
rect 21980 28466 22036 28476
rect 22092 28532 22148 28542
rect 21756 27748 21812 27758
rect 21532 27746 21812 27748
rect 21532 27694 21758 27746
rect 21810 27694 21812 27746
rect 21532 27692 21812 27694
rect 21756 27076 21812 27692
rect 22092 27636 22148 28476
rect 22204 27860 22260 28924
rect 22316 28420 22372 28430
rect 22316 28082 22372 28364
rect 22316 28030 22318 28082
rect 22370 28030 22372 28082
rect 22316 28018 22372 28030
rect 22204 27858 22372 27860
rect 22204 27806 22206 27858
rect 22258 27806 22372 27858
rect 22204 27804 22372 27806
rect 22204 27794 22260 27804
rect 22316 27748 22372 27804
rect 22092 27580 22260 27636
rect 22092 27300 22148 27310
rect 21980 27076 22036 27086
rect 22092 27076 22148 27244
rect 21308 27020 21700 27076
rect 21756 27020 21924 27076
rect 21644 26908 21700 27020
rect 20188 26852 20468 26908
rect 20188 26628 20244 26638
rect 20188 25284 20244 26572
rect 20300 26292 20356 26302
rect 20300 26198 20356 26236
rect 20188 25282 20356 25284
rect 20188 25230 20190 25282
rect 20242 25230 20356 25282
rect 20188 25228 20356 25230
rect 20188 25218 20244 25228
rect 20300 23716 20356 25228
rect 20300 23650 20356 23660
rect 20300 23044 20356 23054
rect 20188 23042 20356 23044
rect 20188 22990 20302 23042
rect 20354 22990 20356 23042
rect 20188 22988 20356 22990
rect 19964 21186 20020 21196
rect 20076 22148 20132 22158
rect 19852 20972 20020 21028
rect 19740 20850 19796 20860
rect 19852 20692 19908 20702
rect 19740 20690 19908 20692
rect 19740 20638 19854 20690
rect 19906 20638 19908 20690
rect 19740 20636 19908 20638
rect 19292 20524 19684 20580
rect 19516 20356 19572 20366
rect 19292 20244 19348 20254
rect 19292 20150 19348 20188
rect 19180 19964 19348 20020
rect 17836 19796 17892 19806
rect 17836 19702 17892 19740
rect 17388 19458 18452 19460
rect 17388 19406 17390 19458
rect 17442 19406 18452 19458
rect 17388 19404 18452 19406
rect 17388 19394 17444 19404
rect 17052 16818 17108 16828
rect 17164 19348 17220 19358
rect 17164 19012 17220 19292
rect 17276 19236 17332 19246
rect 17276 19142 17332 19180
rect 17164 17780 17220 18956
rect 17612 19124 17668 19134
rect 17500 18788 17556 18798
rect 17500 18340 17556 18732
rect 17612 18564 17668 19068
rect 17724 19012 17780 19022
rect 17724 18918 17780 18956
rect 17948 19012 18004 19022
rect 17948 19010 18116 19012
rect 17948 18958 17950 19010
rect 18002 18958 18116 19010
rect 17948 18956 18116 18958
rect 17948 18946 18004 18956
rect 17612 18508 17780 18564
rect 17612 18340 17668 18350
rect 17500 18338 17668 18340
rect 17500 18286 17614 18338
rect 17666 18286 17668 18338
rect 17500 18284 17668 18286
rect 17612 18274 17668 18284
rect 17276 17780 17332 17790
rect 17164 17778 17332 17780
rect 17164 17726 17278 17778
rect 17330 17726 17332 17778
rect 17164 17724 17332 17726
rect 16940 15922 16996 15932
rect 17164 15540 17220 17724
rect 17276 17714 17332 17724
rect 17724 17668 17780 18508
rect 17948 18452 18004 18462
rect 17948 18358 18004 18396
rect 18060 18340 18116 18956
rect 18060 18274 18116 18284
rect 17724 17666 18228 17668
rect 17724 17614 17726 17666
rect 17778 17614 18228 17666
rect 17724 17612 18228 17614
rect 17724 17602 17780 17612
rect 18172 17556 18228 17612
rect 18172 17500 18340 17556
rect 17836 17442 17892 17454
rect 17836 17390 17838 17442
rect 17890 17390 17892 17442
rect 17836 16996 17892 17390
rect 18060 17444 18116 17454
rect 18060 17350 18116 17388
rect 17836 16930 17892 16940
rect 18172 17108 18228 17118
rect 18172 16994 18228 17052
rect 18172 16942 18174 16994
rect 18226 16942 18228 16994
rect 18172 16930 18228 16942
rect 17164 15474 17220 15484
rect 17500 16882 17556 16894
rect 17500 16830 17502 16882
rect 17554 16830 17556 16882
rect 16716 15362 16772 15372
rect 16828 15202 16884 15214
rect 16828 15150 16830 15202
rect 16882 15150 16884 15202
rect 16828 15148 16884 15150
rect 16604 15092 16772 15148
rect 16828 15092 16996 15148
rect 16604 14532 16660 14542
rect 16380 14530 16660 14532
rect 16380 14478 16606 14530
rect 16658 14478 16660 14530
rect 16380 14476 16660 14478
rect 16268 14420 16324 14430
rect 16268 14326 16324 14364
rect 16380 14308 16436 14318
rect 16380 14214 16436 14252
rect 16044 13694 16046 13746
rect 16098 13694 16100 13746
rect 16044 13682 16100 13694
rect 16156 14196 16212 14206
rect 15036 13522 15316 13524
rect 15036 13470 15038 13522
rect 15090 13470 15316 13522
rect 15036 13468 15316 13470
rect 15708 13522 15764 13534
rect 15708 13470 15710 13522
rect 15762 13470 15764 13522
rect 15036 13458 15092 13468
rect 14924 13244 15316 13300
rect 15260 13186 15316 13244
rect 15260 13134 15262 13186
rect 15314 13134 15316 13186
rect 15260 13122 15316 13134
rect 15372 13188 15428 13198
rect 15260 12964 15316 12974
rect 15372 12964 15428 13132
rect 15260 12962 15428 12964
rect 15260 12910 15262 12962
rect 15314 12910 15428 12962
rect 15260 12908 15428 12910
rect 14252 12740 14308 12750
rect 14252 12646 14308 12684
rect 14812 12738 14868 12750
rect 14812 12686 14814 12738
rect 14866 12686 14868 12738
rect 14476 12066 14532 12078
rect 14476 12014 14478 12066
rect 14530 12014 14532 12066
rect 13916 11732 14196 11788
rect 14140 11620 14196 11732
rect 14140 11554 14196 11564
rect 14364 11732 14420 11742
rect 14364 11396 14420 11676
rect 14364 11302 14420 11340
rect 13468 11282 13636 11284
rect 13468 11230 13470 11282
rect 13522 11230 13636 11282
rect 13468 11228 13636 11230
rect 12684 10388 12740 10444
rect 12460 10332 12740 10388
rect 12460 9938 12516 10332
rect 12460 9886 12462 9938
rect 12514 9886 12516 9938
rect 12012 9604 12068 9614
rect 12012 9510 12068 9548
rect 12460 8484 12516 9886
rect 12012 8428 12460 8484
rect 11900 8370 11956 8382
rect 11900 8318 11902 8370
rect 11954 8318 11956 8370
rect 11900 8260 11956 8318
rect 11900 8194 11956 8204
rect 11900 6468 11956 6478
rect 11788 6466 11956 6468
rect 11788 6414 11902 6466
rect 11954 6414 11956 6466
rect 11788 6412 11956 6414
rect 11340 6300 11732 6356
rect 11228 6188 11396 6244
rect 11116 6132 11172 6142
rect 11116 6018 11172 6076
rect 11116 5966 11118 6018
rect 11170 5966 11172 6018
rect 11116 5908 11172 5966
rect 11228 6020 11284 6030
rect 11228 5926 11284 5964
rect 11116 5842 11172 5852
rect 11228 5684 11284 5694
rect 11004 5070 11006 5122
rect 11058 5070 11060 5122
rect 11004 5058 11060 5070
rect 11116 5682 11284 5684
rect 11116 5630 11230 5682
rect 11282 5630 11284 5682
rect 11116 5628 11284 5630
rect 11004 4900 11060 4910
rect 10668 4386 10724 4396
rect 10892 4450 10948 4462
rect 10892 4398 10894 4450
rect 10946 4398 10948 4450
rect 10220 4174 10222 4226
rect 10274 4174 10276 4226
rect 10220 4162 10276 4174
rect 10556 4338 10612 4350
rect 10556 4286 10558 4338
rect 10610 4286 10612 4338
rect 8876 3836 9380 3892
rect 9324 3666 9380 3836
rect 10556 3780 10612 4286
rect 10892 4004 10948 4398
rect 10892 3938 10948 3948
rect 10556 3714 10612 3724
rect 9324 3614 9326 3666
rect 9378 3614 9380 3666
rect 9324 3602 9380 3614
rect 7868 3442 8036 3444
rect 7868 3390 7870 3442
rect 7922 3390 8036 3442
rect 7868 3388 8036 3390
rect 8092 3554 8148 3566
rect 8092 3502 8094 3554
rect 8146 3502 8148 3554
rect 8092 3444 8148 3502
rect 7868 3378 7924 3388
rect 7756 3266 7812 3276
rect 2716 3164 3220 3220
rect 2716 800 2772 3164
rect 8092 2212 8148 3388
rect 8876 3444 8932 3482
rect 8876 3378 8932 3388
rect 11004 2324 11060 4844
rect 11116 2548 11172 5628
rect 11228 5618 11284 5628
rect 11340 5012 11396 6188
rect 11340 4946 11396 4956
rect 11228 4898 11284 4910
rect 11228 4846 11230 4898
rect 11282 4846 11284 4898
rect 11228 3444 11284 4846
rect 11340 4788 11396 4798
rect 11340 4562 11396 4732
rect 11340 4510 11342 4562
rect 11394 4510 11396 4562
rect 11340 4498 11396 4510
rect 11452 4340 11508 4350
rect 11452 4246 11508 4284
rect 11452 4116 11508 4126
rect 11452 3666 11508 4060
rect 11564 4114 11620 4126
rect 11564 4062 11566 4114
rect 11618 4062 11620 4114
rect 11564 4004 11620 4062
rect 11564 3938 11620 3948
rect 11452 3614 11454 3666
rect 11506 3614 11508 3666
rect 11452 3602 11508 3614
rect 11228 2996 11284 3388
rect 11228 2930 11284 2940
rect 11676 2772 11732 6300
rect 11788 4676 11844 6412
rect 11900 6402 11956 6412
rect 11900 6020 11956 6030
rect 11900 5926 11956 5964
rect 11788 4610 11844 4620
rect 12012 5234 12068 8428
rect 12460 8418 12516 8428
rect 12572 10164 12628 10174
rect 12460 8260 12516 8270
rect 12572 8260 12628 10108
rect 12796 9940 12852 9950
rect 12796 9846 12852 9884
rect 12908 9714 12964 9726
rect 12908 9662 12910 9714
rect 12962 9662 12964 9714
rect 12908 9044 12964 9662
rect 13132 9044 13188 9054
rect 12908 8988 13132 9044
rect 13132 8930 13188 8988
rect 13132 8878 13134 8930
rect 13186 8878 13188 8930
rect 13132 8866 13188 8878
rect 12460 8258 12628 8260
rect 12460 8206 12462 8258
rect 12514 8206 12628 8258
rect 12460 8204 12628 8206
rect 13020 8820 13076 8830
rect 13020 8258 13076 8764
rect 13020 8206 13022 8258
rect 13074 8206 13076 8258
rect 12460 8194 12516 8204
rect 13020 8194 13076 8206
rect 13356 8372 13412 8382
rect 12684 8148 12740 8158
rect 12684 8054 12740 8092
rect 12796 8036 12852 8046
rect 12796 7942 12852 7980
rect 13356 7924 13412 8316
rect 13244 7868 13356 7924
rect 12460 7362 12516 7374
rect 12460 7310 12462 7362
rect 12514 7310 12516 7362
rect 12124 6692 12180 6702
rect 12124 6020 12180 6636
rect 12236 6692 12292 6702
rect 12460 6692 12516 7310
rect 13244 7362 13300 7868
rect 13356 7858 13412 7868
rect 13244 7310 13246 7362
rect 13298 7310 13300 7362
rect 13244 7298 13300 7310
rect 13468 7140 13524 11228
rect 13804 11172 13860 11182
rect 14476 11172 14532 12014
rect 14812 12068 14868 12686
rect 14812 12002 14868 12012
rect 15036 12738 15092 12750
rect 15036 12686 15038 12738
rect 15090 12686 15092 12738
rect 15036 11506 15092 12686
rect 15260 12180 15316 12908
rect 15596 12852 15652 12862
rect 15596 12758 15652 12796
rect 15708 12740 15764 13470
rect 15820 13412 15876 13422
rect 15820 12962 15876 13356
rect 16156 13076 16212 14140
rect 16492 13970 16548 13982
rect 16492 13918 16494 13970
rect 16546 13918 16548 13970
rect 16268 13748 16324 13758
rect 16268 13522 16324 13692
rect 16268 13470 16270 13522
rect 16322 13470 16324 13522
rect 16268 13458 16324 13470
rect 16156 13010 16212 13020
rect 16380 13412 16436 13422
rect 15820 12910 15822 12962
rect 15874 12910 15876 12962
rect 15820 12898 15876 12910
rect 16380 12962 16436 13356
rect 16492 13076 16548 13918
rect 16604 13972 16660 14476
rect 16604 13906 16660 13916
rect 16604 13748 16660 13758
rect 16604 13654 16660 13692
rect 16604 13076 16660 13086
rect 16492 13020 16604 13076
rect 16604 13010 16660 13020
rect 16380 12910 16382 12962
rect 16434 12910 16436 12962
rect 16380 12898 16436 12910
rect 15708 12674 15764 12684
rect 16492 12852 16548 12862
rect 16492 12628 16548 12796
rect 15518 12572 15782 12582
rect 15574 12516 15622 12572
rect 15678 12516 15726 12572
rect 15518 12506 15782 12516
rect 15820 12404 15876 12414
rect 15596 12292 15652 12302
rect 15596 12198 15652 12236
rect 15820 12290 15876 12348
rect 15820 12238 15822 12290
rect 15874 12238 15876 12290
rect 15820 12226 15876 12238
rect 15260 12114 15316 12124
rect 16492 12178 16548 12572
rect 16492 12126 16494 12178
rect 16546 12126 16548 12178
rect 16492 12114 16548 12126
rect 16604 12068 16660 12078
rect 16604 11974 16660 12012
rect 15036 11454 15038 11506
rect 15090 11454 15092 11506
rect 15036 11442 15092 11454
rect 13804 11170 14532 11172
rect 13804 11118 13806 11170
rect 13858 11118 14532 11170
rect 13804 11116 14532 11118
rect 13580 10722 13636 10734
rect 13580 10670 13582 10722
rect 13634 10670 13636 10722
rect 13580 10612 13636 10670
rect 13580 10546 13636 10556
rect 13580 9044 13636 9054
rect 13580 9042 13748 9044
rect 13580 8990 13582 9042
rect 13634 8990 13748 9042
rect 13580 8988 13748 8990
rect 13580 8978 13636 8988
rect 13692 8372 13748 8988
rect 13804 8596 13860 11116
rect 15518 11004 15782 11014
rect 15574 10948 15622 11004
rect 15678 10948 15726 11004
rect 15518 10938 15782 10948
rect 15932 10836 15988 10846
rect 14700 10722 14756 10734
rect 14700 10670 14702 10722
rect 14754 10670 14756 10722
rect 14252 10610 14308 10622
rect 14252 10558 14254 10610
rect 14306 10558 14308 10610
rect 13916 9940 13972 9950
rect 13916 9714 13972 9884
rect 13916 9662 13918 9714
rect 13970 9662 13972 9714
rect 13916 9650 13972 9662
rect 14252 9604 14308 10558
rect 14476 10388 14532 10398
rect 13916 9044 13972 9054
rect 13916 8950 13972 8988
rect 14252 8708 14308 9548
rect 14252 8642 14308 8652
rect 14364 10164 14420 10174
rect 13804 8530 13860 8540
rect 14364 8372 14420 10108
rect 14476 9826 14532 10332
rect 14476 9774 14478 9826
rect 14530 9774 14532 9826
rect 14476 9762 14532 9774
rect 14700 9044 14756 10670
rect 14700 8978 14756 8988
rect 14924 10610 14980 10622
rect 14924 10558 14926 10610
rect 14978 10558 14980 10610
rect 14924 8372 14980 10558
rect 15260 10500 15316 10510
rect 15260 10406 15316 10444
rect 15932 10498 15988 10780
rect 15932 10446 15934 10498
rect 15986 10446 15988 10498
rect 15148 9826 15204 9838
rect 15148 9774 15150 9826
rect 15202 9774 15204 9826
rect 15036 9716 15092 9726
rect 15036 9154 15092 9660
rect 15036 9102 15038 9154
rect 15090 9102 15092 9154
rect 15036 9090 15092 9102
rect 15148 8820 15204 9774
rect 15932 9828 15988 10446
rect 16380 10836 16436 10846
rect 16380 10276 16436 10780
rect 16380 10210 16436 10220
rect 16716 10052 16772 15092
rect 16828 13746 16884 13758
rect 16828 13694 16830 13746
rect 16882 13694 16884 13746
rect 16828 13524 16884 13694
rect 16828 13458 16884 13468
rect 16828 12180 16884 12190
rect 16940 12180 16996 15092
rect 17052 14644 17108 14654
rect 17108 14588 17444 14644
rect 17052 14550 17108 14588
rect 17388 13746 17444 14588
rect 17388 13694 17390 13746
rect 17442 13694 17444 13746
rect 17388 13682 17444 13694
rect 17500 13412 17556 16830
rect 18060 16884 18116 16894
rect 17724 16212 17780 16222
rect 17724 16118 17780 16156
rect 17612 15540 17668 15550
rect 17612 15446 17668 15484
rect 18060 15538 18116 16828
rect 18284 16098 18340 17500
rect 18284 16046 18286 16098
rect 18338 16046 18340 16098
rect 18284 16034 18340 16046
rect 18396 15986 18452 19404
rect 18956 19236 19012 19852
rect 19180 19796 19236 19806
rect 19180 19702 19236 19740
rect 18956 19170 19012 19180
rect 19068 19234 19124 19246
rect 19068 19182 19070 19234
rect 19122 19182 19124 19234
rect 18732 19012 18788 19022
rect 18732 18918 18788 18956
rect 19068 18788 19124 19182
rect 19068 18722 19124 18732
rect 19292 18676 19348 19964
rect 19404 20018 19460 20030
rect 19404 19966 19406 20018
rect 19458 19966 19460 20018
rect 19404 19012 19460 19966
rect 19404 18946 19460 18956
rect 19516 19234 19572 20300
rect 19516 19182 19518 19234
rect 19570 19182 19572 19234
rect 19516 18900 19572 19182
rect 19516 18834 19572 18844
rect 19292 18620 19460 18676
rect 18844 18508 19012 18564
rect 18508 18450 18564 18462
rect 18508 18398 18510 18450
rect 18562 18398 18564 18450
rect 18508 16548 18564 18398
rect 18844 18450 18900 18508
rect 18844 18398 18846 18450
rect 18898 18398 18900 18450
rect 18844 18340 18900 18398
rect 18956 18452 19012 18508
rect 19292 18452 19348 18462
rect 18956 18450 19348 18452
rect 18956 18398 19294 18450
rect 19346 18398 19348 18450
rect 18956 18396 19348 18398
rect 19292 18386 19348 18396
rect 18620 18284 18900 18340
rect 18620 17778 18676 18284
rect 19404 18228 19460 18620
rect 19628 18338 19684 20524
rect 19740 20468 19796 20636
rect 19852 20626 19908 20636
rect 19740 20130 19796 20412
rect 19740 20078 19742 20130
rect 19794 20078 19796 20130
rect 19740 20066 19796 20078
rect 19852 19572 19908 19582
rect 19852 19346 19908 19516
rect 19852 19294 19854 19346
rect 19906 19294 19908 19346
rect 19852 19282 19908 19294
rect 19628 18286 19630 18338
rect 19682 18286 19684 18338
rect 19628 18274 19684 18286
rect 19740 18562 19796 18574
rect 19740 18510 19742 18562
rect 19794 18510 19796 18562
rect 18620 17726 18622 17778
rect 18674 17726 18676 17778
rect 18620 17714 18676 17726
rect 18732 18172 19460 18228
rect 18620 16548 18676 16558
rect 18508 16492 18620 16548
rect 18620 16482 18676 16492
rect 18396 15934 18398 15986
rect 18450 15934 18452 15986
rect 18396 15876 18452 15934
rect 18396 15764 18452 15820
rect 18060 15486 18062 15538
rect 18114 15486 18116 15538
rect 18060 15474 18116 15486
rect 18284 15708 18452 15764
rect 18620 15874 18676 15886
rect 18620 15822 18622 15874
rect 18674 15822 18676 15874
rect 17724 15204 17780 15214
rect 17724 14530 17780 15148
rect 17724 14478 17726 14530
rect 17778 14478 17780 14530
rect 17724 14466 17780 14478
rect 18284 14532 18340 15708
rect 18396 15428 18452 15438
rect 18396 14642 18452 15372
rect 18620 15092 18676 15822
rect 18620 15026 18676 15036
rect 18396 14590 18398 14642
rect 18450 14590 18452 14642
rect 18396 14578 18452 14590
rect 18284 14466 18340 14476
rect 17612 14308 17668 14318
rect 17612 13522 17668 14252
rect 17948 13746 18004 13758
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 17948 13636 18004 13694
rect 18172 13746 18228 13758
rect 18172 13694 18174 13746
rect 18226 13694 18228 13746
rect 17948 13570 18004 13580
rect 18060 13634 18116 13646
rect 18060 13582 18062 13634
rect 18114 13582 18116 13634
rect 17612 13470 17614 13522
rect 17666 13470 17668 13522
rect 17612 13458 17668 13470
rect 17500 13346 17556 13356
rect 17164 13076 17220 13086
rect 17164 12982 17220 13020
rect 17612 12740 17668 12750
rect 17388 12404 17444 12414
rect 17388 12402 17556 12404
rect 17388 12350 17390 12402
rect 17442 12350 17556 12402
rect 17388 12348 17556 12350
rect 17388 12338 17444 12348
rect 16884 12124 16996 12180
rect 17388 12180 17444 12190
rect 16828 12114 16884 12124
rect 17388 12086 17444 12124
rect 16940 11732 16996 11742
rect 16940 11396 16996 11676
rect 16828 10498 16884 10510
rect 16828 10446 16830 10498
rect 16882 10446 16884 10498
rect 16828 10276 16884 10446
rect 16828 10210 16884 10220
rect 16604 9996 16772 10052
rect 16380 9828 16436 9838
rect 15932 9772 16380 9828
rect 16380 9734 16436 9772
rect 15820 9716 15876 9726
rect 15820 9714 15988 9716
rect 15820 9662 15822 9714
rect 15874 9662 15988 9714
rect 15820 9660 15988 9662
rect 15820 9650 15876 9660
rect 15518 9436 15782 9446
rect 15574 9380 15622 9436
rect 15678 9380 15726 9436
rect 15518 9370 15782 9380
rect 15932 9156 15988 9660
rect 16492 9156 16548 9166
rect 15932 9154 16548 9156
rect 15932 9102 16494 9154
rect 16546 9102 16548 9154
rect 15932 9100 16548 9102
rect 16492 9090 16548 9100
rect 15484 8932 15540 8942
rect 15484 8838 15540 8876
rect 15596 8932 15652 8942
rect 16044 8932 16100 8942
rect 15596 8930 15764 8932
rect 15596 8878 15598 8930
rect 15650 8878 15764 8930
rect 15596 8876 15764 8878
rect 15596 8866 15652 8876
rect 15148 8754 15204 8764
rect 13692 8306 13748 8316
rect 14252 8316 14644 8372
rect 13580 8260 13636 8270
rect 14252 8260 14308 8316
rect 13580 8166 13636 8204
rect 13804 8204 14308 8260
rect 13804 8148 13860 8204
rect 13692 8146 13860 8148
rect 13692 8094 13806 8146
rect 13858 8094 13860 8146
rect 13692 8092 13860 8094
rect 13580 7476 13636 7486
rect 13692 7476 13748 8092
rect 13804 8082 13860 8092
rect 14252 8146 14308 8204
rect 14252 8094 14254 8146
rect 14306 8094 14308 8146
rect 14252 8082 14308 8094
rect 14364 8146 14420 8158
rect 14364 8094 14366 8146
rect 14418 8094 14420 8146
rect 14028 8036 14084 8046
rect 14028 7942 14084 7980
rect 14364 7924 14420 8094
rect 14364 7858 14420 7868
rect 14476 8036 14532 8046
rect 13580 7474 13748 7476
rect 13580 7422 13582 7474
rect 13634 7422 13748 7474
rect 13580 7420 13748 7422
rect 14028 7588 14084 7598
rect 14476 7588 14532 7980
rect 13580 7410 13636 7420
rect 13468 7084 13636 7140
rect 13468 6916 13524 6926
rect 12796 6804 12852 6814
rect 12572 6692 12628 6702
rect 12236 6690 12628 6692
rect 12236 6638 12238 6690
rect 12290 6638 12574 6690
rect 12626 6638 12628 6690
rect 12236 6636 12628 6638
rect 12236 6626 12292 6636
rect 12572 6626 12628 6636
rect 12796 6356 12852 6748
rect 13468 6690 13524 6860
rect 13468 6638 13470 6690
rect 13522 6638 13524 6690
rect 13468 6626 13524 6638
rect 12124 5796 12180 5964
rect 12236 6300 12852 6356
rect 12236 6018 12292 6300
rect 12236 5966 12238 6018
rect 12290 5966 12292 6018
rect 12236 5954 12292 5966
rect 12348 6020 12404 6030
rect 12348 5926 12404 5964
rect 12572 5908 12628 5918
rect 12572 5814 12628 5852
rect 12796 5906 12852 6300
rect 12908 6466 12964 6478
rect 12908 6414 12910 6466
rect 12962 6414 12964 6466
rect 12908 6020 12964 6414
rect 13020 6020 13076 6030
rect 12964 6018 13076 6020
rect 12964 5966 13022 6018
rect 13074 5966 13076 6018
rect 12964 5964 13076 5966
rect 12908 5926 12964 5964
rect 12796 5854 12798 5906
rect 12850 5854 12852 5906
rect 12796 5842 12852 5854
rect 12124 5740 12516 5796
rect 12012 5182 12014 5234
rect 12066 5182 12068 5234
rect 11900 4340 11956 4350
rect 11900 4246 11956 4284
rect 12012 3668 12068 5182
rect 12460 5236 12516 5740
rect 13020 5460 13076 5964
rect 13356 5908 13412 5918
rect 13356 5814 13412 5852
rect 13132 5796 13188 5806
rect 13132 5702 13188 5740
rect 13132 5460 13188 5470
rect 13020 5404 13132 5460
rect 13132 5394 13188 5404
rect 12908 5348 12964 5358
rect 12908 5254 12964 5292
rect 12460 5142 12516 5180
rect 13580 5124 13636 7084
rect 14028 6690 14084 7532
rect 14364 7532 14532 7588
rect 14364 6804 14420 7532
rect 14476 7364 14532 7374
rect 14588 7364 14644 8316
rect 14924 8306 14980 8316
rect 15036 8370 15092 8382
rect 15036 8318 15038 8370
rect 15090 8318 15092 8370
rect 14700 8148 14756 8158
rect 14700 8146 14868 8148
rect 14700 8094 14702 8146
rect 14754 8094 14868 8146
rect 14700 8092 14868 8094
rect 14700 8082 14756 8092
rect 14476 7362 14644 7364
rect 14476 7310 14478 7362
rect 14530 7310 14644 7362
rect 14476 7308 14644 7310
rect 14476 7298 14532 7308
rect 14028 6638 14030 6690
rect 14082 6638 14084 6690
rect 14028 6626 14084 6638
rect 14140 6802 14420 6804
rect 14140 6750 14366 6802
rect 14418 6750 14420 6802
rect 14140 6748 14420 6750
rect 14140 6468 14196 6748
rect 14364 6738 14420 6748
rect 14700 7250 14756 7262
rect 14700 7198 14702 7250
rect 14754 7198 14756 7250
rect 14700 6804 14756 7198
rect 14700 6738 14756 6748
rect 13916 6412 14196 6468
rect 13916 6130 13972 6412
rect 13916 6078 13918 6130
rect 13970 6078 13972 6130
rect 13916 6066 13972 6078
rect 14476 6132 14532 6142
rect 14476 6038 14532 6076
rect 14812 6132 14868 8092
rect 14924 8034 14980 8046
rect 14924 7982 14926 8034
rect 14978 7982 14980 8034
rect 14924 6356 14980 7982
rect 15036 7924 15092 8318
rect 15708 8260 15764 8876
rect 15708 8194 15764 8204
rect 15260 8148 15316 8158
rect 15260 8054 15316 8092
rect 15596 8148 15652 8158
rect 15596 8054 15652 8092
rect 15932 8148 15988 8158
rect 15484 8036 15540 8046
rect 15372 8034 15540 8036
rect 15372 7982 15486 8034
rect 15538 7982 15540 8034
rect 15372 7980 15540 7982
rect 15036 7868 15316 7924
rect 15036 7700 15092 7710
rect 15036 7606 15092 7644
rect 15260 7140 15316 7868
rect 15372 7588 15428 7980
rect 15484 7970 15540 7980
rect 15518 7868 15782 7878
rect 15574 7812 15622 7868
rect 15678 7812 15726 7868
rect 15518 7802 15782 7812
rect 15372 7522 15428 7532
rect 15932 7588 15988 8092
rect 15932 7522 15988 7532
rect 15932 7362 15988 7374
rect 15932 7310 15934 7362
rect 15986 7310 15988 7362
rect 15260 7074 15316 7084
rect 15372 7250 15428 7262
rect 15372 7198 15374 7250
rect 15426 7198 15428 7250
rect 15372 7028 15428 7198
rect 15708 7252 15764 7262
rect 15708 7158 15764 7196
rect 15372 6962 15428 6972
rect 14924 6290 14980 6300
rect 15148 6804 15204 6814
rect 15148 6466 15204 6748
rect 15484 6804 15540 6814
rect 15484 6690 15540 6748
rect 15484 6638 15486 6690
rect 15538 6638 15540 6690
rect 15484 6626 15540 6638
rect 15148 6414 15150 6466
rect 15202 6414 15204 6466
rect 14812 6038 14868 6076
rect 13468 5068 13636 5124
rect 13804 5906 13860 5918
rect 13804 5854 13806 5906
rect 13858 5854 13860 5906
rect 12796 5012 12852 5022
rect 12796 4918 12852 4956
rect 12684 4900 12740 4910
rect 12124 4452 12180 4462
rect 12124 3892 12180 4396
rect 12684 4338 12740 4844
rect 13468 4788 13524 5068
rect 13692 5012 13748 5022
rect 13804 5012 13860 5854
rect 14028 5906 14084 5918
rect 14028 5854 14030 5906
rect 14082 5854 14084 5906
rect 14028 5796 14084 5854
rect 14028 5730 14084 5740
rect 13692 5010 13860 5012
rect 13692 4958 13694 5010
rect 13746 4958 13860 5010
rect 13692 4956 13860 4958
rect 14700 5572 14756 5582
rect 13580 4900 13636 4910
rect 13580 4806 13636 4844
rect 12908 4452 12964 4462
rect 12908 4358 12964 4396
rect 13468 4452 13524 4732
rect 13468 4386 13524 4396
rect 12684 4286 12686 4338
rect 12738 4286 12740 4338
rect 12684 4274 12740 4286
rect 13244 4338 13300 4350
rect 13244 4286 13246 4338
rect 13298 4286 13300 4338
rect 12236 4116 12292 4126
rect 13244 4116 13300 4286
rect 13692 4226 13748 4956
rect 14028 4452 14084 4462
rect 13916 4396 14028 4452
rect 13692 4174 13694 4226
rect 13746 4174 13748 4226
rect 13692 4162 13748 4174
rect 13804 4338 13860 4350
rect 13804 4286 13806 4338
rect 13858 4286 13860 4338
rect 13804 4228 13860 4286
rect 12236 4114 13300 4116
rect 12236 4062 12238 4114
rect 12290 4062 13300 4114
rect 12236 4060 13300 4062
rect 12236 4050 12292 4060
rect 13468 4004 13524 4014
rect 13804 4004 13860 4172
rect 13524 3948 13860 4004
rect 12124 3836 12292 3892
rect 12012 3556 12068 3612
rect 12124 3556 12180 3566
rect 12012 3554 12180 3556
rect 12012 3502 12126 3554
rect 12178 3502 12180 3554
rect 12012 3500 12180 3502
rect 12124 3490 12180 3500
rect 12236 3556 12292 3836
rect 12236 3490 12292 3500
rect 12572 3780 12628 3790
rect 11676 2706 11732 2716
rect 11116 2482 11172 2492
rect 11116 2324 11172 2334
rect 11004 2268 11116 2324
rect 11116 2258 11172 2268
rect 7644 2156 8148 2212
rect 7644 800 7700 2156
rect 12572 800 12628 3724
rect 13468 3666 13524 3948
rect 13468 3614 13470 3666
rect 13522 3614 13524 3666
rect 13468 3602 13524 3614
rect 13692 3556 13748 3566
rect 13916 3556 13972 4396
rect 14028 4358 14084 4396
rect 14700 4452 14756 5516
rect 15036 5236 15092 5246
rect 15148 5236 15204 6414
rect 15518 6300 15782 6310
rect 15574 6244 15622 6300
rect 15678 6244 15726 6300
rect 15518 6234 15782 6244
rect 15820 6132 15876 6142
rect 15820 5906 15876 6076
rect 15820 5854 15822 5906
rect 15874 5854 15876 5906
rect 15484 5236 15540 5246
rect 15148 5234 15540 5236
rect 15148 5182 15486 5234
rect 15538 5182 15540 5234
rect 15148 5180 15540 5182
rect 15036 5124 15092 5180
rect 15484 5170 15540 5180
rect 15596 5236 15652 5246
rect 15036 5068 15204 5124
rect 15148 5010 15204 5068
rect 15148 4958 15150 5010
rect 15202 4958 15204 5010
rect 15148 4900 15204 4958
rect 15596 4900 15652 5180
rect 15820 5124 15876 5854
rect 15932 5684 15988 7310
rect 16044 6692 16100 8876
rect 16268 8932 16324 8942
rect 16268 8838 16324 8876
rect 16492 8258 16548 8270
rect 16492 8206 16494 8258
rect 16546 8206 16548 8258
rect 16492 7700 16548 8206
rect 16492 7634 16548 7644
rect 16380 7474 16436 7486
rect 16380 7422 16382 7474
rect 16434 7422 16436 7474
rect 16268 6692 16324 6702
rect 16044 6690 16324 6692
rect 16044 6638 16270 6690
rect 16322 6638 16324 6690
rect 16044 6636 16324 6638
rect 16268 6626 16324 6636
rect 16380 6692 16436 7422
rect 16436 6636 16548 6692
rect 16380 6626 16436 6636
rect 16156 5906 16212 5918
rect 16156 5854 16158 5906
rect 16210 5854 16212 5906
rect 16156 5796 16212 5854
rect 16156 5730 16212 5740
rect 15932 5618 15988 5628
rect 15820 5058 15876 5068
rect 16492 5010 16548 6636
rect 16492 4958 16494 5010
rect 16546 4958 16548 5010
rect 16492 4946 16548 4958
rect 15148 4834 15204 4844
rect 15260 4844 15652 4900
rect 15036 4452 15092 4462
rect 14700 4450 14868 4452
rect 14700 4398 14702 4450
rect 14754 4398 14868 4450
rect 14700 4396 14868 4398
rect 14700 4386 14756 4396
rect 13692 3554 13972 3556
rect 13692 3502 13694 3554
rect 13746 3502 13972 3554
rect 13692 3500 13972 3502
rect 14700 3556 14756 3566
rect 13692 3490 13748 3500
rect 14700 3462 14756 3500
rect 14812 3444 14868 4396
rect 15036 4358 15092 4396
rect 15260 4340 15316 4844
rect 15518 4732 15782 4742
rect 15574 4676 15622 4732
rect 15678 4676 15726 4732
rect 15518 4666 15782 4676
rect 15932 4676 15988 4686
rect 15932 4562 15988 4620
rect 15932 4510 15934 4562
rect 15986 4510 15988 4562
rect 15932 4498 15988 4510
rect 16044 4452 16100 4462
rect 15372 4340 15428 4350
rect 15260 4338 15428 4340
rect 15260 4286 15374 4338
rect 15426 4286 15428 4338
rect 15260 4284 15428 4286
rect 15372 4274 15428 4284
rect 15820 4004 15876 4014
rect 15820 3666 15876 3948
rect 16044 3778 16100 4396
rect 16268 4228 16324 4238
rect 16324 4172 16548 4228
rect 16268 4134 16324 4172
rect 16044 3726 16046 3778
rect 16098 3726 16100 3778
rect 16044 3714 16100 3726
rect 16380 3780 16436 3790
rect 16380 3686 16436 3724
rect 15820 3614 15822 3666
rect 15874 3614 15876 3666
rect 15820 3602 15876 3614
rect 14812 3378 14868 3388
rect 15260 3442 15316 3454
rect 15260 3390 15262 3442
rect 15314 3390 15316 3442
rect 15260 2436 15316 3390
rect 15518 3164 15782 3174
rect 15574 3108 15622 3164
rect 15678 3108 15726 3164
rect 15518 3098 15782 3108
rect 16492 2884 16548 4172
rect 16492 2818 16548 2828
rect 15260 2370 15316 2380
rect 16604 2212 16660 9996
rect 16828 9828 16884 9838
rect 16940 9828 16996 11340
rect 16828 9826 16996 9828
rect 16828 9774 16830 9826
rect 16882 9774 16996 9826
rect 16828 9772 16996 9774
rect 17164 11506 17220 11518
rect 17164 11454 17166 11506
rect 17218 11454 17220 11506
rect 16828 9762 16884 9772
rect 17164 9492 17220 11454
rect 17164 9426 17220 9436
rect 17388 10276 17444 10286
rect 16828 9156 16884 9166
rect 16828 9062 16884 9100
rect 16828 8372 16884 8382
rect 16716 7362 16772 7374
rect 16716 7310 16718 7362
rect 16770 7310 16772 7362
rect 16716 6356 16772 7310
rect 16828 6804 16884 8316
rect 17164 8260 17220 8270
rect 17388 8260 17444 10220
rect 17500 9938 17556 12348
rect 17612 11954 17668 12684
rect 17836 12292 17892 12302
rect 17836 12178 17892 12236
rect 18060 12292 18116 13582
rect 18060 12226 18116 12236
rect 18172 13524 18228 13694
rect 18172 12290 18228 13468
rect 18620 13636 18676 13646
rect 18732 13636 18788 18172
rect 19292 17780 19348 17790
rect 19292 17666 19348 17724
rect 19628 17780 19684 17790
rect 19292 17614 19294 17666
rect 19346 17614 19348 17666
rect 19292 17602 19348 17614
rect 19516 17666 19572 17678
rect 19516 17614 19518 17666
rect 19570 17614 19572 17666
rect 18956 15876 19012 15886
rect 18956 15782 19012 15820
rect 19516 15876 19572 17614
rect 19516 15810 19572 15820
rect 19628 16210 19684 17724
rect 19740 16548 19796 18510
rect 19740 16482 19796 16492
rect 19628 16158 19630 16210
rect 19682 16158 19684 16210
rect 19628 15540 19684 16158
rect 19628 15474 19684 15484
rect 19068 15202 19124 15214
rect 19068 15150 19070 15202
rect 19122 15150 19124 15202
rect 19068 13972 19124 15150
rect 19068 13916 19348 13972
rect 18620 13634 18788 13636
rect 18620 13582 18622 13634
rect 18674 13582 18788 13634
rect 18620 13580 18788 13582
rect 18956 13748 19012 13758
rect 18956 13636 19012 13692
rect 19068 13636 19124 13646
rect 18956 13634 19124 13636
rect 18956 13582 19070 13634
rect 19122 13582 19124 13634
rect 18956 13580 19124 13582
rect 18620 13524 18676 13580
rect 18620 13458 18676 13468
rect 18172 12238 18174 12290
rect 18226 12238 18228 12290
rect 18172 12226 18228 12238
rect 17836 12126 17838 12178
rect 17890 12126 17892 12178
rect 17836 12114 17892 12126
rect 18844 12068 18900 12078
rect 18844 11974 18900 12012
rect 17612 11902 17614 11954
rect 17666 11902 17668 11954
rect 17612 11890 17668 11902
rect 18172 11956 18228 11966
rect 17948 11508 18004 11518
rect 17836 11396 17892 11406
rect 17836 11302 17892 11340
rect 17948 11282 18004 11452
rect 18172 11394 18228 11900
rect 18620 11844 18676 11854
rect 18620 11618 18676 11788
rect 18956 11844 19012 13580
rect 19068 13570 19124 13580
rect 19180 13522 19236 13534
rect 19180 13470 19182 13522
rect 19234 13470 19236 13522
rect 18956 11778 19012 11788
rect 19068 12178 19124 12190
rect 19068 12126 19070 12178
rect 19122 12126 19124 12178
rect 19068 11732 19124 12126
rect 19068 11666 19124 11676
rect 18620 11566 18622 11618
rect 18674 11566 18676 11618
rect 18620 11554 18676 11566
rect 19068 11508 19124 11518
rect 19180 11508 19236 13470
rect 19068 11506 19236 11508
rect 19068 11454 19070 11506
rect 19122 11454 19236 11506
rect 19068 11452 19236 11454
rect 19292 13074 19348 13916
rect 19292 13022 19294 13074
rect 19346 13022 19348 13074
rect 19068 11442 19124 11452
rect 18172 11342 18174 11394
rect 18226 11342 18228 11394
rect 18172 11330 18228 11342
rect 18732 11394 18788 11406
rect 18732 11342 18734 11394
rect 18786 11342 18788 11394
rect 17948 11230 17950 11282
rect 18002 11230 18004 11282
rect 17948 11218 18004 11230
rect 18284 11172 18340 11182
rect 17500 9886 17502 9938
rect 17554 9886 17556 9938
rect 17500 9874 17556 9886
rect 17836 10498 17892 10510
rect 17836 10446 17838 10498
rect 17890 10446 17892 10498
rect 17836 10276 17892 10446
rect 17500 9042 17556 9054
rect 17500 8990 17502 9042
rect 17554 8990 17556 9042
rect 17500 8484 17556 8990
rect 17836 8932 17892 10220
rect 18172 10498 18228 10510
rect 18172 10446 18174 10498
rect 18226 10446 18228 10498
rect 18172 10164 18228 10446
rect 18172 10098 18228 10108
rect 18060 9156 18116 9166
rect 18116 9100 18228 9156
rect 18060 9090 18116 9100
rect 18172 9042 18228 9100
rect 18172 8990 18174 9042
rect 18226 8990 18228 9042
rect 18172 8978 18228 8990
rect 17836 8866 17892 8876
rect 17500 8418 17556 8428
rect 18172 8820 18228 8830
rect 17724 8372 17780 8382
rect 17500 8260 17556 8270
rect 17388 8204 17500 8260
rect 17164 8166 17220 8204
rect 17500 7698 17556 8204
rect 17724 8258 17780 8316
rect 17724 8206 17726 8258
rect 17778 8206 17780 8258
rect 17724 8194 17780 8206
rect 17836 8146 17892 8158
rect 17836 8094 17838 8146
rect 17890 8094 17892 8146
rect 17836 7812 17892 8094
rect 17836 7746 17892 7756
rect 17500 7646 17502 7698
rect 17554 7646 17556 7698
rect 17500 6916 17556 7646
rect 17500 6850 17556 6860
rect 18060 7474 18116 7486
rect 18060 7422 18062 7474
rect 18114 7422 18116 7474
rect 16828 6690 16884 6748
rect 16828 6638 16830 6690
rect 16882 6638 16884 6690
rect 16828 6626 16884 6638
rect 17836 6692 17892 6702
rect 17500 6580 17556 6590
rect 17500 6486 17556 6524
rect 17836 6578 17892 6636
rect 17836 6526 17838 6578
rect 17890 6526 17892 6578
rect 17836 6514 17892 6526
rect 16716 6290 16772 6300
rect 17052 6132 17108 6142
rect 16716 5908 16772 5918
rect 16716 5794 16772 5852
rect 16716 5742 16718 5794
rect 16770 5742 16772 5794
rect 16716 5122 16772 5742
rect 17052 5234 17108 6076
rect 17052 5182 17054 5234
rect 17106 5182 17108 5234
rect 17052 5170 17108 5182
rect 17836 5906 17892 5918
rect 17836 5854 17838 5906
rect 17890 5854 17892 5906
rect 16716 5070 16718 5122
rect 16770 5070 16772 5122
rect 16716 5058 16772 5070
rect 17388 5124 17444 5134
rect 17388 5030 17444 5068
rect 16828 5012 16884 5022
rect 16828 4564 16884 4956
rect 17724 4788 17780 4798
rect 16828 4508 16996 4564
rect 16716 4338 16772 4350
rect 16716 4286 16718 4338
rect 16770 4286 16772 4338
rect 16716 4228 16772 4286
rect 16716 4162 16772 4172
rect 16940 3666 16996 4508
rect 17724 4562 17780 4732
rect 17724 4510 17726 4562
rect 17778 4510 17780 4562
rect 17724 4498 17780 4510
rect 17500 4340 17556 4350
rect 17500 4004 17556 4284
rect 17500 3938 17556 3948
rect 16940 3614 16942 3666
rect 16994 3614 16996 3666
rect 16940 3602 16996 3614
rect 16604 2146 16660 2156
rect 17500 3444 17556 3454
rect 17500 800 17556 3388
rect 17836 3332 17892 5854
rect 18060 5348 18116 7422
rect 18060 5282 18116 5292
rect 18172 4564 18228 8764
rect 18284 7140 18340 11116
rect 18732 11172 18788 11342
rect 18732 11106 18788 11116
rect 19292 11172 19348 13022
rect 19740 13634 19796 13646
rect 19740 13582 19742 13634
rect 19794 13582 19796 13634
rect 19740 12628 19796 13582
rect 19964 13522 20020 20972
rect 20076 20802 20132 22092
rect 20188 21924 20244 22988
rect 20300 22978 20356 22988
rect 20412 22372 20468 26852
rect 20524 26852 20580 26862
rect 20636 26852 20804 26908
rect 21532 26852 21588 26862
rect 21644 26852 21812 26908
rect 20524 26402 20580 26796
rect 20748 26628 20804 26852
rect 20748 26562 20804 26572
rect 21196 26850 21588 26852
rect 21196 26798 21534 26850
rect 21586 26798 21588 26850
rect 21196 26796 21588 26798
rect 20524 26350 20526 26402
rect 20578 26350 20580 26402
rect 20524 25396 20580 26350
rect 20636 26404 20692 26414
rect 21196 26404 21252 26796
rect 21532 26786 21588 26796
rect 20636 26402 21252 26404
rect 20636 26350 20638 26402
rect 20690 26350 21252 26402
rect 20636 26348 21252 26350
rect 20636 26338 20692 26348
rect 20524 25330 20580 25340
rect 21084 23940 21140 23950
rect 20636 23380 20692 23390
rect 20636 23378 21028 23380
rect 20636 23326 20638 23378
rect 20690 23326 21028 23378
rect 20636 23324 21028 23326
rect 20636 23314 20692 23324
rect 20412 22306 20468 22316
rect 20860 23154 20916 23166
rect 20860 23102 20862 23154
rect 20914 23102 20916 23154
rect 20188 21858 20244 21868
rect 20300 22146 20356 22158
rect 20300 22094 20302 22146
rect 20354 22094 20356 22146
rect 20300 21700 20356 22094
rect 20860 21700 20916 23102
rect 20300 21644 20916 21700
rect 20300 21476 20356 21486
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20738 20132 20750
rect 20188 21474 20356 21476
rect 20188 21422 20302 21474
rect 20354 21422 20356 21474
rect 20188 21420 20356 21422
rect 20188 20578 20244 21420
rect 20300 21410 20356 21420
rect 20300 21140 20356 21150
rect 20300 21026 20356 21084
rect 20300 20974 20302 21026
rect 20354 20974 20356 21026
rect 20300 20962 20356 20974
rect 20524 20580 20580 21644
rect 20972 20916 21028 23324
rect 21084 22260 21140 23884
rect 21196 22596 21252 26348
rect 21308 26290 21364 26302
rect 21308 26238 21310 26290
rect 21362 26238 21364 26290
rect 21308 25508 21364 26238
rect 21532 26290 21588 26302
rect 21532 26238 21534 26290
rect 21586 26238 21588 26290
rect 21420 26178 21476 26190
rect 21420 26126 21422 26178
rect 21474 26126 21476 26178
rect 21420 25508 21476 26126
rect 21532 26180 21588 26238
rect 21532 26114 21588 26124
rect 21756 25956 21812 26852
rect 21868 26628 21924 27020
rect 21980 27074 22148 27076
rect 21980 27022 21982 27074
rect 22034 27022 22148 27074
rect 21980 27020 22148 27022
rect 21980 27010 22036 27020
rect 21868 26562 21924 26572
rect 21980 26290 22036 26302
rect 21980 26238 21982 26290
rect 22034 26238 22036 26290
rect 21756 25900 21924 25956
rect 21532 25844 21588 25854
rect 21532 25620 21588 25788
rect 21532 25564 21812 25620
rect 21420 25452 21588 25508
rect 21308 25442 21364 25452
rect 21420 25282 21476 25294
rect 21420 25230 21422 25282
rect 21474 25230 21476 25282
rect 21420 24834 21476 25230
rect 21420 24782 21422 24834
rect 21474 24782 21476 24834
rect 21420 24770 21476 24782
rect 21532 24724 21588 25452
rect 21756 25506 21812 25564
rect 21756 25454 21758 25506
rect 21810 25454 21812 25506
rect 21756 25442 21812 25454
rect 21644 25396 21700 25406
rect 21644 25302 21700 25340
rect 21868 25284 21924 25900
rect 21756 25228 21924 25284
rect 21644 24724 21700 24734
rect 21532 24722 21700 24724
rect 21532 24670 21646 24722
rect 21698 24670 21700 24722
rect 21532 24668 21700 24670
rect 21644 24658 21700 24668
rect 21420 24052 21476 24062
rect 21420 23958 21476 23996
rect 21420 23828 21476 23838
rect 21196 22530 21252 22540
rect 21308 23716 21364 23726
rect 21084 22194 21140 22204
rect 20972 20850 21028 20860
rect 20188 20526 20190 20578
rect 20242 20526 20244 20578
rect 20188 20514 20244 20526
rect 20300 20524 20580 20580
rect 20636 20802 20692 20814
rect 20636 20750 20638 20802
rect 20690 20750 20692 20802
rect 20188 19908 20244 19918
rect 20188 19814 20244 19852
rect 20188 19572 20244 19582
rect 20076 19236 20132 19246
rect 20076 15876 20132 19180
rect 20188 17780 20244 19516
rect 20188 17686 20244 17724
rect 20300 17220 20356 20524
rect 20636 19908 20692 20750
rect 21308 20692 21364 23660
rect 21420 21028 21476 23772
rect 21756 23826 21812 25228
rect 21980 24948 22036 26238
rect 22092 25620 22148 27020
rect 22204 27188 22260 27580
rect 22316 27524 22372 27692
rect 22316 27458 22372 27468
rect 22204 27074 22260 27132
rect 22204 27022 22206 27074
rect 22258 27022 22260 27074
rect 22204 27010 22260 27022
rect 22428 26908 22484 30716
rect 22672 30604 22936 30614
rect 22728 30548 22776 30604
rect 22832 30548 22880 30604
rect 22672 30538 22936 30548
rect 23100 29988 23156 30940
rect 23996 30930 24052 30940
rect 23324 30772 23380 30782
rect 23324 30098 23380 30716
rect 23324 30046 23326 30098
rect 23378 30046 23380 30098
rect 23324 30034 23380 30046
rect 23548 30660 23604 30670
rect 23548 30212 23604 30604
rect 23996 30436 24052 30446
rect 24108 30436 24164 31502
rect 23996 30434 24164 30436
rect 23996 30382 23998 30434
rect 24050 30382 24164 30434
rect 23996 30380 24164 30382
rect 24332 31554 24388 31566
rect 24332 31502 24334 31554
rect 24386 31502 24388 31554
rect 24332 30436 24388 31502
rect 24444 31554 24500 31566
rect 24444 31502 24446 31554
rect 24498 31502 24500 31554
rect 24444 30772 24500 31502
rect 24444 30706 24500 30716
rect 24556 31554 24612 31566
rect 24556 31502 24558 31554
rect 24610 31502 24612 31554
rect 24556 30660 24612 31502
rect 24556 30594 24612 30604
rect 24332 30380 24612 30436
rect 23996 30370 24052 30380
rect 23212 29988 23268 29998
rect 23100 29986 23268 29988
rect 23100 29934 23214 29986
rect 23266 29934 23268 29986
rect 23100 29932 23268 29934
rect 23212 29922 23268 29932
rect 23548 29428 23604 30156
rect 23884 30100 23940 30110
rect 23660 30098 23940 30100
rect 23660 30046 23886 30098
rect 23938 30046 23940 30098
rect 23660 30044 23940 30046
rect 23660 29538 23716 30044
rect 23884 30034 23940 30044
rect 23996 29988 24052 29998
rect 23996 29894 24052 29932
rect 23660 29486 23662 29538
rect 23714 29486 23716 29538
rect 23660 29474 23716 29486
rect 24332 29652 24388 30380
rect 24556 30322 24612 30380
rect 24556 30270 24558 30322
rect 24610 30270 24612 30322
rect 24556 30258 24612 30270
rect 24780 30098 24836 30110
rect 24780 30046 24782 30098
rect 24834 30046 24836 30098
rect 24780 29988 24836 30046
rect 23548 29362 23604 29372
rect 23772 29428 23828 29438
rect 23772 29334 23828 29372
rect 24332 29426 24388 29596
rect 24332 29374 24334 29426
rect 24386 29374 24388 29426
rect 24332 29362 24388 29374
rect 24668 29932 24780 29988
rect 24220 29316 24276 29326
rect 23324 29092 23380 29102
rect 22672 29036 22936 29046
rect 22728 28980 22776 29036
rect 22832 28980 22880 29036
rect 22672 28970 22936 28980
rect 22988 28756 23044 28766
rect 22540 28644 22596 28654
rect 22540 28082 22596 28588
rect 22988 28642 23044 28700
rect 22988 28590 22990 28642
rect 23042 28590 23044 28642
rect 22988 28578 23044 28590
rect 23324 28644 23380 29036
rect 23436 28980 23492 28990
rect 23436 28754 23492 28924
rect 23436 28702 23438 28754
rect 23490 28702 23492 28754
rect 23436 28690 23492 28702
rect 23324 28550 23380 28588
rect 23996 28644 24052 28654
rect 23996 28550 24052 28588
rect 24220 28532 24276 29260
rect 24668 29092 24724 29932
rect 24780 29922 24836 29932
rect 24444 29036 24724 29092
rect 24444 28754 24500 29036
rect 24444 28702 24446 28754
rect 24498 28702 24500 28754
rect 24444 28690 24500 28702
rect 24892 28756 24948 28766
rect 24892 28662 24948 28700
rect 24332 28532 24388 28542
rect 24220 28530 24388 28532
rect 24220 28478 24334 28530
rect 24386 28478 24388 28530
rect 24220 28476 24388 28478
rect 22540 28030 22542 28082
rect 22594 28030 22596 28082
rect 22540 28018 22596 28030
rect 23324 28196 23380 28206
rect 22876 27748 22932 27758
rect 22932 27692 23268 27748
rect 22876 27654 22932 27692
rect 22672 27468 22936 27478
rect 22728 27412 22776 27468
rect 22832 27412 22880 27468
rect 22672 27402 22936 27412
rect 22876 27300 22932 27310
rect 22540 27076 22596 27114
rect 22540 27010 22596 27020
rect 22652 26964 22708 27002
rect 22316 26852 22372 26862
rect 22428 26852 22596 26908
rect 22316 26758 22372 26796
rect 22316 26628 22372 26638
rect 22316 26180 22372 26572
rect 22316 26178 22484 26180
rect 22316 26126 22318 26178
rect 22370 26126 22484 26178
rect 22316 26124 22484 26126
rect 22316 26114 22372 26124
rect 22428 25844 22484 26124
rect 22092 25564 22372 25620
rect 22316 25060 22372 25564
rect 22428 25396 22484 25788
rect 22428 25330 22484 25340
rect 22316 24994 22372 25004
rect 21980 24882 22036 24892
rect 21756 23774 21758 23826
rect 21810 23774 21812 23826
rect 21532 22372 21588 22382
rect 21532 22278 21588 22316
rect 21644 22146 21700 22158
rect 21644 22094 21646 22146
rect 21698 22094 21700 22146
rect 21644 22036 21700 22094
rect 21644 21970 21700 21980
rect 21644 21812 21700 21822
rect 21420 20972 21588 21028
rect 21308 20626 21364 20636
rect 21420 20804 21476 20814
rect 20636 19842 20692 19852
rect 20972 19906 21028 19918
rect 20972 19854 20974 19906
rect 21026 19854 21028 19906
rect 20972 19236 21028 19854
rect 20972 19170 21028 19180
rect 20412 19010 20468 19022
rect 20412 18958 20414 19010
rect 20466 18958 20468 19010
rect 20412 18450 20468 18958
rect 21196 18562 21252 18574
rect 21196 18510 21198 18562
rect 21250 18510 21252 18562
rect 20412 18398 20414 18450
rect 20466 18398 20468 18450
rect 20412 18386 20468 18398
rect 20636 18452 20692 18462
rect 21084 18452 21140 18462
rect 20524 17668 20580 17678
rect 20524 17574 20580 17612
rect 20076 15782 20132 15820
rect 20188 17164 20356 17220
rect 20412 17556 20468 17566
rect 20188 14980 20244 17164
rect 20300 16772 20356 16782
rect 20300 16678 20356 16716
rect 20188 14196 20244 14924
rect 20188 14130 20244 14140
rect 20300 16548 20356 16558
rect 19964 13470 19966 13522
rect 20018 13470 20020 13522
rect 19964 13458 20020 13470
rect 20188 13634 20244 13646
rect 20188 13582 20190 13634
rect 20242 13582 20244 13634
rect 19740 12404 19796 12572
rect 19740 12338 19796 12348
rect 19964 12850 20020 12862
rect 19964 12798 19966 12850
rect 20018 12798 20020 12850
rect 19852 12292 19908 12302
rect 19852 12198 19908 12236
rect 19964 11956 20020 12798
rect 19964 11890 20020 11900
rect 20076 12738 20132 12750
rect 20076 12686 20078 12738
rect 20130 12686 20132 12738
rect 20076 11844 20132 12686
rect 20076 11778 20132 11788
rect 20188 12180 20244 13582
rect 20300 12962 20356 16492
rect 20300 12910 20302 12962
rect 20354 12910 20356 12962
rect 20300 12898 20356 12910
rect 20412 15538 20468 17500
rect 20636 17554 20692 18396
rect 20860 18450 21140 18452
rect 20860 18398 21086 18450
rect 21138 18398 21140 18450
rect 20860 18396 21140 18398
rect 20860 17666 20916 18396
rect 21084 18386 21140 18396
rect 20860 17614 20862 17666
rect 20914 17614 20916 17666
rect 20860 17602 20916 17614
rect 20636 17502 20638 17554
rect 20690 17502 20692 17554
rect 20636 17490 20692 17502
rect 20860 17108 20916 17118
rect 20748 17052 20860 17108
rect 20636 16882 20692 16894
rect 20636 16830 20638 16882
rect 20690 16830 20692 16882
rect 20524 16100 20580 16110
rect 20636 16100 20692 16830
rect 20524 16098 20692 16100
rect 20524 16046 20526 16098
rect 20578 16046 20692 16098
rect 20524 16044 20692 16046
rect 20524 16034 20580 16044
rect 20412 15486 20414 15538
rect 20466 15486 20468 15538
rect 20188 11620 20244 12124
rect 20300 11956 20356 11966
rect 20300 11732 20356 11900
rect 20300 11666 20356 11676
rect 20188 11554 20244 11564
rect 19740 11508 19796 11518
rect 19740 11394 19796 11452
rect 19740 11342 19742 11394
rect 19794 11342 19796 11394
rect 19740 11330 19796 11342
rect 19964 11396 20020 11406
rect 19964 11302 20020 11340
rect 19292 11106 19348 11116
rect 19740 10724 19796 10734
rect 19292 10612 19348 10622
rect 19292 10518 19348 10556
rect 19740 10610 19796 10668
rect 19740 10558 19742 10610
rect 19794 10558 19796 10610
rect 19180 10500 19236 10510
rect 19180 10406 19236 10444
rect 19628 10498 19684 10510
rect 19628 10446 19630 10498
rect 19682 10446 19684 10498
rect 18396 10386 18452 10398
rect 18396 10334 18398 10386
rect 18450 10334 18452 10386
rect 18396 8372 18452 10334
rect 18732 10386 18788 10398
rect 18732 10334 18734 10386
rect 18786 10334 18788 10386
rect 18620 8708 18676 8718
rect 18396 7362 18452 8316
rect 18396 7310 18398 7362
rect 18450 7310 18452 7362
rect 18396 7298 18452 7310
rect 18508 8370 18564 8382
rect 18508 8318 18510 8370
rect 18562 8318 18564 8370
rect 18284 7084 18452 7140
rect 18284 5796 18340 5806
rect 18284 5122 18340 5740
rect 18284 5070 18286 5122
rect 18338 5070 18340 5122
rect 18284 5058 18340 5070
rect 18284 4564 18340 4574
rect 18172 4508 18284 4564
rect 18284 4498 18340 4508
rect 18060 4340 18116 4350
rect 18060 4246 18116 4284
rect 17836 3266 17892 3276
rect 18396 2660 18452 7084
rect 18508 5236 18564 8318
rect 18508 5170 18564 5180
rect 18620 8258 18676 8652
rect 18620 8206 18622 8258
rect 18674 8206 18676 8258
rect 18620 6690 18676 8206
rect 18732 7252 18788 10334
rect 19628 10388 19684 10446
rect 19628 10322 19684 10332
rect 19628 9938 19684 9950
rect 19628 9886 19630 9938
rect 19682 9886 19684 9938
rect 19068 9380 19124 9390
rect 18956 7588 19012 7598
rect 19068 7588 19124 9324
rect 19628 9268 19684 9886
rect 19740 9604 19796 10558
rect 19740 9538 19796 9548
rect 20076 10722 20132 10734
rect 20076 10670 20078 10722
rect 20130 10670 20132 10722
rect 20076 9380 20132 10670
rect 20412 9940 20468 15486
rect 20636 15874 20692 15886
rect 20636 15822 20638 15874
rect 20690 15822 20692 15874
rect 20524 14642 20580 14654
rect 20524 14590 20526 14642
rect 20578 14590 20580 14642
rect 20524 13636 20580 14590
rect 20636 14308 20692 15822
rect 20748 15426 20804 17052
rect 20860 17014 20916 17052
rect 20972 16996 21028 17006
rect 20972 16902 21028 16940
rect 21196 16884 21252 18510
rect 21420 18450 21476 20748
rect 21532 19572 21588 20972
rect 21532 19506 21588 19516
rect 21644 19458 21700 21756
rect 21756 20130 21812 23774
rect 21980 23042 22036 23054
rect 21980 22990 21982 23042
rect 22034 22990 22036 23042
rect 21868 22146 21924 22158
rect 21868 22094 21870 22146
rect 21922 22094 21924 22146
rect 21868 20914 21924 22094
rect 21980 22036 22036 22990
rect 22092 22372 22148 22382
rect 22092 22258 22148 22316
rect 22428 22372 22484 22382
rect 22428 22278 22484 22316
rect 22092 22206 22094 22258
rect 22146 22206 22148 22258
rect 22092 22194 22148 22206
rect 22092 22036 22148 22046
rect 21980 21980 22092 22036
rect 21868 20862 21870 20914
rect 21922 20862 21924 20914
rect 21868 20850 21924 20862
rect 21980 20804 22036 20814
rect 21980 20710 22036 20748
rect 21756 20078 21758 20130
rect 21810 20078 21812 20130
rect 21756 20066 21812 20078
rect 22092 20132 22148 21980
rect 22428 21700 22484 21710
rect 22428 21474 22484 21644
rect 22428 21422 22430 21474
rect 22482 21422 22484 21474
rect 22428 21410 22484 21422
rect 22092 20066 22148 20076
rect 21644 19406 21646 19458
rect 21698 19406 21700 19458
rect 21644 19394 21700 19406
rect 22316 20018 22372 20030
rect 22316 19966 22318 20018
rect 22370 19966 22372 20018
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 21420 18386 21476 18398
rect 22204 18452 22260 18462
rect 22204 18358 22260 18396
rect 21308 18340 21364 18350
rect 21308 17668 21364 18284
rect 21980 18340 22036 18350
rect 21980 18246 22036 18284
rect 22316 17892 22372 19966
rect 22316 17826 22372 17836
rect 21308 16994 21364 17612
rect 21532 17556 21588 17566
rect 21532 17462 21588 17500
rect 22540 17108 22596 26852
rect 22652 26290 22708 26908
rect 22876 26962 22932 27244
rect 22988 27188 23044 27198
rect 22988 27074 23044 27132
rect 22988 27022 22990 27074
rect 23042 27022 23044 27074
rect 22988 27010 23044 27022
rect 22876 26910 22878 26962
rect 22930 26910 22932 26962
rect 22876 26898 22932 26910
rect 23212 26628 23268 27692
rect 23324 27412 23380 28140
rect 24220 27860 24276 28476
rect 24332 28466 24388 28476
rect 24556 28420 24612 28430
rect 24556 28326 24612 28364
rect 23324 27346 23380 27356
rect 23996 27858 24276 27860
rect 23996 27806 24222 27858
rect 24274 27806 24276 27858
rect 23996 27804 24276 27806
rect 23884 27188 23940 27198
rect 23660 27074 23716 27086
rect 23660 27022 23662 27074
rect 23714 27022 23716 27074
rect 23212 26562 23268 26572
rect 23548 26964 23604 26974
rect 23660 26908 23716 27022
rect 23548 26852 23716 26908
rect 23548 26402 23604 26852
rect 23548 26350 23550 26402
rect 23602 26350 23604 26402
rect 23548 26338 23604 26350
rect 22652 26238 22654 26290
rect 22706 26238 22708 26290
rect 22652 26226 22708 26238
rect 22876 26292 22932 26302
rect 22876 26198 22932 26236
rect 23772 26292 23828 26302
rect 23772 26198 23828 26236
rect 23212 26068 23268 26078
rect 23212 26066 23492 26068
rect 23212 26014 23214 26066
rect 23266 26014 23492 26066
rect 23212 26012 23492 26014
rect 23212 26002 23268 26012
rect 22672 25900 22936 25910
rect 22728 25844 22776 25900
rect 22832 25844 22880 25900
rect 22672 25834 22936 25844
rect 22876 25172 22932 25182
rect 23436 25172 23492 26012
rect 23884 25618 23940 27132
rect 23884 25566 23886 25618
rect 23938 25566 23940 25618
rect 23884 25554 23940 25566
rect 23436 25116 23716 25172
rect 22876 24946 22932 25116
rect 22876 24894 22878 24946
rect 22930 24894 22932 24946
rect 22876 24882 22932 24894
rect 23660 24946 23716 25116
rect 23660 24894 23662 24946
rect 23714 24894 23716 24946
rect 23660 24882 23716 24894
rect 23884 24948 23940 24958
rect 23996 24948 24052 27804
rect 24220 27794 24276 27804
rect 24332 27746 24388 27758
rect 24332 27694 24334 27746
rect 24386 27694 24388 27746
rect 24220 27074 24276 27086
rect 24220 27022 24222 27074
rect 24274 27022 24276 27074
rect 24220 26516 24276 27022
rect 24332 26964 24388 27694
rect 24668 27748 24724 27758
rect 24668 27654 24724 27692
rect 24892 27188 24948 27198
rect 25004 27188 25060 34972
rect 25228 34802 25284 34972
rect 25564 35028 25620 35038
rect 25676 35028 25732 35532
rect 26796 35588 26852 35598
rect 26796 35586 27300 35588
rect 26796 35534 26798 35586
rect 26850 35534 27300 35586
rect 26796 35532 27300 35534
rect 26796 35522 26852 35532
rect 25564 35026 25732 35028
rect 25564 34974 25566 35026
rect 25618 34974 25732 35026
rect 25564 34972 25732 34974
rect 25900 35476 25956 35486
rect 25564 34962 25620 34972
rect 25900 34914 25956 35420
rect 25900 34862 25902 34914
rect 25954 34862 25956 34914
rect 25900 34850 25956 34862
rect 26348 35028 26404 35038
rect 26348 34804 26404 34972
rect 26460 34916 26516 34926
rect 26460 34822 26516 34860
rect 25228 34750 25230 34802
rect 25282 34750 25284 34802
rect 25228 34738 25284 34750
rect 26236 34802 26404 34804
rect 26236 34750 26350 34802
rect 26402 34750 26404 34802
rect 26236 34748 26404 34750
rect 26124 34692 26180 34702
rect 26124 34598 26180 34636
rect 25228 34132 25284 34142
rect 25228 33346 25284 34076
rect 25676 34130 25732 34142
rect 25676 34078 25678 34130
rect 25730 34078 25732 34130
rect 25340 33908 25396 33918
rect 25340 33814 25396 33852
rect 25676 33908 25732 34078
rect 26012 34132 26068 34142
rect 26012 34018 26068 34076
rect 26012 33966 26014 34018
rect 26066 33966 26068 34018
rect 26012 33954 26068 33966
rect 25228 33294 25230 33346
rect 25282 33294 25284 33346
rect 25228 33282 25284 33294
rect 25116 33124 25172 33134
rect 25676 33124 25732 33852
rect 26124 33460 26180 33470
rect 26236 33460 26292 34748
rect 26348 34738 26404 34748
rect 27244 34802 27300 35532
rect 27244 34750 27246 34802
rect 27298 34750 27300 34802
rect 27244 34738 27300 34750
rect 27580 34802 27636 34814
rect 27580 34750 27582 34802
rect 27634 34750 27636 34802
rect 27580 34356 27636 34750
rect 27580 34290 27636 34300
rect 27580 34130 27636 34142
rect 27580 34078 27582 34130
rect 27634 34078 27636 34130
rect 26908 34018 26964 34030
rect 26908 33966 26910 34018
rect 26962 33966 26964 34018
rect 26908 33908 26964 33966
rect 26908 33842 26964 33852
rect 27580 33908 27636 34078
rect 27580 33842 27636 33852
rect 26124 33458 26292 33460
rect 26124 33406 26126 33458
rect 26178 33406 26292 33458
rect 26124 33404 26292 33406
rect 27356 33684 27412 33694
rect 26124 33394 26180 33404
rect 27244 33348 27300 33358
rect 27244 33254 27300 33292
rect 25116 33122 25732 33124
rect 25116 33070 25118 33122
rect 25170 33070 25678 33122
rect 25730 33070 25732 33122
rect 25116 33068 25732 33070
rect 25116 33058 25172 33068
rect 25676 32340 25732 33068
rect 26572 33124 26628 33134
rect 27356 33124 27412 33628
rect 27692 33572 27748 37212
rect 28812 37156 28868 37166
rect 28476 36482 28532 36494
rect 28476 36430 28478 36482
rect 28530 36430 28532 36482
rect 28364 36372 28420 36382
rect 27804 36258 27860 36270
rect 27804 36206 27806 36258
rect 27858 36206 27860 36258
rect 27804 35588 27860 36206
rect 27804 35522 27860 35532
rect 28140 34916 28196 34926
rect 28140 34914 28308 34916
rect 28140 34862 28142 34914
rect 28194 34862 28308 34914
rect 28140 34860 28308 34862
rect 28140 34850 28196 34860
rect 28252 34242 28308 34860
rect 28364 34802 28420 36316
rect 28476 36260 28532 36430
rect 28476 35364 28532 36204
rect 28476 35298 28532 35308
rect 28364 34750 28366 34802
rect 28418 34750 28420 34802
rect 28364 34738 28420 34750
rect 28252 34190 28254 34242
rect 28306 34190 28308 34242
rect 28252 34178 28308 34190
rect 28812 34354 28868 37100
rect 29148 36372 29204 36382
rect 29148 36278 29204 36316
rect 29820 36260 29876 39200
rect 32060 36932 32116 39200
rect 33292 37044 33348 37054
rect 33348 36988 33460 37044
rect 33292 36978 33348 36988
rect 32060 36866 32116 36876
rect 31276 36594 31332 36606
rect 31276 36542 31278 36594
rect 31330 36542 31332 36594
rect 29820 36204 30212 36260
rect 29825 36092 30089 36102
rect 29881 36036 29929 36092
rect 29985 36036 30033 36092
rect 29825 36026 30089 36036
rect 30156 35812 30212 36204
rect 30156 35756 30548 35812
rect 29596 35698 29652 35710
rect 29596 35646 29598 35698
rect 29650 35646 29652 35698
rect 28924 35588 28980 35598
rect 28924 35494 28980 35532
rect 29596 35364 29652 35646
rect 30380 35588 30436 35598
rect 29596 35298 29652 35308
rect 29708 35586 30436 35588
rect 29708 35534 30382 35586
rect 30434 35534 30436 35586
rect 29708 35532 30436 35534
rect 29372 34802 29428 34814
rect 29372 34750 29374 34802
rect 29426 34750 29428 34802
rect 29372 34580 29428 34750
rect 29708 34802 29764 35532
rect 30380 35522 30436 35532
rect 30156 35364 30212 35374
rect 30156 35026 30212 35308
rect 30492 35138 30548 35756
rect 30492 35086 30494 35138
rect 30546 35086 30548 35138
rect 30492 35074 30548 35086
rect 30156 34974 30158 35026
rect 30210 34974 30212 35026
rect 30156 34962 30212 34974
rect 31276 34914 31332 36542
rect 32620 36484 32676 36494
rect 32172 36428 32620 36484
rect 31836 36148 31892 36158
rect 31276 34862 31278 34914
rect 31330 34862 31332 34914
rect 31276 34850 31332 34862
rect 31724 34916 31780 34926
rect 29708 34750 29710 34802
rect 29762 34750 29764 34802
rect 29708 34738 29764 34750
rect 31612 34580 31668 34590
rect 29372 34514 29428 34524
rect 29825 34524 30089 34534
rect 29881 34468 29929 34524
rect 29985 34468 30033 34524
rect 29825 34458 30089 34468
rect 28812 34302 28814 34354
rect 28866 34302 28868 34354
rect 27580 33516 27748 33572
rect 27916 34018 27972 34030
rect 27916 33966 27918 34018
rect 27970 33966 27972 34018
rect 27580 33460 27636 33516
rect 27580 33394 27636 33404
rect 27916 33460 27972 33966
rect 28476 33908 28532 33918
rect 28252 33460 28308 33470
rect 27916 33458 28308 33460
rect 27916 33406 27918 33458
rect 27970 33406 28254 33458
rect 28306 33406 28308 33458
rect 27916 33404 28308 33406
rect 27916 33394 27972 33404
rect 28252 33394 28308 33404
rect 26572 33030 26628 33068
rect 27244 33068 27412 33124
rect 27692 33348 27748 33358
rect 26236 32676 26292 32686
rect 26236 32674 26404 32676
rect 26236 32622 26238 32674
rect 26290 32622 26404 32674
rect 26236 32620 26404 32622
rect 26236 32610 26292 32620
rect 26124 32564 26180 32574
rect 25676 32004 25732 32284
rect 25676 31938 25732 31948
rect 25900 32562 26180 32564
rect 25900 32510 26126 32562
rect 26178 32510 26180 32562
rect 25900 32508 26180 32510
rect 25900 31778 25956 32508
rect 26124 32498 26180 32508
rect 26236 32340 26292 32350
rect 25900 31726 25902 31778
rect 25954 31726 25956 31778
rect 25900 31714 25956 31726
rect 26124 32338 26292 32340
rect 26124 32286 26238 32338
rect 26290 32286 26292 32338
rect 26124 32284 26292 32286
rect 26124 31780 26180 32284
rect 26236 32274 26292 32284
rect 26124 31714 26180 31724
rect 26236 31778 26292 31790
rect 26236 31726 26238 31778
rect 26290 31726 26292 31778
rect 25564 31666 25620 31678
rect 25564 31614 25566 31666
rect 25618 31614 25620 31666
rect 25564 31108 25620 31614
rect 25676 31556 25732 31566
rect 25676 31462 25732 31500
rect 26012 31108 26068 31118
rect 26236 31108 26292 31726
rect 26348 31780 26404 32620
rect 27132 32564 27188 32574
rect 26348 31714 26404 31724
rect 26460 32004 26516 32014
rect 25564 31106 26292 31108
rect 25564 31054 26014 31106
rect 26066 31054 26292 31106
rect 25564 31052 26292 31054
rect 26012 31042 26068 31052
rect 26012 30212 26068 30222
rect 26012 30118 26068 30156
rect 25676 29652 25732 29662
rect 25676 29558 25732 29596
rect 25788 29314 25844 29326
rect 25788 29262 25790 29314
rect 25842 29262 25844 29314
rect 25116 29092 25172 29102
rect 25116 28866 25172 29036
rect 25116 28814 25118 28866
rect 25170 28814 25172 28866
rect 25116 28802 25172 28814
rect 25788 28756 25844 29262
rect 25788 28690 25844 28700
rect 25900 28980 25956 28990
rect 25900 28754 25956 28924
rect 25900 28702 25902 28754
rect 25954 28702 25956 28754
rect 25900 28690 25956 28702
rect 25452 28644 25508 28654
rect 25452 28418 25508 28588
rect 25452 28366 25454 28418
rect 25506 28366 25508 28418
rect 25452 28354 25508 28366
rect 25788 28420 25844 28430
rect 25788 28326 25844 28364
rect 25452 27970 25508 27982
rect 25452 27918 25454 27970
rect 25506 27918 25508 27970
rect 25228 27748 25284 27758
rect 25228 27654 25284 27692
rect 25452 27524 25508 27918
rect 25900 27860 25956 27870
rect 25788 27858 25956 27860
rect 25788 27806 25902 27858
rect 25954 27806 25956 27858
rect 25788 27804 25956 27806
rect 25564 27748 25620 27758
rect 25788 27748 25844 27804
rect 25900 27794 25956 27804
rect 25564 27746 25844 27748
rect 25564 27694 25566 27746
rect 25618 27694 25844 27746
rect 25564 27692 25844 27694
rect 26012 27748 26068 27758
rect 25564 27682 25620 27692
rect 25900 27636 25956 27646
rect 25900 27542 25956 27580
rect 25452 27458 25508 27468
rect 24948 27132 25060 27188
rect 26012 27186 26068 27692
rect 26236 27636 26292 27646
rect 26236 27542 26292 27580
rect 26012 27134 26014 27186
rect 26066 27134 26068 27186
rect 24892 27122 24948 27132
rect 26012 27122 26068 27134
rect 24332 26898 24388 26908
rect 26236 26964 26292 27002
rect 26236 26898 26292 26908
rect 26460 26908 26516 31948
rect 27132 31890 27188 32508
rect 27132 31838 27134 31890
rect 27186 31838 27188 31890
rect 27132 31826 27188 31838
rect 26572 31778 26628 31790
rect 26572 31726 26574 31778
rect 26626 31726 26628 31778
rect 26572 31556 26628 31726
rect 27244 31668 27300 33068
rect 27692 32786 27748 33292
rect 28476 33122 28532 33852
rect 28588 33460 28644 33470
rect 28588 33366 28644 33404
rect 28812 33348 28868 34302
rect 29372 34356 29428 34366
rect 29372 34262 29428 34300
rect 29932 34356 29988 34366
rect 29932 34018 29988 34300
rect 30940 34356 30996 34366
rect 30940 34262 30996 34300
rect 31500 34132 31556 34142
rect 31500 34038 31556 34076
rect 29932 33966 29934 34018
rect 29986 33966 29988 34018
rect 29708 33906 29764 33918
rect 29708 33854 29710 33906
rect 29762 33854 29764 33906
rect 29596 33460 29652 33470
rect 28812 33282 28868 33292
rect 29148 33348 29204 33358
rect 28476 33070 28478 33122
rect 28530 33070 28532 33122
rect 27692 32734 27694 32786
rect 27746 32734 27748 32786
rect 27692 32452 27748 32734
rect 27692 32386 27748 32396
rect 28028 32788 28084 32798
rect 28028 32450 28084 32732
rect 28028 32398 28030 32450
rect 28082 32398 28084 32450
rect 28028 32004 28084 32398
rect 28252 32452 28308 32462
rect 28252 32358 28308 32396
rect 28028 31948 28420 32004
rect 27916 31892 27972 31902
rect 27692 31836 27916 31892
rect 27356 31780 27412 31790
rect 27356 31686 27412 31724
rect 27692 31778 27748 31836
rect 27916 31826 27972 31836
rect 27692 31726 27694 31778
rect 27746 31726 27748 31778
rect 26572 29986 26628 31500
rect 27020 31612 27300 31668
rect 26684 31220 26740 31230
rect 26684 30994 26740 31164
rect 26684 30942 26686 30994
rect 26738 30942 26740 30994
rect 26684 30930 26740 30942
rect 26908 31108 26964 31118
rect 26908 30994 26964 31052
rect 26908 30942 26910 30994
rect 26962 30942 26964 30994
rect 26908 30930 26964 30942
rect 26572 29934 26574 29986
rect 26626 29934 26628 29986
rect 26572 29922 26628 29934
rect 26908 28532 26964 28542
rect 26908 27972 26964 28476
rect 27020 28308 27076 31612
rect 27580 31556 27636 31566
rect 27580 31462 27636 31500
rect 27692 31108 27748 31726
rect 28364 31668 28420 31948
rect 28476 31780 28532 33070
rect 28588 32564 28644 32574
rect 28924 32564 28980 32574
rect 29148 32564 29204 33292
rect 29484 33348 29540 33358
rect 29484 33254 29540 33292
rect 28588 32562 29204 32564
rect 28588 32510 28590 32562
rect 28642 32510 28926 32562
rect 28978 32510 29204 32562
rect 28588 32508 29204 32510
rect 29372 33124 29428 33134
rect 29372 32562 29428 33068
rect 29372 32510 29374 32562
rect 29426 32510 29428 32562
rect 28588 32498 28644 32508
rect 28924 32498 28980 32508
rect 29372 32498 29428 32510
rect 29148 32340 29204 32350
rect 29148 32246 29204 32284
rect 29596 32340 29652 33404
rect 29708 32788 29764 33854
rect 29932 33460 29988 33966
rect 30492 34018 30548 34030
rect 30492 33966 30494 34018
rect 30546 33966 30548 34018
rect 30156 33460 30212 33470
rect 29932 33458 30212 33460
rect 29932 33406 30158 33458
rect 30210 33406 30212 33458
rect 29932 33404 30212 33406
rect 29825 32956 30089 32966
rect 29881 32900 29929 32956
rect 29985 32900 30033 32956
rect 29825 32890 30089 32900
rect 29820 32788 29876 32798
rect 29708 32786 29876 32788
rect 29708 32734 29822 32786
rect 29874 32734 29876 32786
rect 29708 32732 29876 32734
rect 29820 32722 29876 32732
rect 29596 32274 29652 32284
rect 30156 32004 30212 33404
rect 30492 33346 30548 33966
rect 30492 33294 30494 33346
rect 30546 33294 30548 33346
rect 30492 33124 30548 33294
rect 30492 33058 30548 33068
rect 30940 33124 30996 33134
rect 30940 33030 30996 33068
rect 30604 33012 30660 33022
rect 30380 32676 30436 32686
rect 30380 32582 30436 32620
rect 30604 32674 30660 32956
rect 30604 32622 30606 32674
rect 30658 32622 30660 32674
rect 30604 32610 30660 32622
rect 30268 32564 30324 32574
rect 30268 32470 30324 32508
rect 30828 32564 30884 32574
rect 30828 32470 30884 32508
rect 31388 32452 31444 32462
rect 31388 32358 31444 32396
rect 30156 31938 30212 31948
rect 31612 31892 31668 34524
rect 31388 31836 31668 31892
rect 28476 31724 28868 31780
rect 28364 31612 28644 31668
rect 28588 31554 28644 31612
rect 28588 31502 28590 31554
rect 28642 31502 28644 31554
rect 27692 31042 27748 31052
rect 28252 31106 28308 31118
rect 28252 31054 28254 31106
rect 28306 31054 28308 31106
rect 28252 30548 28308 31054
rect 28364 30884 28420 30894
rect 28364 30790 28420 30828
rect 28252 30482 28308 30492
rect 28476 30770 28532 30782
rect 28476 30718 28478 30770
rect 28530 30718 28532 30770
rect 28476 30436 28532 30718
rect 28588 30436 28644 31502
rect 28588 30380 28756 30436
rect 28476 30370 28532 30380
rect 27692 30324 27748 30334
rect 27580 30322 27748 30324
rect 27580 30270 27694 30322
rect 27746 30270 27748 30322
rect 27580 30268 27748 30270
rect 27580 29428 27636 30268
rect 27692 30258 27748 30268
rect 27468 29316 27524 29326
rect 27132 29314 27524 29316
rect 27132 29262 27470 29314
rect 27522 29262 27524 29314
rect 27132 29260 27524 29262
rect 27132 28754 27188 29260
rect 27132 28702 27134 28754
rect 27186 28702 27188 28754
rect 27132 28690 27188 28702
rect 27132 28532 27188 28542
rect 27132 28438 27188 28476
rect 27020 28252 27188 28308
rect 27020 27972 27076 27982
rect 26908 27916 27020 27972
rect 27020 27906 27076 27916
rect 27132 26908 27188 28252
rect 24780 26852 24836 26862
rect 26460 26852 26628 26908
rect 24556 26850 24836 26852
rect 24556 26798 24782 26850
rect 24834 26798 24836 26850
rect 24556 26796 24836 26798
rect 24332 26516 24388 26526
rect 24220 26514 24388 26516
rect 24220 26462 24334 26514
rect 24386 26462 24388 26514
rect 24220 26460 24388 26462
rect 24220 26292 24276 26460
rect 24332 26450 24388 26460
rect 24220 26226 24276 26236
rect 24556 26402 24612 26796
rect 24780 26786 24836 26796
rect 24892 26628 24948 26638
rect 24556 26350 24558 26402
rect 24610 26350 24612 26402
rect 23884 24946 24052 24948
rect 23884 24894 23886 24946
rect 23938 24894 24052 24946
rect 23884 24892 24052 24894
rect 24108 26066 24164 26078
rect 24108 26014 24110 26066
rect 24162 26014 24164 26066
rect 24108 24946 24164 26014
rect 24556 25956 24612 26350
rect 24780 26572 24892 26628
rect 24668 26292 24724 26302
rect 24668 26198 24724 26236
rect 24556 25620 24612 25900
rect 24556 25554 24612 25564
rect 24108 24894 24110 24946
rect 24162 24894 24164 24946
rect 23884 24882 23940 24892
rect 24108 24882 24164 24894
rect 24332 24948 24388 24958
rect 22988 24836 23044 24846
rect 22988 24834 23156 24836
rect 22988 24782 22990 24834
rect 23042 24782 23156 24834
rect 22988 24780 23156 24782
rect 22988 24770 23044 24780
rect 22672 24332 22936 24342
rect 22728 24276 22776 24332
rect 22832 24276 22880 24332
rect 22672 24266 22936 24276
rect 23100 23716 23156 24780
rect 23772 24724 23828 24734
rect 23772 24630 23828 24668
rect 23212 24276 23268 24286
rect 23212 23940 23268 24220
rect 23212 23874 23268 23884
rect 24332 23938 24388 24892
rect 24332 23886 24334 23938
rect 24386 23886 24388 23938
rect 24332 23874 24388 23886
rect 24668 24612 24724 24622
rect 24668 23938 24724 24556
rect 24668 23886 24670 23938
rect 24722 23886 24724 23938
rect 24668 23874 24724 23886
rect 23324 23828 23380 23838
rect 23324 23826 23492 23828
rect 23324 23774 23326 23826
rect 23378 23774 23492 23826
rect 23324 23772 23492 23774
rect 23324 23762 23380 23772
rect 23212 23716 23268 23726
rect 23100 23714 23268 23716
rect 23100 23662 23214 23714
rect 23266 23662 23268 23714
rect 23100 23660 23268 23662
rect 23212 23650 23268 23660
rect 23436 23268 23492 23772
rect 24556 23716 24612 23726
rect 24556 23622 24612 23660
rect 24444 23604 24500 23614
rect 23548 23268 23604 23278
rect 23436 23266 23604 23268
rect 23436 23214 23550 23266
rect 23602 23214 23604 23266
rect 23436 23212 23604 23214
rect 23548 23202 23604 23212
rect 23100 23156 23156 23166
rect 22672 22764 22936 22774
rect 22728 22708 22776 22764
rect 22832 22708 22880 22764
rect 22672 22698 22936 22708
rect 23100 22596 23156 23100
rect 22876 22372 22932 22382
rect 22876 22278 22932 22316
rect 23100 22258 23156 22540
rect 24108 23154 24164 23166
rect 24108 23102 24110 23154
rect 24162 23102 24164 23154
rect 24108 22482 24164 23102
rect 24332 23156 24388 23166
rect 24108 22430 24110 22482
rect 24162 22430 24164 22482
rect 24108 22418 24164 22430
rect 24220 22596 24276 22606
rect 23100 22206 23102 22258
rect 23154 22206 23156 22258
rect 23100 22194 23156 22206
rect 23996 22260 24052 22270
rect 23996 22166 24052 22204
rect 24220 22148 24276 22540
rect 24220 22054 24276 22092
rect 24332 21924 24388 23100
rect 24444 23042 24500 23548
rect 24444 22990 24446 23042
rect 24498 22990 24500 23042
rect 24444 22978 24500 22990
rect 24444 22148 24500 22158
rect 24444 22054 24500 22092
rect 24332 21868 24500 21924
rect 22764 21812 22820 21822
rect 22764 21718 22820 21756
rect 22988 21812 23044 21822
rect 22988 21810 23828 21812
rect 22988 21758 22990 21810
rect 23042 21758 23828 21810
rect 22988 21756 23828 21758
rect 22988 21746 23044 21756
rect 23436 21586 23492 21598
rect 23436 21534 23438 21586
rect 23490 21534 23492 21586
rect 22876 21474 22932 21486
rect 22876 21422 22878 21474
rect 22930 21422 22932 21474
rect 22876 21364 22932 21422
rect 22876 21308 23380 21364
rect 22672 21196 22936 21206
rect 22728 21140 22776 21196
rect 22832 21140 22880 21196
rect 22672 21130 22936 21140
rect 22652 20690 22708 20702
rect 22652 20638 22654 20690
rect 22706 20638 22708 20690
rect 22652 20020 22708 20638
rect 23100 20132 23156 20142
rect 22988 20020 23044 20030
rect 22652 20018 23044 20020
rect 22652 19966 22990 20018
rect 23042 19966 23044 20018
rect 22652 19964 23044 19966
rect 22988 19954 23044 19964
rect 22672 19628 22936 19638
rect 22728 19572 22776 19628
rect 22832 19572 22880 19628
rect 22672 19562 22936 19572
rect 22764 19346 22820 19358
rect 22764 19294 22766 19346
rect 22818 19294 22820 19346
rect 22764 19236 22820 19294
rect 22764 18562 22820 19180
rect 22876 19348 22932 19358
rect 22876 19234 22932 19292
rect 22876 19182 22878 19234
rect 22930 19182 22932 19234
rect 22876 19170 22932 19182
rect 22764 18510 22766 18562
rect 22818 18510 22820 18562
rect 22764 18498 22820 18510
rect 23100 18450 23156 20076
rect 23324 20018 23380 21308
rect 23324 19966 23326 20018
rect 23378 19966 23380 20018
rect 23324 19954 23380 19966
rect 23436 19458 23492 21534
rect 23772 21474 23828 21756
rect 23772 21422 23774 21474
rect 23826 21422 23828 21474
rect 23772 20692 23828 21422
rect 23772 20626 23828 20636
rect 24332 20130 24388 20142
rect 24332 20078 24334 20130
rect 24386 20078 24388 20130
rect 24332 19908 24388 20078
rect 24332 19842 24388 19852
rect 23436 19406 23438 19458
rect 23490 19406 23492 19458
rect 23436 19394 23492 19406
rect 23996 19348 24052 19358
rect 23996 19254 24052 19292
rect 24444 19346 24500 21868
rect 24668 20132 24724 20142
rect 24668 20038 24724 20076
rect 24780 19348 24836 26572
rect 24892 26562 24948 26572
rect 25228 26628 25284 26638
rect 25228 26514 25284 26572
rect 25228 26462 25230 26514
rect 25282 26462 25284 26514
rect 25228 26450 25284 26462
rect 25564 26292 25620 26302
rect 25564 26198 25620 26236
rect 25228 25508 25284 25518
rect 25228 24834 25284 25452
rect 26460 25506 26516 25518
rect 26460 25454 26462 25506
rect 26514 25454 26516 25506
rect 25228 24782 25230 24834
rect 25282 24782 25284 24834
rect 25228 24770 25284 24782
rect 25788 25396 25844 25406
rect 25340 24722 25396 24734
rect 25340 24670 25342 24722
rect 25394 24670 25396 24722
rect 25340 24612 25396 24670
rect 25340 24546 25396 24556
rect 25676 24722 25732 24734
rect 25676 24670 25678 24722
rect 25730 24670 25732 24722
rect 25004 24500 25060 24510
rect 25004 22482 25060 24444
rect 25340 23828 25396 23838
rect 25676 23828 25732 24670
rect 25340 23826 25732 23828
rect 25340 23774 25342 23826
rect 25394 23774 25732 23826
rect 25340 23772 25732 23774
rect 25228 23716 25284 23726
rect 25228 23622 25284 23660
rect 25340 23044 25396 23772
rect 25788 23716 25844 25340
rect 26124 24612 26180 24622
rect 26124 23938 26180 24556
rect 26124 23886 26126 23938
rect 26178 23886 26180 23938
rect 26124 23874 26180 23886
rect 25340 22978 25396 22988
rect 25452 23714 26068 23716
rect 25452 23662 25790 23714
rect 25842 23662 26068 23714
rect 25452 23660 26068 23662
rect 25004 22430 25006 22482
rect 25058 22430 25060 22482
rect 25004 22418 25060 22430
rect 25228 22708 25284 22718
rect 25228 22372 25284 22652
rect 24892 22260 24948 22270
rect 24892 22166 24948 22204
rect 25116 22146 25172 22158
rect 25116 22094 25118 22146
rect 25170 22094 25172 22146
rect 25116 21924 25172 22094
rect 25116 21858 25172 21868
rect 25228 21476 25284 22316
rect 25340 22148 25396 22158
rect 25340 22054 25396 22092
rect 25228 21410 25284 21420
rect 25228 20916 25284 20926
rect 25228 20018 25284 20860
rect 25228 19966 25230 20018
rect 25282 19966 25284 20018
rect 25228 19954 25284 19966
rect 25452 19908 25508 23660
rect 25788 23650 25844 23660
rect 25900 23268 25956 23278
rect 25788 23266 25956 23268
rect 25788 23214 25902 23266
rect 25954 23214 25956 23266
rect 25788 23212 25956 23214
rect 25564 23044 25620 23054
rect 25788 23044 25844 23212
rect 25900 23202 25956 23212
rect 26012 23266 26068 23660
rect 26012 23214 26014 23266
rect 26066 23214 26068 23266
rect 26012 23202 26068 23214
rect 25564 23042 25844 23044
rect 25564 22990 25566 23042
rect 25618 22990 25844 23042
rect 25564 22988 25844 22990
rect 25564 22036 25620 22988
rect 25900 22930 25956 22942
rect 25900 22878 25902 22930
rect 25954 22878 25956 22930
rect 25788 22372 25844 22382
rect 25900 22372 25956 22878
rect 25788 22370 25956 22372
rect 25788 22318 25790 22370
rect 25842 22318 25956 22370
rect 25788 22316 25956 22318
rect 26124 22372 26180 22382
rect 26348 22372 26404 22382
rect 26124 22370 26404 22372
rect 26124 22318 26126 22370
rect 26178 22318 26350 22370
rect 26402 22318 26404 22370
rect 26124 22316 26404 22318
rect 25788 22306 25844 22316
rect 26124 22306 26180 22316
rect 26348 22306 26404 22316
rect 26012 22260 26068 22270
rect 25900 22204 26012 22260
rect 25900 22146 25956 22204
rect 26012 22194 26068 22204
rect 25900 22094 25902 22146
rect 25954 22094 25956 22146
rect 25900 22082 25956 22094
rect 25788 22036 25844 22046
rect 25564 21980 25788 22036
rect 25788 21810 25844 21980
rect 26124 22036 26180 22046
rect 25788 21758 25790 21810
rect 25842 21758 25844 21810
rect 25788 21746 25844 21758
rect 25900 21924 25956 21934
rect 25900 21810 25956 21868
rect 25900 21758 25902 21810
rect 25954 21758 25956 21810
rect 25900 21746 25956 21758
rect 26124 21810 26180 21980
rect 26124 21758 26126 21810
rect 26178 21758 26180 21810
rect 26124 21746 26180 21758
rect 26236 21586 26292 21598
rect 26236 21534 26238 21586
rect 26290 21534 26292 21586
rect 26236 21476 26292 21534
rect 26236 21410 26292 21420
rect 26348 21252 26404 21262
rect 26012 20244 26068 20254
rect 26012 20130 26068 20188
rect 26012 20078 26014 20130
rect 26066 20078 26068 20130
rect 26012 20066 26068 20078
rect 26348 20132 26404 21196
rect 26460 20916 26516 25454
rect 26572 21028 26628 26852
rect 27020 26852 27188 26908
rect 27356 27860 27412 27870
rect 27356 27524 27412 27804
rect 27356 26908 27412 27468
rect 27468 27300 27524 29260
rect 27580 28980 27636 29372
rect 27580 28914 27636 28924
rect 27916 30210 27972 30222
rect 27916 30158 27918 30210
rect 27970 30158 27972 30210
rect 27916 29316 27972 30158
rect 28588 30212 28644 30222
rect 28588 30118 28644 30156
rect 28252 29764 28308 29774
rect 28028 29708 28252 29764
rect 28308 29708 28532 29764
rect 28028 29538 28084 29708
rect 28252 29698 28308 29708
rect 28028 29486 28030 29538
rect 28082 29486 28084 29538
rect 28028 29474 28084 29486
rect 27916 28866 27972 29260
rect 27916 28814 27918 28866
rect 27970 28814 27972 28866
rect 27916 28802 27972 28814
rect 28476 28754 28532 29708
rect 28700 28868 28756 30380
rect 28812 29316 28868 31724
rect 30156 31778 30212 31790
rect 30156 31726 30158 31778
rect 30210 31726 30212 31778
rect 29148 31668 29204 31678
rect 29148 31574 29204 31612
rect 29825 31388 30089 31398
rect 29881 31332 29929 31388
rect 29985 31332 30033 31388
rect 29825 31322 30089 31332
rect 29372 31220 29428 31230
rect 29260 31164 29372 31220
rect 29148 30994 29204 31006
rect 29148 30942 29150 30994
rect 29202 30942 29204 30994
rect 28924 30882 28980 30894
rect 28924 30830 28926 30882
rect 28978 30830 28980 30882
rect 28924 30772 28980 30830
rect 28924 30706 28980 30716
rect 29148 30210 29204 30942
rect 29148 30158 29150 30210
rect 29202 30158 29204 30210
rect 29148 30146 29204 30158
rect 29260 29650 29316 31164
rect 29372 31154 29428 31164
rect 29820 30994 29876 31006
rect 29820 30942 29822 30994
rect 29874 30942 29876 30994
rect 29372 30884 29428 30894
rect 29372 30790 29428 30828
rect 29820 30884 29876 30942
rect 29820 30818 29876 30828
rect 29372 30548 29428 30558
rect 29372 30098 29428 30492
rect 29484 30436 29540 30446
rect 29484 30210 29540 30380
rect 30156 30436 30212 31726
rect 30604 30884 30660 30894
rect 30604 30790 30660 30828
rect 31388 30436 31444 31836
rect 31724 31780 31780 34860
rect 31836 34804 31892 36092
rect 32172 35364 32228 36428
rect 32620 36390 32676 36428
rect 33292 36372 33348 36382
rect 33180 36370 33348 36372
rect 33180 36318 33294 36370
rect 33346 36318 33348 36370
rect 33180 36316 33348 36318
rect 33068 35700 33124 35710
rect 32508 35698 33124 35700
rect 32508 35646 33070 35698
rect 33122 35646 33124 35698
rect 32508 35644 33124 35646
rect 32508 35586 32564 35644
rect 33068 35634 33124 35644
rect 32508 35534 32510 35586
rect 32562 35534 32564 35586
rect 32508 35522 32564 35534
rect 32172 35026 32228 35308
rect 32172 34974 32174 35026
rect 32226 34974 32228 35026
rect 32172 34962 32228 34974
rect 32956 34914 33012 34926
rect 32956 34862 32958 34914
rect 33010 34862 33012 34914
rect 31836 34738 31892 34748
rect 32732 34802 32788 34814
rect 32732 34750 32734 34802
rect 32786 34750 32788 34802
rect 32172 34132 32228 34142
rect 32172 34038 32228 34076
rect 32396 34020 32452 34030
rect 32396 33926 32452 33964
rect 32732 34020 32788 34750
rect 32732 33954 32788 33964
rect 32844 34690 32900 34702
rect 32844 34638 32846 34690
rect 32898 34638 32900 34690
rect 32844 33908 32900 34638
rect 32956 34692 33012 34862
rect 32956 34132 33012 34636
rect 33180 34354 33236 36316
rect 33292 36306 33348 36316
rect 33180 34302 33182 34354
rect 33234 34302 33236 34354
rect 33180 34290 33236 34302
rect 33292 34802 33348 34814
rect 33292 34750 33294 34802
rect 33346 34750 33348 34802
rect 32956 34066 33012 34076
rect 32844 33842 32900 33852
rect 33292 33460 33348 34750
rect 33404 33572 33460 36988
rect 33740 36932 33796 36942
rect 33740 35586 33796 36876
rect 33740 35534 33742 35586
rect 33794 35534 33796 35586
rect 33740 35522 33796 35534
rect 33964 35476 34020 35486
rect 33740 35028 33796 35038
rect 33740 34914 33796 34972
rect 33740 34862 33742 34914
rect 33794 34862 33796 34914
rect 33740 34850 33796 34862
rect 33964 34914 34020 35420
rect 34300 35252 34356 39200
rect 34524 37044 34580 37054
rect 34524 35586 34580 36988
rect 35308 36596 35364 36606
rect 35308 36036 35364 36540
rect 35420 36596 35476 36606
rect 35420 36594 35812 36596
rect 35420 36542 35422 36594
rect 35474 36542 35812 36594
rect 35420 36540 35812 36542
rect 35420 36530 35476 36540
rect 35308 35980 35588 36036
rect 35532 35922 35588 35980
rect 35532 35870 35534 35922
rect 35586 35870 35588 35922
rect 35532 35812 35588 35870
rect 35532 35746 35588 35756
rect 34524 35534 34526 35586
rect 34578 35534 34580 35586
rect 34524 35476 34580 35534
rect 34524 35410 34580 35420
rect 34300 35186 34356 35196
rect 35084 35252 35140 35262
rect 35084 35138 35140 35196
rect 35084 35086 35086 35138
rect 35138 35086 35140 35138
rect 35084 35074 35140 35086
rect 35308 35140 35364 35150
rect 33964 34862 33966 34914
rect 34018 34862 34020 34914
rect 33964 34850 34020 34862
rect 33852 34692 33908 34702
rect 33852 34598 33908 34636
rect 34188 34692 34244 34702
rect 34188 34598 34244 34636
rect 34860 34690 34916 34702
rect 34860 34638 34862 34690
rect 34914 34638 34916 34690
rect 33516 34356 33572 34366
rect 33516 34242 33572 34300
rect 33516 34190 33518 34242
rect 33570 34190 33572 34242
rect 33516 34178 33572 34190
rect 34860 34356 34916 34638
rect 34748 34130 34804 34142
rect 34748 34078 34750 34130
rect 34802 34078 34804 34130
rect 33964 34020 34020 34030
rect 33964 33926 34020 33964
rect 34076 34018 34132 34030
rect 34076 33966 34078 34018
rect 34130 33966 34132 34018
rect 33404 33516 33572 33572
rect 33292 33394 33348 33404
rect 32620 33346 32676 33358
rect 32620 33294 32622 33346
rect 32674 33294 32676 33346
rect 32172 33234 32228 33246
rect 32172 33182 32174 33234
rect 32226 33182 32228 33234
rect 31836 33012 31892 33022
rect 31836 32562 31892 32956
rect 31836 32510 31838 32562
rect 31890 32510 31892 32562
rect 31836 32498 31892 32510
rect 32172 32788 32228 33182
rect 32620 33012 32676 33294
rect 32620 32946 32676 32956
rect 33404 33346 33460 33358
rect 33404 33294 33406 33346
rect 33458 33294 33460 33346
rect 33292 32788 33348 32798
rect 32172 32786 33348 32788
rect 32172 32734 33294 32786
rect 33346 32734 33348 32786
rect 32172 32732 33348 32734
rect 32172 32004 32228 32732
rect 33292 32722 33348 32732
rect 32284 32564 32340 32574
rect 33068 32564 33124 32574
rect 32284 32562 33124 32564
rect 32284 32510 32286 32562
rect 32338 32510 33070 32562
rect 33122 32510 33124 32562
rect 32284 32508 33124 32510
rect 32284 32498 32340 32508
rect 33068 32498 33124 32508
rect 33180 32564 33236 32574
rect 33180 32470 33236 32508
rect 33292 32452 33348 32462
rect 33404 32452 33460 33294
rect 33516 32788 33572 33516
rect 33964 33460 34020 33470
rect 34076 33460 34132 33966
rect 34748 33684 34804 34078
rect 34860 34020 34916 34300
rect 35308 34242 35364 35084
rect 35756 34914 35812 36540
rect 36540 36594 36596 39200
rect 36979 36876 37243 36886
rect 37035 36820 37083 36876
rect 37139 36820 37187 36876
rect 36979 36810 37243 36820
rect 36540 36542 36542 36594
rect 36594 36542 36596 36594
rect 36540 36530 36596 36542
rect 37212 36596 37268 36606
rect 37212 36482 37268 36540
rect 37212 36430 37214 36482
rect 37266 36430 37268 36482
rect 37212 36418 37268 36430
rect 37996 36482 38052 36494
rect 37996 36430 37998 36482
rect 38050 36430 38052 36482
rect 35868 35812 35924 35822
rect 35868 35698 35924 35756
rect 35868 35646 35870 35698
rect 35922 35646 35924 35698
rect 35868 35634 35924 35646
rect 36428 35812 36484 35822
rect 36428 35698 36484 35756
rect 36428 35646 36430 35698
rect 36482 35646 36484 35698
rect 36428 35634 36484 35646
rect 37772 35810 37828 35822
rect 37772 35758 37774 35810
rect 37826 35758 37828 35810
rect 37772 35700 37828 35758
rect 37772 35634 37828 35644
rect 37436 35588 37492 35598
rect 37436 35494 37492 35532
rect 35756 34862 35758 34914
rect 35810 34862 35812 34914
rect 35756 34850 35812 34862
rect 36428 35476 36484 35486
rect 36428 34690 36484 35420
rect 37996 35476 38052 36430
rect 38556 36482 38612 36494
rect 38556 36430 38558 36482
rect 38610 36430 38612 36482
rect 38556 36372 38612 36430
rect 38556 36306 38612 36316
rect 37996 35410 38052 35420
rect 37660 35364 37716 35374
rect 36979 35308 37243 35318
rect 37035 35252 37083 35308
rect 37139 35252 37187 35308
rect 36979 35242 37243 35252
rect 36988 35028 37044 35038
rect 37212 35028 37268 35038
rect 36988 34934 37044 34972
rect 37100 34972 37212 35028
rect 37100 34804 37156 34972
rect 37212 34962 37268 34972
rect 36764 34802 37156 34804
rect 36764 34750 37102 34802
rect 37154 34750 37156 34802
rect 36764 34748 37156 34750
rect 36428 34638 36430 34690
rect 36482 34638 36484 34690
rect 35308 34190 35310 34242
rect 35362 34190 35364 34242
rect 35308 34178 35364 34190
rect 35980 34356 36036 34366
rect 35980 34130 36036 34300
rect 35980 34078 35982 34130
rect 36034 34078 36036 34130
rect 35980 34066 36036 34078
rect 36204 34020 36260 34030
rect 34860 33964 35140 34020
rect 34748 33628 34916 33684
rect 34636 33460 34692 33470
rect 33964 33458 34356 33460
rect 33964 33406 33966 33458
rect 34018 33406 34356 33458
rect 33964 33404 34356 33406
rect 33964 33394 34020 33404
rect 34300 33346 34356 33404
rect 34300 33294 34302 33346
rect 34354 33294 34356 33346
rect 34300 33282 34356 33294
rect 34524 33236 34580 33246
rect 34524 33142 34580 33180
rect 34636 33122 34692 33404
rect 34860 33460 34916 33628
rect 34860 33394 34916 33404
rect 34972 33348 35028 33358
rect 34972 33254 35028 33292
rect 34636 33070 34638 33122
rect 34690 33070 34692 33122
rect 34636 33058 34692 33070
rect 33516 32732 33684 32788
rect 33348 32396 33460 32452
rect 33516 32564 33572 32574
rect 33292 32386 33348 32396
rect 33516 32116 33572 32508
rect 33404 32060 33572 32116
rect 32396 32004 32452 32014
rect 32172 32002 32452 32004
rect 32172 31950 32398 32002
rect 32450 31950 32452 32002
rect 32172 31948 32452 31950
rect 32396 31938 32452 31948
rect 33404 32002 33460 32060
rect 33628 32004 33684 32732
rect 34412 32674 34468 32686
rect 34412 32622 34414 32674
rect 34466 32622 34468 32674
rect 34300 32564 34356 32574
rect 34412 32564 34468 32622
rect 34412 32508 34916 32564
rect 34300 32470 34356 32508
rect 33404 31950 33406 32002
rect 33458 31950 33460 32002
rect 33404 31938 33460 31950
rect 33516 31948 33684 32004
rect 34412 32338 34468 32350
rect 34412 32286 34414 32338
rect 34466 32286 34468 32338
rect 31724 31714 31780 31724
rect 31836 31890 31892 31902
rect 31836 31838 31838 31890
rect 31890 31838 31892 31890
rect 31500 31666 31556 31678
rect 31500 31614 31502 31666
rect 31554 31614 31556 31666
rect 31500 30884 31556 31614
rect 31724 31556 31780 31566
rect 31500 30818 31556 30828
rect 31612 30994 31668 31006
rect 31612 30942 31614 30994
rect 31666 30942 31668 30994
rect 31388 30380 31556 30436
rect 30044 30212 30100 30222
rect 29484 30158 29486 30210
rect 29538 30158 29540 30210
rect 29484 30146 29540 30158
rect 29596 30210 30100 30212
rect 29596 30158 30046 30210
rect 30098 30158 30100 30210
rect 29596 30156 30100 30158
rect 29372 30046 29374 30098
rect 29426 30046 29428 30098
rect 29372 30034 29428 30046
rect 29596 29764 29652 30156
rect 30044 30146 30100 30156
rect 29596 29698 29652 29708
rect 29708 29988 29764 29998
rect 29260 29598 29262 29650
rect 29314 29598 29316 29650
rect 29260 29586 29316 29598
rect 29036 29428 29092 29438
rect 29036 29334 29092 29372
rect 28812 29250 28868 29260
rect 29596 29316 29652 29326
rect 28700 28812 28980 28868
rect 28476 28702 28478 28754
rect 28530 28702 28532 28754
rect 28476 28532 28532 28702
rect 28476 28466 28532 28476
rect 28812 28084 28868 28094
rect 27692 27860 27748 27870
rect 27692 27766 27748 27804
rect 28028 27858 28084 27870
rect 28028 27806 28030 27858
rect 28082 27806 28084 27858
rect 28028 27748 28084 27806
rect 28812 27858 28868 28028
rect 28812 27806 28814 27858
rect 28866 27806 28868 27858
rect 28028 27524 28084 27692
rect 28140 27748 28196 27758
rect 28476 27748 28532 27758
rect 28140 27746 28532 27748
rect 28140 27694 28142 27746
rect 28194 27694 28478 27746
rect 28530 27694 28532 27746
rect 28140 27692 28532 27694
rect 28140 27682 28196 27692
rect 28476 27682 28532 27692
rect 28588 27748 28644 27758
rect 28588 27654 28644 27692
rect 28028 27458 28084 27468
rect 27468 27244 28196 27300
rect 27468 27074 27524 27244
rect 27468 27022 27470 27074
rect 27522 27022 27524 27074
rect 27468 27010 27524 27022
rect 27916 26964 27972 27002
rect 27356 26852 27748 26908
rect 27916 26898 27972 26908
rect 27020 24836 27076 26852
rect 27580 26178 27636 26190
rect 27580 26126 27582 26178
rect 27634 26126 27636 26178
rect 27580 25396 27636 26126
rect 27580 25330 27636 25340
rect 27132 25284 27188 25294
rect 27132 24946 27188 25228
rect 27132 24894 27134 24946
rect 27186 24894 27188 24946
rect 27132 24882 27188 24894
rect 27692 24948 27748 26852
rect 28140 25732 28196 27244
rect 28812 26908 28868 27806
rect 28476 26852 28868 26908
rect 28476 26402 28532 26852
rect 28476 26350 28478 26402
rect 28530 26350 28532 26402
rect 28476 26338 28532 26350
rect 28140 25666 28196 25676
rect 28476 26178 28532 26190
rect 28476 26126 28478 26178
rect 28530 26126 28532 26178
rect 27916 25508 27972 25518
rect 27916 25414 27972 25452
rect 27804 25396 27860 25406
rect 27804 25302 27860 25340
rect 28028 25394 28084 25406
rect 28028 25342 28030 25394
rect 28082 25342 28084 25394
rect 27692 24882 27748 24892
rect 27916 25284 27972 25294
rect 27020 24770 27076 24780
rect 27580 24836 27636 24846
rect 27580 24724 27636 24780
rect 27468 24722 27636 24724
rect 27468 24670 27582 24722
rect 27634 24670 27636 24722
rect 27468 24668 27636 24670
rect 27020 24052 27076 24062
rect 27020 23958 27076 23996
rect 26796 23938 26852 23950
rect 26796 23886 26798 23938
rect 26850 23886 26852 23938
rect 26796 23548 26852 23886
rect 27468 23604 27524 24668
rect 27580 24658 27636 24668
rect 27916 24610 27972 25228
rect 27916 24558 27918 24610
rect 27970 24558 27972 24610
rect 27916 24546 27972 24558
rect 28028 24724 28084 25342
rect 28476 24948 28532 26126
rect 28588 25732 28644 25742
rect 28588 25060 28644 25676
rect 28700 25284 28756 25294
rect 28700 25282 28868 25284
rect 28700 25230 28702 25282
rect 28754 25230 28868 25282
rect 28700 25228 28868 25230
rect 28700 25218 28756 25228
rect 28812 25172 28868 25228
rect 28588 25004 28756 25060
rect 28476 24882 28532 24892
rect 28028 24498 28084 24668
rect 28028 24446 28030 24498
rect 28082 24446 28084 24498
rect 28028 24434 28084 24446
rect 27132 23548 27524 23604
rect 27580 24052 27636 24062
rect 27580 23714 27636 23996
rect 27804 23940 27860 23950
rect 28476 23940 28532 23950
rect 27804 23938 28532 23940
rect 27804 23886 27806 23938
rect 27858 23886 28478 23938
rect 28530 23886 28532 23938
rect 27804 23884 28532 23886
rect 27804 23874 27860 23884
rect 27580 23662 27582 23714
rect 27634 23662 27636 23714
rect 26796 23492 27076 23548
rect 27020 23380 27076 23492
rect 27020 23314 27076 23324
rect 26684 23154 26740 23166
rect 26684 23102 26686 23154
rect 26738 23102 26740 23154
rect 26684 21924 26740 23102
rect 26908 23044 26964 23054
rect 26684 21858 26740 21868
rect 26796 23042 26964 23044
rect 26796 22990 26910 23042
rect 26962 22990 26964 23042
rect 26796 22988 26964 22990
rect 26796 22484 26852 22988
rect 26908 22978 26964 22988
rect 26796 21474 26852 22428
rect 26796 21422 26798 21474
rect 26850 21422 26852 21474
rect 26796 21410 26852 21422
rect 26572 20972 26740 21028
rect 26460 20914 26628 20916
rect 26460 20862 26462 20914
rect 26514 20862 26628 20914
rect 26460 20860 26628 20862
rect 26460 20850 26516 20860
rect 25676 19908 25732 19918
rect 25452 19852 25676 19908
rect 24892 19348 24948 19358
rect 24444 19294 24446 19346
rect 24498 19294 24500 19346
rect 23772 19236 23828 19246
rect 23772 19142 23828 19180
rect 23772 19012 23828 19022
rect 23100 18398 23102 18450
rect 23154 18398 23156 18450
rect 23100 18386 23156 18398
rect 23212 18564 23268 18574
rect 22672 18060 22936 18070
rect 22728 18004 22776 18060
rect 22832 18004 22880 18060
rect 22672 17994 22936 18004
rect 23100 17108 23156 17118
rect 22540 17052 22820 17108
rect 21308 16942 21310 16994
rect 21362 16942 21364 16994
rect 21308 16930 21364 16942
rect 22204 16940 22708 16996
rect 21196 16818 21252 16828
rect 21756 16882 21812 16894
rect 21756 16830 21758 16882
rect 21810 16830 21812 16882
rect 21756 16660 21812 16830
rect 21756 16594 21812 16604
rect 21868 16884 21924 16894
rect 21756 16210 21812 16222
rect 21756 16158 21758 16210
rect 21810 16158 21812 16210
rect 20860 16100 20916 16110
rect 20860 16006 20916 16044
rect 21756 16100 21812 16158
rect 21756 16034 21812 16044
rect 20748 15374 20750 15426
rect 20802 15374 20804 15426
rect 20748 15362 20804 15374
rect 21084 15876 21140 15886
rect 20636 14242 20692 14252
rect 20524 13570 20580 13580
rect 20636 13634 20692 13646
rect 20636 13582 20638 13634
rect 20690 13582 20692 13634
rect 20636 12740 20692 13582
rect 20972 13636 21028 13646
rect 20972 13542 21028 13580
rect 21084 13076 21140 15820
rect 21644 15764 21700 15774
rect 21420 15428 21476 15438
rect 21420 15314 21476 15372
rect 21420 15262 21422 15314
rect 21474 15262 21476 15314
rect 21420 15250 21476 15262
rect 21532 15202 21588 15214
rect 21532 15150 21534 15202
rect 21586 15150 21588 15202
rect 21532 15148 21588 15150
rect 21308 15092 21588 15148
rect 21308 14532 21364 15092
rect 21644 14980 21700 15708
rect 21868 15540 21924 16828
rect 22204 16882 22260 16940
rect 22204 16830 22206 16882
rect 22258 16830 22260 16882
rect 22204 16818 22260 16830
rect 22092 16660 22148 16670
rect 21980 15540 22036 15550
rect 21868 15538 22036 15540
rect 21868 15486 21982 15538
rect 22034 15486 22036 15538
rect 21868 15484 22036 15486
rect 22092 15540 22148 16604
rect 22204 15988 22260 15998
rect 22204 15894 22260 15932
rect 22204 15540 22260 15550
rect 22092 15538 22260 15540
rect 22092 15486 22206 15538
rect 22258 15486 22260 15538
rect 22092 15484 22260 15486
rect 21980 15474 22036 15484
rect 22204 15474 22260 15484
rect 22316 15426 22372 16940
rect 22652 16882 22708 16940
rect 22652 16830 22654 16882
rect 22706 16830 22708 16882
rect 22652 16818 22708 16830
rect 22764 16660 22820 17052
rect 23100 16882 23156 17052
rect 23100 16830 23102 16882
rect 23154 16830 23156 16882
rect 23100 16818 23156 16830
rect 22316 15374 22318 15426
rect 22370 15374 22372 15426
rect 22316 15362 22372 15374
rect 22428 16604 22820 16660
rect 21644 14914 21700 14924
rect 21308 14438 21364 14476
rect 21756 14644 21812 14654
rect 21756 14530 21812 14588
rect 21756 14478 21758 14530
rect 21810 14478 21812 14530
rect 21756 14466 21812 14478
rect 22204 14530 22260 14542
rect 22204 14478 22206 14530
rect 22258 14478 22260 14530
rect 21084 13010 21140 13020
rect 21196 14420 21252 14430
rect 20636 12674 20692 12684
rect 20860 12738 20916 12750
rect 20860 12686 20862 12738
rect 20914 12686 20916 12738
rect 20636 12404 20692 12414
rect 20524 11508 20580 11518
rect 20524 11414 20580 11452
rect 20524 11172 20580 11182
rect 20636 11172 20692 12348
rect 20860 12068 20916 12686
rect 20748 11620 20804 11630
rect 20748 11526 20804 11564
rect 20860 11508 20916 12012
rect 20860 11442 20916 11452
rect 20524 11170 20692 11172
rect 20524 11118 20526 11170
rect 20578 11118 20692 11170
rect 20524 11116 20692 11118
rect 20524 10164 20580 11116
rect 20524 10098 20580 10108
rect 20636 10836 20692 10846
rect 20636 10724 20692 10780
rect 21196 10724 21252 14364
rect 21644 13858 21700 13870
rect 21644 13806 21646 13858
rect 21698 13806 21700 13858
rect 21420 13746 21476 13758
rect 21420 13694 21422 13746
rect 21474 13694 21476 13746
rect 21420 13636 21476 13694
rect 21644 13748 21700 13806
rect 22204 13860 22260 14478
rect 22204 13794 22260 13804
rect 22092 13748 22148 13758
rect 21644 13746 22148 13748
rect 21644 13694 22094 13746
rect 22146 13694 22148 13746
rect 21644 13692 22148 13694
rect 21420 13570 21476 13580
rect 21868 13524 21924 13534
rect 21756 12964 21812 12974
rect 21644 12908 21756 12964
rect 21308 11396 21364 11406
rect 21308 11302 21364 11340
rect 20636 10668 21252 10724
rect 20412 9884 20580 9940
rect 20188 9604 20244 9614
rect 20188 9510 20244 9548
rect 20076 9324 20468 9380
rect 19628 9202 19684 9212
rect 20412 9266 20468 9324
rect 20412 9214 20414 9266
rect 20466 9214 20468 9266
rect 20412 9156 20468 9214
rect 20412 9090 20468 9100
rect 19740 8484 19796 8494
rect 18956 7586 19124 7588
rect 18956 7534 18958 7586
rect 19010 7534 19124 7586
rect 18956 7532 19124 7534
rect 19180 8146 19236 8158
rect 19180 8094 19182 8146
rect 19234 8094 19236 8146
rect 19180 7588 19236 8094
rect 19292 8148 19348 8158
rect 19292 7698 19348 8092
rect 19292 7646 19294 7698
rect 19346 7646 19348 7698
rect 19292 7634 19348 7646
rect 18844 7476 18900 7486
rect 18844 7382 18900 7420
rect 18732 7186 18788 7196
rect 18620 6638 18622 6690
rect 18674 6638 18676 6690
rect 18620 5124 18676 6638
rect 18620 5058 18676 5068
rect 18956 5906 19012 7532
rect 19180 7522 19236 7532
rect 18956 5854 18958 5906
rect 19010 5854 19012 5906
rect 18508 4676 18564 4686
rect 18508 4450 18564 4620
rect 18956 4564 19012 5854
rect 19068 6690 19124 6702
rect 19068 6638 19070 6690
rect 19122 6638 19124 6690
rect 19068 5124 19124 6638
rect 19180 5124 19236 5134
rect 19068 5122 19236 5124
rect 19068 5070 19182 5122
rect 19234 5070 19236 5122
rect 19068 5068 19236 5070
rect 19180 4676 19236 5068
rect 19292 5124 19348 5134
rect 19516 5124 19572 5134
rect 19348 5122 19572 5124
rect 19348 5070 19518 5122
rect 19570 5070 19572 5122
rect 19348 5068 19572 5070
rect 19292 5058 19348 5068
rect 19516 5058 19572 5068
rect 19180 4610 19236 4620
rect 18956 4508 19124 4564
rect 18508 4398 18510 4450
rect 18562 4398 18564 4450
rect 18508 4386 18564 4398
rect 19068 4340 19124 4508
rect 19404 4452 19460 4462
rect 19404 4340 19460 4396
rect 19068 4338 19460 4340
rect 19068 4286 19406 4338
rect 19458 4286 19460 4338
rect 19068 4284 19460 4286
rect 19404 4274 19460 4284
rect 19068 4116 19124 4126
rect 19068 3666 19124 4060
rect 19068 3614 19070 3666
rect 19122 3614 19124 3666
rect 19068 3602 19124 3614
rect 19740 3556 19796 8428
rect 20412 8484 20468 8494
rect 20524 8484 20580 9884
rect 20468 8428 20580 8484
rect 20636 9826 20692 10668
rect 21644 10610 21700 12908
rect 21756 12898 21812 12908
rect 21756 12738 21812 12750
rect 21756 12686 21758 12738
rect 21810 12686 21812 12738
rect 21756 11956 21812 12686
rect 21868 12628 21924 13468
rect 22092 13188 22148 13692
rect 22428 13636 22484 16604
rect 23212 16548 23268 18508
rect 23660 18450 23716 18462
rect 23660 18398 23662 18450
rect 23714 18398 23716 18450
rect 23548 17892 23604 17902
rect 23324 17108 23380 17118
rect 23324 16772 23380 17052
rect 23324 16706 23380 16716
rect 23436 16996 23492 17006
rect 23436 16770 23492 16940
rect 23436 16718 23438 16770
rect 23490 16718 23492 16770
rect 23436 16706 23492 16718
rect 22672 16492 22936 16502
rect 23212 16492 23492 16548
rect 22728 16436 22776 16492
rect 22832 16436 22880 16492
rect 22672 16426 22936 16436
rect 23324 16100 23380 16110
rect 23324 16006 23380 16044
rect 22540 15428 22596 15438
rect 22540 14756 22596 15372
rect 22764 15314 22820 15326
rect 22764 15262 22766 15314
rect 22818 15262 22820 15314
rect 22764 15204 22820 15262
rect 22764 15138 22820 15148
rect 23100 15314 23156 15326
rect 23100 15262 23102 15314
rect 23154 15262 23156 15314
rect 22672 14924 22936 14934
rect 22728 14868 22776 14924
rect 22832 14868 22880 14924
rect 22672 14858 22936 14868
rect 22540 14700 22820 14756
rect 22652 14532 22708 14542
rect 22652 14438 22708 14476
rect 22764 14418 22820 14700
rect 23100 14532 23156 15262
rect 23212 15316 23268 15326
rect 23212 15222 23268 15260
rect 23324 15314 23380 15326
rect 23324 15262 23326 15314
rect 23378 15262 23380 15314
rect 23100 14466 23156 14476
rect 23324 14420 23380 15262
rect 23436 15316 23492 16492
rect 23548 15874 23604 17836
rect 23660 17780 23716 18398
rect 23660 17714 23716 17724
rect 23548 15822 23550 15874
rect 23602 15822 23604 15874
rect 23548 15810 23604 15822
rect 23660 15988 23716 15998
rect 23660 15426 23716 15932
rect 23660 15374 23662 15426
rect 23714 15374 23716 15426
rect 23660 15362 23716 15374
rect 23436 15260 23604 15316
rect 23548 15148 23604 15260
rect 23436 15092 23604 15148
rect 23436 14980 23492 15092
rect 23436 14914 23492 14924
rect 22764 14366 22766 14418
rect 22818 14366 22820 14418
rect 22764 14354 22820 14366
rect 23212 14364 23380 14420
rect 23548 14418 23604 14430
rect 23548 14366 23550 14418
rect 23602 14366 23604 14418
rect 22988 14308 23044 14318
rect 22988 14214 23044 14252
rect 23212 14306 23268 14364
rect 23436 14308 23492 14318
rect 23212 14254 23214 14306
rect 23266 14254 23268 14306
rect 23100 13636 23156 13646
rect 23212 13636 23268 14254
rect 22428 13634 22596 13636
rect 22428 13582 22430 13634
rect 22482 13582 22596 13634
rect 22428 13580 22596 13582
rect 22428 13570 22484 13580
rect 22540 13188 22596 13580
rect 23100 13634 23268 13636
rect 23100 13582 23102 13634
rect 23154 13582 23268 13634
rect 23100 13580 23268 13582
rect 23324 14306 23492 14308
rect 23324 14254 23438 14306
rect 23490 14254 23492 14306
rect 23324 14252 23492 14254
rect 23100 13570 23156 13580
rect 22672 13356 22936 13366
rect 22728 13300 22776 13356
rect 22832 13300 22880 13356
rect 22672 13290 22936 13300
rect 23324 13188 23380 14252
rect 23436 14242 23492 14252
rect 23548 13972 23604 14366
rect 23548 13906 23604 13916
rect 23436 13748 23492 13758
rect 23436 13654 23492 13692
rect 22540 13132 23380 13188
rect 22092 13122 22148 13132
rect 22764 13074 22820 13132
rect 22764 13022 22766 13074
rect 22818 13022 22820 13074
rect 22764 13010 22820 13022
rect 23548 12964 23604 12974
rect 23436 12962 23604 12964
rect 23436 12910 23550 12962
rect 23602 12910 23604 12962
rect 23436 12908 23604 12910
rect 21868 12562 21924 12572
rect 22204 12740 22260 12750
rect 21980 12292 22036 12302
rect 21980 12066 22036 12236
rect 21980 12014 21982 12066
rect 22034 12014 22036 12066
rect 21980 12002 22036 12014
rect 21756 11890 21812 11900
rect 21980 11396 22036 11406
rect 21980 11302 22036 11340
rect 22204 11394 22260 12684
rect 22428 12740 22484 12750
rect 22428 12292 22484 12684
rect 22428 12198 22484 12236
rect 22988 12738 23044 12750
rect 22988 12686 22990 12738
rect 23042 12686 23044 12738
rect 22540 12180 22596 12190
rect 22988 12180 23044 12686
rect 23436 12628 23492 12908
rect 23548 12898 23604 12908
rect 23436 12562 23492 12572
rect 22540 12178 23044 12180
rect 22540 12126 22542 12178
rect 22594 12126 22990 12178
rect 23042 12126 23044 12178
rect 22540 12124 23044 12126
rect 22540 12114 22596 12124
rect 22988 12114 23044 12124
rect 23436 12178 23492 12190
rect 23436 12126 23438 12178
rect 23490 12126 23492 12178
rect 23212 11956 23268 11966
rect 22204 11342 22206 11394
rect 22258 11342 22260 11394
rect 22204 11284 22260 11342
rect 22540 11844 22596 11854
rect 22540 11394 22596 11788
rect 22672 11788 22936 11798
rect 22728 11732 22776 11788
rect 22832 11732 22880 11788
rect 22672 11722 22936 11732
rect 22540 11342 22542 11394
rect 22594 11342 22596 11394
rect 22540 11330 22596 11342
rect 22764 11396 22820 11406
rect 22204 11218 22260 11228
rect 22764 11170 22820 11340
rect 22764 11118 22766 11170
rect 22818 11118 22820 11170
rect 22764 11060 22820 11118
rect 22876 11284 22932 11294
rect 22876 11172 22932 11228
rect 22876 11116 23156 11172
rect 22764 11004 22932 11060
rect 22764 10724 22820 10734
rect 22764 10630 22820 10668
rect 21644 10558 21646 10610
rect 21698 10558 21700 10610
rect 20860 10386 20916 10398
rect 20860 10334 20862 10386
rect 20914 10334 20916 10386
rect 20636 9774 20638 9826
rect 20690 9774 20692 9826
rect 20412 8418 20468 8428
rect 20076 8370 20132 8382
rect 20076 8318 20078 8370
rect 20130 8318 20132 8370
rect 20076 7476 20132 8318
rect 20636 8258 20692 9774
rect 20748 10276 20804 10286
rect 20748 9714 20804 10220
rect 20748 9662 20750 9714
rect 20802 9662 20804 9714
rect 20748 9650 20804 9662
rect 20860 9380 20916 10334
rect 21644 10276 21700 10558
rect 21644 10210 21700 10220
rect 21980 10500 22036 10510
rect 22204 10500 22260 10510
rect 21980 9826 22036 10444
rect 21980 9774 21982 9826
rect 22034 9774 22036 9826
rect 21980 9762 22036 9774
rect 22092 10498 22260 10500
rect 22092 10446 22206 10498
rect 22258 10446 22260 10498
rect 22092 10444 22260 10446
rect 21532 9716 21588 9726
rect 21532 9622 21588 9660
rect 20860 9314 20916 9324
rect 21644 9602 21700 9614
rect 21644 9550 21646 9602
rect 21698 9550 21700 9602
rect 20636 8206 20638 8258
rect 20690 8206 20692 8258
rect 20636 8194 20692 8206
rect 20860 8930 20916 8942
rect 20860 8878 20862 8930
rect 20914 8878 20916 8930
rect 20860 7924 20916 8878
rect 19852 7364 19908 7374
rect 19852 7270 19908 7308
rect 19964 7140 20020 7150
rect 19964 6914 20020 7084
rect 19964 6862 19966 6914
rect 20018 6862 20020 6914
rect 19964 6850 20020 6862
rect 19852 6020 19908 6030
rect 20076 6020 20132 7420
rect 20188 7700 20244 7710
rect 20188 7252 20244 7644
rect 20860 7700 20916 7868
rect 20860 7634 20916 7644
rect 21084 8818 21140 8830
rect 21084 8766 21086 8818
rect 21138 8766 21140 8818
rect 20188 6914 20244 7196
rect 20188 6862 20190 6914
rect 20242 6862 20244 6914
rect 20188 6850 20244 6862
rect 20412 7474 20468 7486
rect 20412 7422 20414 7474
rect 20466 7422 20468 7474
rect 20412 6132 20468 7422
rect 20860 7364 20916 7374
rect 20860 7270 20916 7308
rect 20636 6914 20692 6926
rect 20636 6862 20638 6914
rect 20690 6862 20692 6914
rect 20524 6692 20580 6702
rect 20524 6598 20580 6636
rect 20636 6468 20692 6862
rect 21084 6916 21140 8766
rect 21308 8818 21364 8830
rect 21308 8766 21310 8818
rect 21362 8766 21364 8818
rect 21308 7028 21364 8766
rect 21644 8820 21700 9550
rect 22092 9044 22148 10444
rect 22204 10434 22260 10444
rect 22316 10500 22372 10510
rect 22316 9266 22372 10444
rect 22876 10500 22932 11004
rect 22876 10434 22932 10444
rect 22988 10948 23044 10958
rect 22988 10610 23044 10892
rect 22988 10558 22990 10610
rect 23042 10558 23044 10610
rect 22988 10388 23044 10558
rect 23100 10388 23156 11116
rect 23212 10724 23268 11900
rect 23324 11394 23380 11406
rect 23324 11342 23326 11394
rect 23378 11342 23380 11394
rect 23324 10948 23380 11342
rect 23324 10882 23380 10892
rect 23436 10836 23492 12126
rect 23548 12180 23604 12190
rect 23548 12086 23604 12124
rect 23660 12178 23716 12190
rect 23660 12126 23662 12178
rect 23714 12126 23716 12178
rect 23212 10668 23380 10724
rect 23212 10388 23268 10398
rect 23100 10332 23212 10388
rect 22988 10322 23044 10332
rect 23212 10322 23268 10332
rect 22672 10220 22936 10230
rect 22728 10164 22776 10220
rect 22832 10164 22880 10220
rect 22672 10154 22936 10164
rect 22988 9828 23044 9838
rect 22316 9214 22318 9266
rect 22370 9214 22372 9266
rect 22316 9202 22372 9214
rect 22540 9714 22596 9726
rect 22540 9662 22542 9714
rect 22594 9662 22596 9714
rect 22428 9044 22484 9054
rect 22540 9044 22596 9662
rect 22092 8988 22372 9044
rect 21644 8754 21700 8764
rect 21756 8818 21812 8830
rect 21756 8766 21758 8818
rect 21810 8766 21812 8818
rect 21756 8428 21812 8766
rect 21756 8372 22260 8428
rect 22204 8258 22260 8372
rect 22204 8206 22206 8258
rect 22258 8206 22260 8258
rect 22204 8194 22260 8206
rect 21308 6962 21364 6972
rect 21420 8034 21476 8046
rect 21420 7982 21422 8034
rect 21474 7982 21476 8034
rect 21084 6850 21140 6860
rect 20636 6402 20692 6412
rect 20748 6578 20804 6590
rect 20748 6526 20750 6578
rect 20802 6526 20804 6578
rect 20412 6066 20468 6076
rect 19852 6018 20132 6020
rect 19852 5966 19854 6018
rect 19906 5966 20132 6018
rect 19852 5964 20132 5966
rect 19852 4340 19908 5964
rect 20300 5236 20356 5246
rect 20300 5142 20356 5180
rect 19852 4274 19908 4284
rect 20412 4450 20468 4462
rect 20412 4398 20414 4450
rect 20466 4398 20468 4450
rect 20412 4340 20468 4398
rect 20412 4274 20468 4284
rect 19852 3556 19908 3566
rect 19740 3500 19852 3556
rect 19852 3462 19908 3500
rect 18396 2594 18452 2604
rect 20748 2548 20804 6526
rect 21084 4900 21140 4910
rect 20972 4452 21028 4490
rect 20972 4386 21028 4396
rect 20860 4340 20916 4350
rect 20860 4246 20916 4284
rect 20972 4228 21028 4238
rect 20972 3666 21028 4172
rect 20972 3614 20974 3666
rect 21026 3614 21028 3666
rect 20972 3602 21028 3614
rect 21084 3554 21140 4844
rect 21420 3780 21476 7982
rect 21756 8036 21812 8046
rect 21756 7942 21812 7980
rect 21644 7476 21700 7486
rect 21644 6018 21700 7420
rect 22316 7474 22372 8988
rect 22428 9042 22596 9044
rect 22428 8990 22430 9042
rect 22482 8990 22596 9042
rect 22428 8988 22596 8990
rect 22876 9716 22932 9726
rect 22428 8482 22484 8988
rect 22876 8820 22932 9660
rect 22988 9042 23044 9772
rect 23324 9604 23380 10668
rect 23436 10498 23492 10780
rect 23436 10446 23438 10498
rect 23490 10446 23492 10498
rect 23436 10434 23492 10446
rect 23660 10052 23716 12126
rect 23772 11620 23828 18956
rect 24444 18674 24500 19294
rect 24444 18622 24446 18674
rect 24498 18622 24500 18674
rect 24444 18610 24500 18622
rect 24556 19346 24948 19348
rect 24556 19294 24894 19346
rect 24946 19294 24948 19346
rect 24556 19292 24948 19294
rect 24108 18450 24164 18462
rect 24108 18398 24110 18450
rect 24162 18398 24164 18450
rect 24108 16548 24164 18398
rect 24556 18228 24612 19292
rect 24892 19282 24948 19292
rect 25452 19346 25508 19358
rect 25452 19294 25454 19346
rect 25506 19294 25508 19346
rect 25452 19012 25508 19294
rect 25452 18946 25508 18956
rect 24668 18676 24724 18686
rect 24668 18582 24724 18620
rect 24780 18564 24836 18574
rect 24780 18450 24836 18508
rect 24780 18398 24782 18450
rect 24834 18398 24836 18450
rect 24780 18386 24836 18398
rect 24444 18172 24612 18228
rect 25228 18338 25284 18350
rect 25228 18286 25230 18338
rect 25282 18286 25284 18338
rect 24220 17780 24276 17790
rect 24220 17106 24276 17724
rect 24220 17054 24222 17106
rect 24274 17054 24276 17106
rect 24220 17042 24276 17054
rect 24444 17106 24500 18172
rect 24444 17054 24446 17106
rect 24498 17054 24500 17106
rect 24444 17042 24500 17054
rect 24556 17556 24612 17566
rect 24556 16770 24612 17500
rect 25228 17108 25284 18286
rect 25676 17332 25732 19852
rect 25788 19234 25844 19246
rect 25788 19182 25790 19234
rect 25842 19182 25844 19234
rect 25788 18676 25844 19182
rect 26348 19236 26404 20076
rect 26460 19236 26516 19246
rect 26348 19234 26516 19236
rect 26348 19182 26462 19234
rect 26514 19182 26516 19234
rect 26348 19180 26516 19182
rect 26460 19170 26516 19180
rect 26124 19012 26180 19022
rect 25788 17444 25844 18620
rect 26012 19010 26180 19012
rect 26012 18958 26126 19010
rect 26178 18958 26180 19010
rect 26012 18956 26180 18958
rect 25900 18452 25956 18462
rect 26012 18452 26068 18956
rect 26124 18946 26180 18956
rect 26348 19012 26404 19022
rect 26348 18918 26404 18956
rect 25900 18450 26068 18452
rect 25900 18398 25902 18450
rect 25954 18398 26068 18450
rect 25900 18396 26068 18398
rect 26124 18452 26180 18462
rect 26460 18452 26516 18462
rect 26124 18450 26516 18452
rect 26124 18398 26126 18450
rect 26178 18398 26462 18450
rect 26514 18398 26516 18450
rect 26124 18396 26516 18398
rect 25900 18386 25956 18396
rect 26124 18386 26180 18396
rect 26460 18386 26516 18396
rect 26572 17666 26628 20860
rect 26684 19124 26740 20972
rect 26684 19058 26740 19068
rect 26908 19124 26964 19134
rect 26908 19030 26964 19068
rect 26684 18564 26740 18574
rect 26684 18470 26740 18508
rect 26572 17614 26574 17666
rect 26626 17614 26628 17666
rect 26572 17602 26628 17614
rect 26796 18450 26852 18462
rect 26796 18398 26798 18450
rect 26850 18398 26852 18450
rect 26796 17556 26852 18398
rect 26796 17490 26852 17500
rect 25900 17444 25956 17454
rect 25788 17388 25900 17444
rect 25900 17378 25956 17388
rect 25676 17276 25844 17332
rect 24556 16718 24558 16770
rect 24610 16718 24612 16770
rect 24556 16706 24612 16718
rect 24668 17052 25284 17108
rect 24108 16482 24164 16492
rect 24444 16324 24500 16334
rect 24332 16212 24388 16222
rect 24108 15316 24164 15326
rect 24108 15222 24164 15260
rect 24220 14530 24276 14542
rect 24220 14478 24222 14530
rect 24274 14478 24276 14530
rect 23884 13860 23940 13870
rect 23884 13766 23940 13804
rect 24220 13748 24276 14478
rect 23996 13692 24220 13748
rect 23884 12740 23940 12750
rect 23884 12646 23940 12684
rect 23996 12402 24052 13692
rect 24220 13682 24276 13692
rect 24332 12404 24388 16156
rect 24444 13524 24500 16268
rect 24556 15316 24612 15326
rect 24668 15316 24724 17052
rect 25340 16996 25396 17006
rect 24780 16884 24836 16894
rect 24780 16322 24836 16828
rect 25340 16770 25396 16940
rect 25676 16884 25732 16894
rect 25676 16790 25732 16828
rect 25340 16718 25342 16770
rect 25394 16718 25396 16770
rect 25340 16706 25396 16718
rect 25452 16772 25508 16782
rect 24780 16270 24782 16322
rect 24834 16270 24836 16322
rect 24780 16258 24836 16270
rect 25340 16548 25396 16558
rect 25116 16212 25172 16222
rect 25116 16118 25172 16156
rect 25340 16100 25396 16492
rect 25228 16098 25396 16100
rect 25228 16046 25342 16098
rect 25394 16046 25396 16098
rect 25228 16044 25396 16046
rect 24556 15314 24724 15316
rect 24556 15262 24558 15314
rect 24610 15262 24724 15314
rect 24556 15260 24724 15262
rect 24780 15876 24836 15886
rect 24556 15250 24612 15260
rect 24444 13458 24500 13468
rect 24556 14532 24612 14542
rect 23996 12350 23998 12402
rect 24050 12350 24052 12402
rect 23996 12338 24052 12350
rect 24220 12348 24388 12404
rect 24444 12962 24500 12974
rect 24444 12910 24446 12962
rect 24498 12910 24500 12962
rect 24220 11620 24276 12348
rect 24332 12180 24388 12190
rect 24332 12086 24388 12124
rect 24444 12068 24500 12910
rect 24556 12292 24612 14476
rect 24668 14530 24724 14542
rect 24668 14478 24670 14530
rect 24722 14478 24724 14530
rect 24668 14308 24724 14478
rect 24668 14242 24724 14252
rect 24780 13970 24836 15820
rect 25116 15204 25172 15214
rect 24892 15092 25172 15148
rect 24892 14642 24948 15092
rect 24892 14590 24894 14642
rect 24946 14590 24948 14642
rect 24892 14578 24948 14590
rect 25228 14644 25284 16044
rect 25340 16034 25396 16044
rect 25340 15876 25396 15886
rect 25452 15876 25508 16716
rect 25396 15820 25508 15876
rect 25564 16770 25620 16782
rect 25564 16718 25566 16770
rect 25618 16718 25620 16770
rect 25340 15538 25396 15820
rect 25340 15486 25342 15538
rect 25394 15486 25396 15538
rect 25340 15474 25396 15486
rect 25452 15316 25508 15326
rect 25452 15222 25508 15260
rect 25564 15148 25620 16718
rect 25340 15092 25620 15148
rect 25340 15090 25396 15092
rect 25340 15038 25342 15090
rect 25394 15038 25396 15090
rect 25340 15026 25396 15038
rect 25340 14644 25396 14654
rect 25228 14642 25396 14644
rect 25228 14590 25342 14642
rect 25394 14590 25396 14642
rect 25228 14588 25396 14590
rect 25340 14578 25396 14588
rect 25452 14532 25508 14542
rect 25452 14438 25508 14476
rect 25228 14308 25284 14318
rect 25228 14214 25284 14252
rect 25788 14084 25844 17276
rect 26908 16100 26964 16110
rect 26012 15986 26068 15998
rect 26012 15934 26014 15986
rect 26066 15934 26068 15986
rect 26012 15314 26068 15934
rect 26012 15262 26014 15314
rect 26066 15262 26068 15314
rect 26012 15204 26068 15262
rect 26012 15138 26068 15148
rect 26124 15874 26180 15886
rect 26124 15822 26126 15874
rect 26178 15822 26180 15874
rect 26124 15540 26180 15822
rect 26348 15876 26404 15886
rect 26348 15782 26404 15820
rect 25900 14868 25956 14878
rect 25900 14530 25956 14812
rect 26124 14644 26180 15484
rect 26908 15426 26964 16044
rect 26908 15374 26910 15426
rect 26962 15374 26964 15426
rect 26908 15362 26964 15374
rect 26460 15316 26516 15326
rect 26460 15314 26628 15316
rect 26460 15262 26462 15314
rect 26514 15262 26628 15314
rect 26460 15260 26628 15262
rect 26460 15250 26516 15260
rect 26572 15148 26628 15260
rect 26124 14578 26180 14588
rect 26460 15092 26628 15148
rect 25900 14478 25902 14530
rect 25954 14478 25956 14530
rect 25900 14466 25956 14478
rect 26460 14308 26516 15092
rect 26572 14644 26628 14654
rect 26628 14588 26852 14644
rect 26572 14578 26628 14588
rect 26460 14214 26516 14252
rect 26572 14420 26628 14430
rect 25788 14018 25844 14028
rect 26348 14084 26404 14094
rect 24780 13918 24782 13970
rect 24834 13918 24836 13970
rect 24780 13906 24836 13918
rect 25228 13972 25284 13982
rect 25228 13878 25284 13916
rect 24668 13860 24724 13870
rect 24668 12964 24724 13804
rect 25564 13746 25620 13758
rect 25564 13694 25566 13746
rect 25618 13694 25620 13746
rect 24668 12870 24724 12908
rect 24780 13524 24836 13534
rect 24780 12852 24836 13468
rect 24892 13412 24948 13422
rect 24892 13074 24948 13356
rect 25564 13188 25620 13694
rect 25900 13746 25956 13758
rect 25900 13694 25902 13746
rect 25954 13694 25956 13746
rect 25900 13188 25956 13694
rect 25564 13132 25956 13188
rect 24892 13022 24894 13074
rect 24946 13022 24948 13074
rect 24892 13010 24948 13022
rect 25676 12964 25732 12974
rect 25676 12870 25732 12908
rect 25116 12852 25172 12862
rect 24780 12796 24948 12852
rect 24556 12198 24612 12236
rect 24444 12002 24500 12012
rect 23772 11564 23940 11620
rect 24220 11564 24724 11620
rect 23772 11394 23828 11406
rect 23772 11342 23774 11394
rect 23826 11342 23828 11394
rect 23772 10612 23828 11342
rect 23772 10518 23828 10556
rect 23660 9986 23716 9996
rect 23660 9828 23716 9838
rect 23660 9734 23716 9772
rect 23324 9538 23380 9548
rect 23548 9714 23604 9726
rect 23548 9662 23550 9714
rect 23602 9662 23604 9714
rect 23100 9156 23156 9166
rect 23548 9156 23604 9662
rect 23156 9100 23604 9156
rect 23100 9062 23156 9100
rect 22988 8990 22990 9042
rect 23042 8990 23044 9042
rect 22988 8978 23044 8990
rect 23436 8932 23492 8942
rect 23436 8838 23492 8876
rect 22876 8764 23156 8820
rect 22672 8652 22936 8662
rect 22728 8596 22776 8652
rect 22832 8596 22880 8652
rect 22672 8586 22936 8596
rect 22428 8430 22430 8482
rect 22482 8430 22484 8482
rect 22428 8418 22484 8430
rect 22764 8260 22820 8270
rect 22764 8166 22820 8204
rect 23100 8258 23156 8764
rect 23100 8206 23102 8258
rect 23154 8206 23156 8258
rect 23100 8148 23156 8206
rect 23100 8082 23156 8092
rect 23324 8484 23380 8494
rect 23100 7700 23156 7710
rect 22316 7422 22318 7474
rect 22370 7422 22372 7474
rect 22316 7410 22372 7422
rect 22988 7476 23044 7486
rect 22988 7382 23044 7420
rect 22672 7084 22936 7094
rect 21868 7028 21924 7038
rect 22728 7028 22776 7084
rect 22832 7028 22880 7084
rect 22672 7018 22936 7028
rect 21868 6578 21924 6972
rect 21868 6526 21870 6578
rect 21922 6526 21924 6578
rect 21868 6514 21924 6526
rect 22764 6916 22820 6926
rect 22764 6690 22820 6860
rect 23100 6802 23156 7644
rect 23100 6750 23102 6802
rect 23154 6750 23156 6802
rect 23100 6738 23156 6750
rect 23212 7250 23268 7262
rect 23212 7198 23214 7250
rect 23266 7198 23268 7250
rect 22764 6638 22766 6690
rect 22818 6638 22820 6690
rect 21644 5966 21646 6018
rect 21698 5966 21700 6018
rect 21644 5954 21700 5966
rect 22428 6468 22484 6478
rect 22092 5908 22148 5918
rect 21980 5906 22148 5908
rect 21980 5854 22094 5906
rect 22146 5854 22148 5906
rect 21980 5852 22148 5854
rect 21980 5572 22036 5852
rect 22092 5842 22148 5852
rect 21420 3714 21476 3724
rect 21756 5516 22036 5572
rect 21756 3666 21812 5516
rect 22316 5122 22372 5134
rect 22316 5070 22318 5122
rect 22370 5070 22372 5122
rect 22316 4676 22372 5070
rect 22316 4610 22372 4620
rect 21980 4340 22036 4350
rect 21980 4246 22036 4284
rect 21756 3614 21758 3666
rect 21810 3614 21812 3666
rect 21756 3602 21812 3614
rect 22316 4004 22372 4014
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 20748 2482 20804 2492
rect 22316 1876 22372 3948
rect 22428 3554 22484 6412
rect 22652 6132 22708 6142
rect 22540 6076 22652 6132
rect 22540 5906 22596 6076
rect 22652 6066 22708 6076
rect 22764 6130 22820 6638
rect 22764 6078 22766 6130
rect 22818 6078 22820 6130
rect 22764 6066 22820 6078
rect 22540 5854 22542 5906
rect 22594 5854 22596 5906
rect 22540 5236 22596 5854
rect 22672 5516 22936 5526
rect 22728 5460 22776 5516
rect 22832 5460 22880 5516
rect 22672 5450 22936 5460
rect 22540 5170 22596 5180
rect 22764 5348 22820 5358
rect 22652 5122 22708 5134
rect 22652 5070 22654 5122
rect 22706 5070 22708 5122
rect 22652 4564 22708 5070
rect 22652 4498 22708 4508
rect 22764 4338 22820 5292
rect 22764 4286 22766 4338
rect 22818 4286 22820 4338
rect 22764 4274 22820 4286
rect 23100 5124 23156 5134
rect 22876 4228 22932 4238
rect 22876 4134 22932 4172
rect 22672 3948 22936 3958
rect 22728 3892 22776 3948
rect 22832 3892 22880 3948
rect 22672 3882 22936 3892
rect 22428 3502 22430 3554
rect 22482 3502 22484 3554
rect 22428 3490 22484 3502
rect 22988 3556 23044 3566
rect 23100 3556 23156 5068
rect 23212 5012 23268 7198
rect 23324 6466 23380 8428
rect 23772 8148 23828 8158
rect 23548 7474 23604 7486
rect 23548 7422 23550 7474
rect 23602 7422 23604 7474
rect 23548 6804 23604 7422
rect 23324 6414 23326 6466
rect 23378 6414 23380 6466
rect 23324 6402 23380 6414
rect 23436 6748 23604 6804
rect 23436 6132 23492 6748
rect 23436 6066 23492 6076
rect 23548 6580 23604 6590
rect 23548 6020 23604 6524
rect 23660 6020 23716 6030
rect 23548 6018 23716 6020
rect 23548 5966 23662 6018
rect 23714 5966 23716 6018
rect 23548 5964 23716 5966
rect 23660 5954 23716 5964
rect 23324 5572 23380 5582
rect 23324 5234 23380 5516
rect 23324 5182 23326 5234
rect 23378 5182 23380 5234
rect 23324 5170 23380 5182
rect 23772 5122 23828 8092
rect 23884 7588 23940 11564
rect 24220 11396 24276 11406
rect 24556 11396 24612 11406
rect 24220 11394 24388 11396
rect 24220 11342 24222 11394
rect 24274 11342 24388 11394
rect 24220 11340 24388 11342
rect 24220 11330 24276 11340
rect 24332 10610 24388 11340
rect 24556 11302 24612 11340
rect 24332 10558 24334 10610
rect 24386 10558 24388 10610
rect 24332 9940 24388 10558
rect 24332 9874 24388 9884
rect 24556 9156 24612 9166
rect 24556 9062 24612 9100
rect 24108 9044 24164 9054
rect 23996 8820 24052 8830
rect 23996 8258 24052 8764
rect 24108 8484 24164 8988
rect 24108 8418 24164 8428
rect 24332 8930 24388 8942
rect 24332 8878 24334 8930
rect 24386 8878 24388 8930
rect 24332 8260 24388 8878
rect 23996 8206 23998 8258
rect 24050 8206 24052 8258
rect 23996 8194 24052 8206
rect 24220 8258 24388 8260
rect 24220 8206 24334 8258
rect 24386 8206 24388 8258
rect 24220 8204 24388 8206
rect 23884 7522 23940 7532
rect 23772 5070 23774 5122
rect 23826 5070 23828 5122
rect 23772 5058 23828 5070
rect 24220 5122 24276 8204
rect 24332 8194 24388 8204
rect 24220 5070 24222 5122
rect 24274 5070 24276 5122
rect 24220 5058 24276 5070
rect 24332 6466 24388 6478
rect 24332 6414 24334 6466
rect 24386 6414 24388 6466
rect 24332 5124 24388 6414
rect 24668 6132 24724 11564
rect 24668 6038 24724 6076
rect 24332 5058 24388 5068
rect 24780 5908 24836 5918
rect 23212 4946 23268 4956
rect 23996 4900 24052 4910
rect 23996 4450 24052 4844
rect 24332 4564 24388 4574
rect 24332 4470 24388 4508
rect 23996 4398 23998 4450
rect 24050 4398 24052 4450
rect 23996 4386 24052 4398
rect 24668 4452 24724 4462
rect 24780 4452 24836 5852
rect 24892 4564 24948 12796
rect 25116 12758 25172 12796
rect 25340 12850 25396 12862
rect 25340 12798 25342 12850
rect 25394 12798 25396 12850
rect 25340 12628 25396 12798
rect 25676 12738 25732 12750
rect 25676 12686 25678 12738
rect 25730 12686 25732 12738
rect 25676 12628 25732 12686
rect 25340 12572 25732 12628
rect 25340 12292 25396 12302
rect 25340 12066 25396 12236
rect 25340 12014 25342 12066
rect 25394 12014 25396 12066
rect 25340 12002 25396 12014
rect 25564 12180 25620 12190
rect 25788 12180 25844 13132
rect 26012 12962 26068 12974
rect 26012 12910 26014 12962
rect 26066 12910 26068 12962
rect 25564 12178 25844 12180
rect 25564 12126 25566 12178
rect 25618 12126 25844 12178
rect 25564 12124 25844 12126
rect 25900 12852 25956 12862
rect 25900 12180 25956 12796
rect 25228 11396 25284 11406
rect 25284 11340 25508 11396
rect 25228 11302 25284 11340
rect 25340 10836 25396 10846
rect 25340 10742 25396 10780
rect 25228 10610 25284 10622
rect 25228 10558 25230 10610
rect 25282 10558 25284 10610
rect 25228 10052 25284 10558
rect 25228 9938 25284 9996
rect 25228 9886 25230 9938
rect 25282 9886 25284 9938
rect 25228 9874 25284 9886
rect 25452 9044 25508 11340
rect 25564 10834 25620 12124
rect 25676 11284 25732 11294
rect 25900 11284 25956 12124
rect 26012 11508 26068 12910
rect 26236 12964 26292 12974
rect 26348 12964 26404 14028
rect 26460 13748 26516 13758
rect 26572 13748 26628 14364
rect 26796 14418 26852 14588
rect 26796 14366 26798 14418
rect 26850 14366 26852 14418
rect 26796 14354 26852 14366
rect 26460 13746 26628 13748
rect 26460 13694 26462 13746
rect 26514 13694 26628 13746
rect 26460 13692 26628 13694
rect 26684 14196 26740 14206
rect 26460 13682 26516 13692
rect 26460 12964 26516 12974
rect 26348 12962 26516 12964
rect 26348 12910 26462 12962
rect 26514 12910 26516 12962
rect 26348 12908 26516 12910
rect 26236 12870 26292 12908
rect 26460 12898 26516 12908
rect 26684 12962 26740 14140
rect 27020 13634 27076 13646
rect 27020 13582 27022 13634
rect 27074 13582 27076 13634
rect 26684 12910 26686 12962
rect 26738 12910 26740 12962
rect 26684 12898 26740 12910
rect 26908 13188 26964 13198
rect 26908 12850 26964 13132
rect 26908 12798 26910 12850
rect 26962 12798 26964 12850
rect 26908 12786 26964 12798
rect 27020 12850 27076 13582
rect 27020 12798 27022 12850
rect 27074 12798 27076 12850
rect 26796 12516 26852 12526
rect 26236 12178 26292 12190
rect 26236 12126 26238 12178
rect 26290 12126 26292 12178
rect 26012 11442 26068 11452
rect 26124 12068 26180 12078
rect 26012 11284 26068 11294
rect 25900 11282 26068 11284
rect 25900 11230 26014 11282
rect 26066 11230 26068 11282
rect 25900 11228 26068 11230
rect 25676 11190 25732 11228
rect 26012 11218 26068 11228
rect 26124 11060 26180 12012
rect 26236 11956 26292 12126
rect 26236 11890 26292 11900
rect 26460 12068 26516 12078
rect 26348 11394 26404 11406
rect 26348 11342 26350 11394
rect 26402 11342 26404 11394
rect 26124 11004 26292 11060
rect 25564 10782 25566 10834
rect 25618 10782 25620 10834
rect 25564 10770 25620 10782
rect 26124 10836 26180 10846
rect 26124 10742 26180 10780
rect 26124 10610 26180 10622
rect 26124 10558 26126 10610
rect 26178 10558 26180 10610
rect 26124 10052 26180 10558
rect 26124 9986 26180 9996
rect 26012 9940 26068 9950
rect 26012 9846 26068 9884
rect 25788 9826 25844 9838
rect 25788 9774 25790 9826
rect 25842 9774 25844 9826
rect 25676 9044 25732 9054
rect 25452 9042 25732 9044
rect 25452 8990 25678 9042
rect 25730 8990 25732 9042
rect 25452 8988 25732 8990
rect 25676 8978 25732 8988
rect 25788 8820 25844 9774
rect 26124 9826 26180 9838
rect 26124 9774 26126 9826
rect 26178 9774 26180 9826
rect 25900 9492 25956 9502
rect 25900 9042 25956 9436
rect 25900 8990 25902 9042
rect 25954 8990 25956 9042
rect 25900 8932 25956 8990
rect 26124 9044 26180 9774
rect 26124 8978 26180 8988
rect 25900 8866 25956 8876
rect 26236 8820 26292 11004
rect 26348 10948 26404 11342
rect 26348 10882 26404 10892
rect 26460 9940 26516 12012
rect 26684 11508 26740 11518
rect 25788 8754 25844 8764
rect 26124 8764 26292 8820
rect 26348 9884 26516 9940
rect 26572 11394 26628 11406
rect 26572 11342 26574 11394
rect 26626 11342 26628 11394
rect 25676 8708 25732 8718
rect 25452 8652 25676 8708
rect 25228 8372 25284 8382
rect 25228 7698 25284 8316
rect 25228 7646 25230 7698
rect 25282 7646 25284 7698
rect 25228 7634 25284 7646
rect 25228 6578 25284 6590
rect 25228 6526 25230 6578
rect 25282 6526 25284 6578
rect 25228 6356 25284 6526
rect 25284 6300 25396 6356
rect 25228 6290 25284 6300
rect 25228 6018 25284 6030
rect 25228 5966 25230 6018
rect 25282 5966 25284 6018
rect 25228 5684 25284 5966
rect 25340 5906 25396 6300
rect 25340 5854 25342 5906
rect 25394 5854 25396 5906
rect 25340 5842 25396 5854
rect 25116 5628 25284 5684
rect 24892 4498 24948 4508
rect 25004 5124 25060 5134
rect 24668 4450 24836 4452
rect 24668 4398 24670 4450
rect 24722 4398 24836 4450
rect 24668 4396 24836 4398
rect 24668 4386 24724 4396
rect 23996 3668 24052 3678
rect 23996 3574 24052 3612
rect 22988 3554 23156 3556
rect 22988 3502 22990 3554
rect 23042 3502 23156 3554
rect 22988 3500 23156 3502
rect 25004 3556 25060 5068
rect 25116 4900 25172 5628
rect 25116 4834 25172 4844
rect 25228 5460 25284 5470
rect 25228 4338 25284 5404
rect 25340 5236 25396 5246
rect 25452 5236 25508 8652
rect 25676 8642 25732 8652
rect 25564 8372 25620 8382
rect 25564 8278 25620 8316
rect 25900 8260 25956 8270
rect 25900 8166 25956 8204
rect 26012 8258 26068 8270
rect 26012 8206 26014 8258
rect 26066 8206 26068 8258
rect 25788 7364 25844 7374
rect 26012 7364 26068 8206
rect 26124 8148 26180 8764
rect 26348 8708 26404 9884
rect 26348 8642 26404 8652
rect 26460 9716 26516 9726
rect 26572 9716 26628 11342
rect 26684 10836 26740 11452
rect 26796 11172 26852 12460
rect 27020 12516 27076 12798
rect 27020 12068 27076 12460
rect 27132 12964 27188 23548
rect 27580 23492 27636 23662
rect 27692 23716 27748 23726
rect 27692 23622 27748 23660
rect 28028 23716 28084 23726
rect 28028 23622 28084 23660
rect 27916 23604 27972 23614
rect 27244 23436 27636 23492
rect 27804 23548 27916 23604
rect 27244 22708 27300 23436
rect 27356 23268 27412 23278
rect 27692 23268 27748 23278
rect 27804 23268 27860 23548
rect 27916 23538 27972 23548
rect 27356 23266 27860 23268
rect 27356 23214 27358 23266
rect 27410 23214 27694 23266
rect 27746 23214 27860 23266
rect 27356 23212 27860 23214
rect 28028 23380 28084 23390
rect 28028 23266 28084 23324
rect 28028 23214 28030 23266
rect 28082 23214 28084 23266
rect 27356 23202 27412 23212
rect 27692 23202 27748 23212
rect 28028 23202 28084 23214
rect 28252 23266 28308 23884
rect 28476 23874 28532 23884
rect 28588 23940 28644 23950
rect 28588 23846 28644 23884
rect 28252 23214 28254 23266
rect 28306 23214 28308 23266
rect 28252 23202 28308 23214
rect 27804 23044 27860 23054
rect 27804 22950 27860 22988
rect 27244 22594 27300 22652
rect 27244 22542 27246 22594
rect 27298 22542 27300 22594
rect 27244 22530 27300 22542
rect 27356 22932 27412 22942
rect 27356 22596 27412 22876
rect 27356 22370 27412 22540
rect 27356 22318 27358 22370
rect 27410 22318 27412 22370
rect 27356 22306 27412 22318
rect 27580 22370 27636 22382
rect 27580 22318 27582 22370
rect 27634 22318 27636 22370
rect 27580 22260 27636 22318
rect 27580 22194 27636 22204
rect 28364 22370 28420 22382
rect 28364 22318 28366 22370
rect 28418 22318 28420 22370
rect 28028 22146 28084 22158
rect 28028 22094 28030 22146
rect 28082 22094 28084 22146
rect 27244 21586 27300 21598
rect 27244 21534 27246 21586
rect 27298 21534 27300 21586
rect 27244 16100 27300 21534
rect 28028 21476 28084 22094
rect 28028 21410 28084 21420
rect 28140 21586 28196 21598
rect 28140 21534 28142 21586
rect 28194 21534 28196 21586
rect 28028 21140 28084 21150
rect 28028 20020 28084 21084
rect 28140 20132 28196 21534
rect 28140 20066 28196 20076
rect 28028 19954 28084 19964
rect 28364 20020 28420 22318
rect 28588 22372 28644 22410
rect 28588 22306 28644 22316
rect 28588 22148 28644 22158
rect 28588 21586 28644 22092
rect 28588 21534 28590 21586
rect 28642 21534 28644 21586
rect 28588 21522 28644 21534
rect 28700 21364 28756 25004
rect 28812 23828 28868 25116
rect 28812 23762 28868 23772
rect 28924 23548 28980 28812
rect 29260 28532 29316 28542
rect 29260 26964 29316 28476
rect 29148 25508 29204 25518
rect 29148 25414 29204 25452
rect 29148 25060 29204 25070
rect 29148 24834 29204 25004
rect 29260 24948 29316 26908
rect 29372 27524 29428 27534
rect 29372 26290 29428 27468
rect 29372 26238 29374 26290
rect 29426 26238 29428 26290
rect 29372 26226 29428 26238
rect 29596 25618 29652 29260
rect 29708 29204 29764 29932
rect 29825 29820 30089 29830
rect 29881 29764 29929 29820
rect 29985 29764 30033 29820
rect 29825 29754 30089 29764
rect 30156 29652 30212 30380
rect 31388 30212 31444 30222
rect 31388 30118 31444 30156
rect 29932 29596 30212 29652
rect 29932 29538 29988 29596
rect 29932 29486 29934 29538
rect 29986 29486 29988 29538
rect 29932 29474 29988 29486
rect 30604 29428 30660 29438
rect 30604 29334 30660 29372
rect 30268 29314 30324 29326
rect 30268 29262 30270 29314
rect 30322 29262 30324 29314
rect 30268 29204 30324 29262
rect 31388 29314 31444 29326
rect 31388 29262 31390 29314
rect 31442 29262 31444 29314
rect 31276 29204 31332 29214
rect 29708 29148 30100 29204
rect 30044 28754 30100 29148
rect 30044 28702 30046 28754
rect 30098 28702 30100 28754
rect 30044 28690 30100 28702
rect 30268 29202 31332 29204
rect 30268 29150 31278 29202
rect 31330 29150 31332 29202
rect 30268 29148 31332 29150
rect 29825 28252 30089 28262
rect 29881 28196 29929 28252
rect 29985 28196 30033 28252
rect 29825 28186 30089 28196
rect 30268 27970 30324 29148
rect 31276 29138 31332 29148
rect 31388 28980 31444 29262
rect 30492 28924 31444 28980
rect 30492 28754 30548 28924
rect 31164 28756 31220 28766
rect 31500 28756 31556 30380
rect 31612 30324 31668 30942
rect 31724 30434 31780 31500
rect 31836 31444 31892 31838
rect 33292 31780 33348 31790
rect 33292 31686 33348 31724
rect 32732 31668 32788 31678
rect 33404 31668 33460 31678
rect 32732 31666 33236 31668
rect 32732 31614 32734 31666
rect 32786 31614 33236 31666
rect 32732 31612 33236 31614
rect 32732 31602 32788 31612
rect 32508 31556 32564 31566
rect 32508 31462 32564 31500
rect 31836 31388 32004 31444
rect 31836 31220 31892 31230
rect 31836 30882 31892 31164
rect 31836 30830 31838 30882
rect 31890 30830 31892 30882
rect 31836 30818 31892 30830
rect 31836 30548 31892 30558
rect 31948 30548 32004 31388
rect 33180 31218 33236 31612
rect 33404 31574 33460 31612
rect 33180 31166 33182 31218
rect 33234 31166 33236 31218
rect 33180 31154 33236 31166
rect 33292 31108 33348 31118
rect 33292 31014 33348 31052
rect 32284 30884 32340 30894
rect 33068 30884 33124 30894
rect 32284 30882 33124 30884
rect 32284 30830 32286 30882
rect 32338 30830 33070 30882
rect 33122 30830 33124 30882
rect 32284 30828 33124 30830
rect 32284 30818 32340 30828
rect 33068 30818 33124 30828
rect 31892 30492 32004 30548
rect 31836 30482 31892 30492
rect 31724 30382 31726 30434
rect 31778 30382 31780 30434
rect 31724 30370 31780 30382
rect 31612 30098 31668 30268
rect 31948 30212 32004 30492
rect 31948 30146 32004 30156
rect 32396 30660 32452 30670
rect 32396 30210 32452 30604
rect 33180 30212 33236 30222
rect 32396 30158 32398 30210
rect 32450 30158 32452 30210
rect 32396 30146 32452 30158
rect 33068 30210 33236 30212
rect 33068 30158 33182 30210
rect 33234 30158 33236 30210
rect 33068 30156 33236 30158
rect 31612 30046 31614 30098
rect 31666 30046 31668 30098
rect 31612 30034 31668 30046
rect 32060 30100 32116 30110
rect 31948 29764 32004 29774
rect 31948 29650 32004 29708
rect 31948 29598 31950 29650
rect 32002 29598 32004 29650
rect 31948 29586 32004 29598
rect 32060 29650 32116 30044
rect 33068 29764 33124 30156
rect 33180 30146 33236 30156
rect 32060 29598 32062 29650
rect 32114 29598 32116 29650
rect 32060 29586 32116 29598
rect 32396 29652 32452 29662
rect 32956 29652 33012 29662
rect 32396 29558 32452 29596
rect 32844 29596 32956 29652
rect 31612 29428 31668 29438
rect 31612 28868 31668 29372
rect 32172 29428 32228 29438
rect 32172 29334 32228 29372
rect 31612 28802 31668 28812
rect 30492 28702 30494 28754
rect 30546 28702 30548 28754
rect 30492 28690 30548 28702
rect 30604 28754 31220 28756
rect 30604 28702 31166 28754
rect 31218 28702 31220 28754
rect 30604 28700 31220 28702
rect 30604 28642 30660 28700
rect 31164 28690 31220 28700
rect 31388 28700 31556 28756
rect 30604 28590 30606 28642
rect 30658 28590 30660 28642
rect 30604 28578 30660 28590
rect 30268 27918 30270 27970
rect 30322 27918 30324 27970
rect 30268 27906 30324 27918
rect 31276 28418 31332 28430
rect 31276 28366 31278 28418
rect 31330 28366 31332 28418
rect 30940 27858 30996 27870
rect 30940 27806 30942 27858
rect 30994 27806 30996 27858
rect 30940 27188 30996 27806
rect 31276 27748 31332 28366
rect 31276 27682 31332 27692
rect 31388 27524 31444 28700
rect 32844 28644 32900 29596
rect 32956 29586 33012 29596
rect 32732 28642 32900 28644
rect 32732 28590 32846 28642
rect 32898 28590 32900 28642
rect 32732 28588 32900 28590
rect 31500 28532 31556 28542
rect 31500 28530 31780 28532
rect 31500 28478 31502 28530
rect 31554 28478 31780 28530
rect 31500 28476 31780 28478
rect 31500 28466 31556 28476
rect 30716 27186 30996 27188
rect 30716 27134 30942 27186
rect 30994 27134 30996 27186
rect 30716 27132 30996 27134
rect 30492 26962 30548 26974
rect 30492 26910 30494 26962
rect 30546 26910 30548 26962
rect 30492 26908 30548 26910
rect 30044 26852 30100 26862
rect 30268 26852 30548 26908
rect 30100 26796 30212 26852
rect 30044 26758 30100 26796
rect 29825 26684 30089 26694
rect 29881 26628 29929 26684
rect 29985 26628 30033 26684
rect 29825 26618 30089 26628
rect 30156 25732 30212 26796
rect 29596 25566 29598 25618
rect 29650 25566 29652 25618
rect 29596 25554 29652 25566
rect 30044 25676 30212 25732
rect 30044 25506 30100 25676
rect 30044 25454 30046 25506
rect 30098 25454 30100 25506
rect 29820 25394 29876 25406
rect 29820 25342 29822 25394
rect 29874 25342 29876 25394
rect 29820 25284 29876 25342
rect 29708 25228 29876 25284
rect 30044 25284 30100 25454
rect 29596 25172 29652 25182
rect 29708 25172 29764 25228
rect 30044 25218 30100 25228
rect 30156 25508 30212 25518
rect 29652 25116 29764 25172
rect 29596 25106 29652 25116
rect 29260 24892 29428 24948
rect 29148 24782 29150 24834
rect 29202 24782 29204 24834
rect 29148 24770 29204 24782
rect 29260 24724 29316 24734
rect 29260 24630 29316 24668
rect 29372 24164 29428 24892
rect 29708 24724 29764 25116
rect 29825 25116 30089 25126
rect 29881 25060 29929 25116
rect 29985 25060 30033 25116
rect 29825 25050 30089 25060
rect 29708 24658 29764 24668
rect 29820 24722 29876 24734
rect 29820 24670 29822 24722
rect 29874 24670 29876 24722
rect 29820 24500 29876 24670
rect 29820 24434 29876 24444
rect 29372 24108 29764 24164
rect 28588 21308 28756 21364
rect 28812 23492 28980 23548
rect 29260 23938 29316 23950
rect 29484 23940 29540 23950
rect 29260 23886 29262 23938
rect 29314 23886 29316 23938
rect 29260 23604 29316 23886
rect 29260 23538 29316 23548
rect 29372 23938 29540 23940
rect 29372 23886 29486 23938
rect 29538 23886 29540 23938
rect 29372 23884 29540 23886
rect 28476 20804 28532 20814
rect 28476 20710 28532 20748
rect 28364 19954 28420 19964
rect 28140 19908 28196 19918
rect 28140 19814 28196 19852
rect 28588 19906 28644 21308
rect 28588 19854 28590 19906
rect 28642 19854 28644 19906
rect 28588 19842 28644 19854
rect 28700 20020 28756 20030
rect 28588 19348 28644 19358
rect 28700 19348 28756 19964
rect 28588 19346 28756 19348
rect 28588 19294 28590 19346
rect 28642 19294 28756 19346
rect 28588 19292 28756 19294
rect 28588 19282 28644 19292
rect 28140 19234 28196 19246
rect 28140 19182 28142 19234
rect 28194 19182 28196 19234
rect 28140 19124 28196 19182
rect 28140 19058 28196 19068
rect 28476 19236 28532 19246
rect 28476 18564 28532 19180
rect 28588 18564 28644 18574
rect 28476 18562 28644 18564
rect 28476 18510 28590 18562
rect 28642 18510 28644 18562
rect 28476 18508 28644 18510
rect 28588 18498 28644 18508
rect 27916 18450 27972 18462
rect 27916 18398 27918 18450
rect 27970 18398 27972 18450
rect 27916 18228 27972 18398
rect 28364 18450 28420 18462
rect 28364 18398 28366 18450
rect 28418 18398 28420 18450
rect 27916 18162 27972 18172
rect 28028 18340 28084 18350
rect 28364 18340 28420 18398
rect 28476 18340 28532 18350
rect 28364 18284 28476 18340
rect 28028 17778 28084 18284
rect 28476 18274 28532 18284
rect 28028 17726 28030 17778
rect 28082 17726 28084 17778
rect 28028 17714 28084 17726
rect 27356 17666 27412 17678
rect 27916 17668 27972 17678
rect 27356 17614 27358 17666
rect 27410 17614 27412 17666
rect 27356 16884 27412 17614
rect 27804 17612 27916 17668
rect 27356 16882 27524 16884
rect 27356 16830 27358 16882
rect 27410 16830 27524 16882
rect 27356 16828 27524 16830
rect 27356 16818 27412 16828
rect 27356 16660 27412 16670
rect 27356 16566 27412 16604
rect 27356 16324 27412 16334
rect 27468 16324 27524 16828
rect 27804 16770 27860 17612
rect 27916 17574 27972 17612
rect 27804 16718 27806 16770
rect 27858 16718 27860 16770
rect 27804 16706 27860 16718
rect 28364 16882 28420 16894
rect 28364 16830 28366 16882
rect 28418 16830 28420 16882
rect 27356 16322 27524 16324
rect 27356 16270 27358 16322
rect 27410 16270 27524 16322
rect 27356 16268 27524 16270
rect 28364 16322 28420 16830
rect 28364 16270 28366 16322
rect 28418 16270 28420 16322
rect 27356 16258 27412 16268
rect 28364 16258 28420 16270
rect 28476 16660 28532 16670
rect 27580 16210 27636 16222
rect 27580 16158 27582 16210
rect 27634 16158 27636 16210
rect 27580 16100 27636 16158
rect 27244 16044 27524 16100
rect 27244 15876 27300 15886
rect 27468 15876 27524 16044
rect 27580 16034 27636 16044
rect 27692 16100 27748 16110
rect 28252 16100 28308 16110
rect 27692 16098 28196 16100
rect 27692 16046 27694 16098
rect 27746 16046 28196 16098
rect 27692 16044 28196 16046
rect 27692 16034 27748 16044
rect 28140 15876 28196 16044
rect 28252 16006 28308 16044
rect 28364 15876 28420 15886
rect 27468 15820 27748 15876
rect 28140 15874 28420 15876
rect 28140 15822 28366 15874
rect 28418 15822 28420 15874
rect 28140 15820 28420 15822
rect 27244 15426 27300 15820
rect 27244 15374 27246 15426
rect 27298 15374 27300 15426
rect 27244 15362 27300 15374
rect 27356 15428 27412 15438
rect 27580 15428 27636 15438
rect 27356 15426 27524 15428
rect 27356 15374 27358 15426
rect 27410 15374 27524 15426
rect 27356 15372 27524 15374
rect 27356 15362 27412 15372
rect 27356 15204 27412 15214
rect 27356 14642 27412 15148
rect 27468 15148 27524 15372
rect 27580 15334 27636 15372
rect 27468 15092 27636 15148
rect 27356 14590 27358 14642
rect 27410 14590 27412 14642
rect 27356 14578 27412 14590
rect 27356 14084 27412 14094
rect 27356 13970 27412 14028
rect 27356 13918 27358 13970
rect 27410 13918 27412 13970
rect 27356 13906 27412 13918
rect 27132 12292 27188 12908
rect 27468 12850 27524 12862
rect 27468 12798 27470 12850
rect 27522 12798 27524 12850
rect 27132 12198 27188 12236
rect 27356 12738 27412 12750
rect 27356 12686 27358 12738
rect 27410 12686 27412 12738
rect 27020 12002 27076 12012
rect 27244 12178 27300 12190
rect 27244 12126 27246 12178
rect 27298 12126 27300 12178
rect 26908 11844 26964 11854
rect 26908 11396 26964 11788
rect 27020 11620 27076 11630
rect 27020 11506 27076 11564
rect 27020 11454 27022 11506
rect 27074 11454 27076 11506
rect 27020 11442 27076 11454
rect 26908 11302 26964 11340
rect 27132 11396 27188 11406
rect 27132 11302 27188 11340
rect 26796 11116 27076 11172
rect 26908 10836 26964 10846
rect 26684 10834 26964 10836
rect 26684 10782 26910 10834
rect 26962 10782 26964 10834
rect 26684 10780 26964 10782
rect 26908 10770 26964 10780
rect 27020 10724 27076 11116
rect 27244 10948 27300 12126
rect 27356 11396 27412 12686
rect 27468 12740 27524 12798
rect 27468 12674 27524 12684
rect 27580 12068 27636 15092
rect 27580 11974 27636 12012
rect 27692 11844 27748 15820
rect 28140 15652 28196 15662
rect 28028 15428 28084 15438
rect 28028 15334 28084 15372
rect 27916 15316 27972 15326
rect 27916 15148 27972 15260
rect 27804 15092 27860 15102
rect 27916 15092 28084 15148
rect 27804 14756 27860 15036
rect 27804 14690 27860 14700
rect 27916 14420 27972 14430
rect 27916 14326 27972 14364
rect 28028 13970 28084 15092
rect 28028 13918 28030 13970
rect 28082 13918 28084 13970
rect 28028 13906 28084 13918
rect 28028 12740 28084 12750
rect 27692 11778 27748 11788
rect 27804 12292 27860 12302
rect 27804 11506 27860 12236
rect 27916 12180 27972 12190
rect 27916 12086 27972 12124
rect 27804 11454 27806 11506
rect 27858 11454 27860 11506
rect 27804 11442 27860 11454
rect 27356 11340 27748 11396
rect 27356 11172 27412 11182
rect 27356 11078 27412 11116
rect 27020 10658 27076 10668
rect 27132 10836 27188 10846
rect 27020 9828 27076 9838
rect 27020 9734 27076 9772
rect 26516 9660 26628 9716
rect 26684 9714 26740 9726
rect 26684 9662 26686 9714
rect 26738 9662 26740 9714
rect 26124 8082 26180 8092
rect 26236 8258 26292 8270
rect 26236 8206 26238 8258
rect 26290 8206 26292 8258
rect 25788 7362 26068 7364
rect 25788 7310 25790 7362
rect 25842 7310 26068 7362
rect 25788 7308 26068 7310
rect 25340 5234 25508 5236
rect 25340 5182 25342 5234
rect 25394 5182 25508 5234
rect 25340 5180 25508 5182
rect 25564 7252 25620 7262
rect 25340 5170 25396 5180
rect 25564 5012 25620 7196
rect 25788 6692 25844 7308
rect 26236 7252 26292 8206
rect 26236 7186 26292 7196
rect 26348 8258 26404 8270
rect 26348 8206 26350 8258
rect 26402 8206 26404 8258
rect 25788 5460 25844 6636
rect 26124 6690 26180 6702
rect 26124 6638 26126 6690
rect 26178 6638 26180 6690
rect 26124 6580 26180 6638
rect 26124 6514 26180 6524
rect 26012 5908 26068 5918
rect 26012 5814 26068 5852
rect 25788 5394 25844 5404
rect 26236 5684 26292 5694
rect 25676 5348 25732 5358
rect 25676 5234 25732 5292
rect 25676 5182 25678 5234
rect 25730 5182 25732 5234
rect 25676 5170 25732 5182
rect 26236 5346 26292 5628
rect 26236 5294 26238 5346
rect 26290 5294 26292 5346
rect 25900 5122 25956 5134
rect 25900 5070 25902 5122
rect 25954 5070 25956 5122
rect 25564 4956 25732 5012
rect 25452 4900 25508 4910
rect 25508 4844 25620 4900
rect 25452 4834 25508 4844
rect 25452 4676 25508 4686
rect 25452 4562 25508 4620
rect 25452 4510 25454 4562
rect 25506 4510 25508 4562
rect 25452 4498 25508 4510
rect 25564 4452 25620 4844
rect 25564 4386 25620 4396
rect 25676 4676 25732 4956
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4274 25284 4286
rect 25564 4228 25620 4238
rect 25676 4228 25732 4620
rect 25564 4226 25732 4228
rect 25564 4174 25566 4226
rect 25618 4174 25732 4226
rect 25564 4172 25732 4174
rect 25564 4162 25620 4172
rect 22988 3490 23044 3500
rect 25004 3462 25060 3500
rect 25676 3444 25732 3482
rect 25676 3378 25732 3388
rect 25900 2884 25956 5070
rect 26236 4338 26292 5294
rect 26348 5682 26404 8206
rect 26460 6020 26516 9660
rect 26684 9156 26740 9662
rect 27132 9714 27188 10780
rect 27244 9938 27300 10892
rect 27692 10836 27748 11340
rect 27356 10780 27636 10836
rect 27692 10780 27972 10836
rect 27356 10724 27412 10780
rect 27356 10630 27412 10668
rect 27468 10610 27524 10622
rect 27468 10558 27470 10610
rect 27522 10558 27524 10610
rect 27244 9886 27246 9938
rect 27298 9886 27300 9938
rect 27244 9874 27300 9886
rect 27356 10164 27412 10174
rect 27132 9662 27134 9714
rect 27186 9662 27188 9714
rect 27132 9650 27188 9662
rect 27020 9604 27076 9614
rect 26460 5954 26516 5964
rect 26572 7812 26628 7822
rect 26572 5906 26628 7756
rect 26684 7028 26740 9100
rect 26908 9380 26964 9390
rect 26908 9042 26964 9324
rect 26908 8990 26910 9042
rect 26962 8990 26964 9042
rect 26908 8978 26964 8990
rect 26796 8820 26852 8830
rect 26796 8726 26852 8764
rect 27020 8146 27076 9548
rect 27020 8094 27022 8146
rect 27074 8094 27076 8146
rect 27020 8082 27076 8094
rect 27132 9268 27188 9278
rect 27132 8036 27188 9212
rect 27356 9044 27412 10108
rect 27132 7970 27188 7980
rect 27244 8988 27412 9044
rect 27244 8260 27300 8988
rect 27356 8820 27412 8830
rect 27468 8820 27524 10558
rect 27580 9268 27636 10780
rect 27804 10610 27860 10622
rect 27804 10558 27806 10610
rect 27858 10558 27860 10610
rect 27804 9492 27860 10558
rect 27916 9938 27972 10780
rect 27916 9886 27918 9938
rect 27970 9886 27972 9938
rect 27916 9604 27972 9886
rect 27916 9538 27972 9548
rect 27804 9426 27860 9436
rect 28028 9268 28084 12684
rect 28140 11396 28196 15596
rect 28252 15314 28308 15326
rect 28252 15262 28254 15314
rect 28306 15262 28308 15314
rect 28252 14530 28308 15262
rect 28364 14754 28420 15820
rect 28364 14702 28366 14754
rect 28418 14702 28420 14754
rect 28364 14690 28420 14702
rect 28476 15314 28532 16604
rect 28812 16212 28868 23492
rect 28924 23380 28980 23390
rect 29372 23380 29428 23884
rect 29484 23874 29540 23884
rect 29596 23940 29652 23950
rect 28980 23324 29428 23380
rect 28924 23286 28980 23324
rect 29484 23156 29540 23166
rect 29596 23156 29652 23884
rect 29484 23154 29652 23156
rect 29484 23102 29486 23154
rect 29538 23102 29652 23154
rect 29484 23100 29652 23102
rect 29484 23090 29540 23100
rect 29260 22932 29316 22942
rect 29260 22838 29316 22876
rect 29260 22372 29316 22382
rect 29036 22258 29092 22270
rect 29036 22206 29038 22258
rect 29090 22206 29092 22258
rect 29036 22148 29092 22206
rect 29036 22082 29092 22092
rect 29148 21476 29204 21486
rect 29148 20802 29204 21420
rect 29260 21364 29316 22316
rect 29372 22258 29428 22270
rect 29708 22260 29764 24108
rect 30156 24050 30212 25452
rect 30268 25396 30324 26852
rect 30716 26514 30772 27132
rect 30716 26462 30718 26514
rect 30770 26462 30772 26514
rect 30716 26450 30772 26462
rect 30828 26964 30884 26974
rect 30492 26292 30548 26302
rect 30548 26236 30660 26292
rect 30492 26226 30548 26236
rect 30492 26068 30548 26078
rect 30268 24500 30324 25340
rect 30268 24434 30324 24444
rect 30380 26012 30492 26068
rect 30156 23998 30158 24050
rect 30210 23998 30212 24050
rect 30156 23986 30212 23998
rect 29825 23548 30089 23558
rect 29881 23492 29929 23548
rect 29985 23492 30033 23548
rect 29825 23482 30089 23492
rect 30156 23156 30212 23166
rect 30156 22370 30212 23100
rect 30268 23044 30324 23054
rect 30268 22950 30324 22988
rect 30156 22318 30158 22370
rect 30210 22318 30212 22370
rect 30156 22306 30212 22318
rect 29372 22206 29374 22258
rect 29426 22206 29428 22258
rect 29372 21588 29428 22206
rect 29372 21522 29428 21532
rect 29596 22204 29764 22260
rect 29932 22258 29988 22270
rect 29932 22206 29934 22258
rect 29986 22206 29988 22258
rect 29596 21476 29652 22204
rect 29932 22148 29988 22206
rect 29596 21410 29652 21420
rect 29708 22092 29988 22148
rect 29708 21586 29764 22092
rect 29825 21980 30089 21990
rect 29881 21924 29929 21980
rect 29985 21924 30033 21980
rect 29825 21914 30089 21924
rect 29708 21534 29710 21586
rect 29762 21534 29764 21586
rect 29260 21308 29428 21364
rect 29148 20750 29150 20802
rect 29202 20750 29204 20802
rect 29148 20738 29204 20750
rect 29260 20692 29316 20702
rect 29260 20598 29316 20636
rect 29372 20018 29428 21308
rect 29708 20244 29764 21534
rect 30268 21588 30324 21598
rect 30268 21474 30324 21532
rect 30268 21422 30270 21474
rect 30322 21422 30324 21474
rect 30268 21410 30324 21422
rect 30380 21252 30436 26012
rect 30492 26002 30548 26012
rect 30604 25172 30660 26236
rect 30716 25508 30772 25518
rect 30828 25508 30884 26908
rect 30940 26908 30996 27132
rect 31164 27468 31444 27524
rect 30940 26852 31108 26908
rect 30940 26404 30996 26414
rect 30940 26310 30996 26348
rect 31052 26290 31108 26852
rect 31052 26238 31054 26290
rect 31106 26238 31108 26290
rect 31052 26226 31108 26238
rect 31164 25732 31220 27468
rect 31724 27186 31780 28476
rect 32172 27970 32228 27982
rect 32172 27918 32174 27970
rect 32226 27918 32228 27970
rect 32172 27748 32228 27918
rect 32172 27682 32228 27692
rect 32284 27746 32340 27758
rect 32284 27694 32286 27746
rect 32338 27694 32340 27746
rect 31724 27134 31726 27186
rect 31778 27134 31780 27186
rect 31724 27122 31780 27134
rect 31276 27074 31332 27086
rect 31276 27022 31278 27074
rect 31330 27022 31332 27074
rect 31276 26908 31332 27022
rect 32060 26964 32116 27002
rect 31276 26852 31556 26908
rect 32060 26898 32116 26908
rect 30772 25452 30884 25508
rect 31052 25676 31220 25732
rect 30716 25414 30772 25452
rect 30492 24836 30548 24846
rect 30492 24742 30548 24780
rect 30492 23828 30548 23838
rect 30604 23828 30660 25116
rect 30940 24724 30996 24734
rect 30492 23826 30660 23828
rect 30492 23774 30494 23826
rect 30546 23774 30660 23826
rect 30492 23772 30660 23774
rect 30716 24612 30772 24622
rect 30716 23938 30772 24556
rect 30940 24610 30996 24668
rect 30940 24558 30942 24610
rect 30994 24558 30996 24610
rect 30940 24546 30996 24558
rect 30716 23886 30718 23938
rect 30770 23886 30772 23938
rect 30492 23762 30548 23772
rect 30604 23380 30660 23390
rect 30492 23268 30548 23278
rect 30492 23174 30548 23212
rect 30604 22708 30660 23324
rect 30604 22642 30660 22652
rect 30604 22260 30660 22270
rect 30604 22166 30660 22204
rect 30268 21196 30436 21252
rect 30492 21476 30548 21486
rect 30268 21028 30324 21196
rect 30156 20972 30324 21028
rect 30156 20804 30212 20972
rect 30492 20916 30548 21420
rect 30716 20916 30772 23886
rect 30828 23156 30884 23166
rect 30828 23062 30884 23100
rect 30940 22596 30996 22606
rect 30828 22484 30884 22494
rect 30828 22370 30884 22428
rect 30828 22318 30830 22370
rect 30882 22318 30884 22370
rect 30828 22306 30884 22318
rect 30940 21588 30996 22540
rect 30716 20860 30884 20916
rect 29825 20412 30089 20422
rect 29881 20356 29929 20412
rect 29985 20356 30033 20412
rect 29825 20346 30089 20356
rect 30156 20244 30212 20748
rect 30268 20804 30324 20814
rect 30268 20802 30436 20804
rect 30268 20750 30270 20802
rect 30322 20750 30436 20802
rect 30268 20748 30436 20750
rect 30268 20738 30324 20748
rect 30380 20244 30436 20748
rect 30492 20802 30548 20860
rect 30492 20750 30494 20802
rect 30546 20750 30548 20802
rect 30492 20738 30548 20750
rect 30716 20692 30772 20702
rect 30604 20636 30716 20692
rect 30492 20244 30548 20254
rect 30156 20188 30324 20244
rect 30380 20242 30548 20244
rect 30380 20190 30494 20242
rect 30546 20190 30548 20242
rect 30380 20188 30548 20190
rect 29708 20178 29764 20188
rect 29372 19966 29374 20018
rect 29426 19966 29428 20018
rect 29372 19908 29428 19966
rect 30156 20020 30212 20030
rect 30156 19926 30212 19964
rect 29932 19908 29988 19918
rect 29372 19906 29988 19908
rect 29372 19854 29934 19906
rect 29986 19854 29988 19906
rect 29372 19852 29988 19854
rect 29932 19460 29988 19852
rect 29932 19394 29988 19404
rect 29260 19348 29316 19358
rect 29260 19254 29316 19292
rect 30268 19346 30324 20188
rect 30492 20178 30548 20188
rect 30604 20020 30660 20636
rect 30716 20626 30772 20636
rect 30268 19294 30270 19346
rect 30322 19294 30324 19346
rect 30268 19282 30324 19294
rect 30492 19964 30660 20020
rect 30716 20132 30772 20142
rect 29036 19236 29092 19246
rect 29036 19142 29092 19180
rect 29484 19124 29540 19134
rect 29484 19030 29540 19068
rect 29708 19122 29764 19134
rect 29708 19070 29710 19122
rect 29762 19070 29764 19122
rect 29708 18676 29764 19070
rect 30268 18900 30324 18910
rect 29825 18844 30089 18854
rect 29881 18788 29929 18844
rect 29985 18788 30033 18844
rect 29825 18778 30089 18788
rect 30156 18844 30268 18900
rect 30044 18676 30100 18686
rect 29708 18674 30100 18676
rect 29708 18622 30046 18674
rect 30098 18622 30100 18674
rect 29708 18620 30100 18622
rect 30044 18610 30100 18620
rect 29148 18450 29204 18462
rect 29148 18398 29150 18450
rect 29202 18398 29204 18450
rect 29148 17892 29204 18398
rect 29260 18452 29316 18462
rect 29260 18358 29316 18396
rect 29372 18452 29428 18462
rect 29820 18452 29876 18462
rect 29372 18450 29540 18452
rect 29372 18398 29374 18450
rect 29426 18398 29540 18450
rect 29372 18396 29540 18398
rect 29372 18386 29428 18396
rect 29148 17826 29204 17836
rect 29148 17668 29204 17678
rect 29148 17574 29204 17612
rect 29484 17444 29540 18396
rect 29820 18358 29876 18396
rect 30156 18116 30212 18844
rect 30268 18834 30324 18844
rect 30380 18340 30436 18350
rect 30380 18246 30436 18284
rect 30156 18050 30212 18060
rect 30044 17892 30100 17902
rect 30044 17780 30100 17836
rect 30044 17778 30212 17780
rect 30044 17726 30046 17778
rect 30098 17726 30212 17778
rect 30044 17724 30212 17726
rect 30044 17714 30100 17724
rect 29596 17666 29652 17678
rect 29596 17614 29598 17666
rect 29650 17614 29652 17666
rect 29596 17444 29652 17614
rect 29372 17388 29652 17444
rect 29036 16996 29092 17006
rect 29372 16996 29428 17388
rect 29825 17276 30089 17286
rect 29881 17220 29929 17276
rect 29985 17220 30033 17276
rect 29825 17210 30089 17220
rect 30156 17108 30212 17724
rect 30492 17220 30548 19964
rect 30604 19348 30660 19358
rect 30716 19348 30772 20076
rect 30604 19346 30772 19348
rect 30604 19294 30606 19346
rect 30658 19294 30772 19346
rect 30604 19292 30772 19294
rect 30604 19012 30660 19292
rect 30604 18946 30660 18956
rect 30716 18452 30772 18462
rect 30604 18338 30660 18350
rect 30604 18286 30606 18338
rect 30658 18286 30660 18338
rect 30604 18228 30660 18286
rect 30604 18162 30660 18172
rect 30716 17890 30772 18396
rect 30716 17838 30718 17890
rect 30770 17838 30772 17890
rect 30716 17826 30772 17838
rect 30828 17666 30884 20860
rect 30940 20244 30996 21532
rect 31052 20692 31108 25676
rect 31500 25620 31556 26852
rect 32172 26850 32228 26862
rect 32172 26798 32174 26850
rect 32226 26798 32228 26850
rect 31612 26292 31668 26302
rect 31612 26198 31668 26236
rect 32060 26292 32116 26302
rect 32060 25730 32116 26236
rect 32060 25678 32062 25730
rect 32114 25678 32116 25730
rect 32060 25666 32116 25678
rect 31612 25620 31668 25630
rect 31948 25620 32004 25630
rect 31500 25618 32004 25620
rect 31500 25566 31614 25618
rect 31666 25566 31950 25618
rect 32002 25566 32004 25618
rect 31500 25564 32004 25566
rect 31612 25554 31668 25564
rect 31948 25554 32004 25564
rect 31164 25508 31220 25518
rect 31164 25414 31220 25452
rect 32172 25508 32228 26798
rect 32284 26292 32340 27694
rect 32284 26226 32340 26236
rect 32396 26850 32452 26862
rect 32396 26798 32398 26850
rect 32450 26798 32452 26850
rect 32396 26290 32452 26798
rect 32396 26238 32398 26290
rect 32450 26238 32452 26290
rect 32396 26226 32452 26238
rect 32172 24948 32228 25452
rect 32732 25282 32788 28588
rect 32844 28578 32900 28588
rect 32956 28644 33012 28654
rect 32956 26908 33012 28588
rect 33068 28196 33124 29708
rect 33180 29428 33236 29438
rect 33180 28644 33236 29372
rect 33292 29316 33348 29326
rect 33292 29314 33460 29316
rect 33292 29262 33294 29314
rect 33346 29262 33460 29314
rect 33292 29260 33460 29262
rect 33292 29250 33348 29260
rect 33292 28756 33348 28766
rect 33292 28662 33348 28700
rect 33180 28550 33236 28588
rect 33404 28644 33460 29260
rect 33516 28756 33572 31948
rect 33852 31892 33908 31902
rect 33852 31798 33908 31836
rect 33740 31780 33796 31790
rect 33628 30210 33684 30222
rect 33628 30158 33630 30210
rect 33682 30158 33684 30210
rect 33628 29426 33684 30158
rect 33628 29374 33630 29426
rect 33682 29374 33684 29426
rect 33628 29204 33684 29374
rect 33740 29428 33796 31724
rect 34412 31444 34468 32286
rect 34860 31892 34916 32508
rect 34972 31892 35028 31902
rect 34860 31836 34972 31892
rect 34524 31778 34580 31790
rect 34524 31726 34526 31778
rect 34578 31726 34580 31778
rect 34524 31668 34580 31726
rect 34524 31602 34580 31612
rect 34748 31778 34804 31790
rect 34748 31726 34750 31778
rect 34802 31726 34804 31778
rect 34412 31378 34468 31388
rect 34748 31108 34804 31726
rect 34188 31106 34804 31108
rect 34188 31054 34750 31106
rect 34802 31054 34804 31106
rect 34188 31052 34804 31054
rect 34076 30996 34132 31006
rect 34076 30902 34132 30940
rect 34076 30324 34132 30334
rect 34188 30324 34244 31052
rect 34748 31042 34804 31052
rect 34412 30884 34468 30894
rect 34860 30884 34916 31836
rect 34972 31826 35028 31836
rect 34412 30882 34916 30884
rect 34412 30830 34414 30882
rect 34466 30830 34916 30882
rect 34412 30828 34916 30830
rect 34412 30818 34468 30828
rect 34076 30322 34244 30324
rect 34076 30270 34078 30322
rect 34130 30270 34244 30322
rect 34076 30268 34244 30270
rect 34076 30258 34132 30268
rect 34636 29652 34692 29662
rect 34524 29540 34580 29550
rect 34188 29538 34580 29540
rect 34188 29486 34526 29538
rect 34578 29486 34580 29538
rect 34188 29484 34580 29486
rect 33740 29372 34132 29428
rect 34076 29314 34132 29372
rect 34076 29262 34078 29314
rect 34130 29262 34132 29314
rect 34076 29250 34132 29262
rect 33740 29204 33796 29214
rect 33628 29148 33740 29204
rect 33740 29138 33796 29148
rect 34188 28980 34244 29484
rect 34524 29474 34580 29484
rect 34636 29538 34692 29596
rect 34636 29486 34638 29538
rect 34690 29486 34692 29538
rect 34636 29474 34692 29486
rect 34524 29204 34580 29214
rect 34524 29110 34580 29148
rect 33852 28924 34244 28980
rect 33852 28866 33908 28924
rect 33852 28814 33854 28866
rect 33906 28814 33908 28866
rect 33852 28802 33908 28814
rect 33516 28700 33684 28756
rect 33404 28642 33572 28644
rect 33404 28590 33406 28642
rect 33458 28590 33572 28642
rect 33404 28588 33572 28590
rect 33404 28578 33460 28588
rect 33068 28140 33460 28196
rect 33292 26962 33348 26974
rect 33292 26910 33294 26962
rect 33346 26910 33348 26962
rect 32844 26850 32900 26862
rect 32956 26852 33236 26908
rect 32844 26798 32846 26850
rect 32898 26798 32900 26850
rect 32844 25844 32900 26798
rect 33180 26628 33236 26852
rect 33180 26562 33236 26572
rect 33292 26516 33348 26910
rect 33292 26450 33348 26460
rect 33404 26514 33460 28140
rect 33404 26462 33406 26514
rect 33458 26462 33460 26514
rect 33404 26450 33460 26462
rect 33516 26514 33572 28588
rect 33628 28420 33684 28700
rect 33740 28644 33796 28654
rect 33740 28550 33796 28588
rect 33628 28364 33908 28420
rect 33740 27746 33796 27758
rect 33740 27694 33742 27746
rect 33794 27694 33796 27746
rect 33740 27076 33796 27694
rect 33740 27010 33796 27020
rect 33852 27186 33908 28364
rect 34524 28418 34580 28430
rect 34524 28366 34526 28418
rect 34578 28366 34580 28418
rect 34188 27860 34244 27870
rect 34188 27858 34356 27860
rect 34188 27806 34190 27858
rect 34242 27806 34356 27858
rect 34188 27804 34356 27806
rect 34188 27794 34244 27804
rect 33852 27134 33854 27186
rect 33906 27134 33908 27186
rect 33852 26908 33908 27134
rect 34076 27076 34132 27114
rect 34076 27010 34132 27020
rect 34300 27076 34356 27804
rect 34524 27636 34580 28366
rect 34636 27860 34692 27870
rect 34972 27860 35028 27870
rect 34636 27766 34692 27804
rect 34748 27858 35028 27860
rect 34748 27806 34974 27858
rect 35026 27806 35028 27858
rect 34748 27804 35028 27806
rect 34524 27570 34580 27580
rect 34748 27412 34804 27804
rect 34972 27794 35028 27804
rect 34412 27356 34804 27412
rect 34860 27412 34916 27422
rect 34412 27298 34468 27356
rect 34412 27246 34414 27298
rect 34466 27246 34468 27298
rect 34412 27234 34468 27246
rect 34636 27076 34692 27086
rect 34300 27074 34692 27076
rect 34300 27022 34638 27074
rect 34690 27022 34692 27074
rect 34300 27020 34692 27022
rect 34300 26962 34356 27020
rect 34636 27010 34692 27020
rect 34300 26910 34302 26962
rect 34354 26910 34356 26962
rect 33852 26852 34132 26908
rect 34300 26898 34356 26910
rect 34860 26962 34916 27356
rect 34860 26910 34862 26962
rect 34914 26910 34916 26962
rect 34860 26898 34916 26910
rect 34972 26964 35028 27002
rect 34972 26898 35028 26908
rect 34076 26740 34132 26852
rect 34076 26684 34468 26740
rect 33964 26628 34020 26638
rect 33516 26462 33518 26514
rect 33570 26462 33572 26514
rect 33516 26450 33572 26462
rect 33852 26516 33908 26526
rect 33180 26402 33236 26414
rect 33180 26350 33182 26402
rect 33234 26350 33236 26402
rect 32844 25778 32900 25788
rect 33068 26290 33124 26302
rect 33068 26238 33070 26290
rect 33122 26238 33124 26290
rect 33068 25620 33124 26238
rect 33180 26292 33236 26350
rect 33740 26404 33796 26414
rect 33740 26292 33796 26348
rect 33180 26236 33796 26292
rect 33852 26290 33908 26460
rect 33852 26238 33854 26290
rect 33906 26238 33908 26290
rect 33180 25844 33236 26236
rect 33180 25778 33236 25788
rect 33852 25620 33908 26238
rect 33964 25730 34020 26572
rect 34300 26404 34356 26414
rect 34300 26310 34356 26348
rect 34188 26292 34244 26302
rect 33964 25678 33966 25730
rect 34018 25678 34020 25730
rect 33964 25666 34020 25678
rect 34076 26290 34244 26292
rect 34076 26238 34190 26290
rect 34242 26238 34244 26290
rect 34076 26236 34244 26238
rect 33068 25564 33348 25620
rect 33292 25508 33348 25564
rect 33740 25564 33908 25620
rect 33516 25508 33572 25518
rect 33292 25506 33572 25508
rect 33292 25454 33518 25506
rect 33570 25454 33572 25506
rect 33292 25452 33572 25454
rect 32732 25230 32734 25282
rect 32786 25230 32788 25282
rect 32732 25218 32788 25230
rect 32956 25394 33012 25406
rect 32956 25342 32958 25394
rect 33010 25342 33012 25394
rect 32956 25284 33012 25342
rect 33180 25396 33236 25406
rect 33180 25302 33236 25340
rect 32956 25218 33012 25228
rect 32284 24948 32340 24958
rect 32172 24946 32340 24948
rect 32172 24894 32286 24946
rect 32338 24894 32340 24946
rect 32172 24892 32340 24894
rect 32284 24882 32340 24892
rect 31724 24722 31780 24734
rect 31724 24670 31726 24722
rect 31778 24670 31780 24722
rect 31500 24612 31556 24622
rect 31500 24518 31556 24556
rect 31724 23940 31780 24670
rect 32172 24724 32228 24734
rect 31724 23874 31780 23884
rect 31948 24276 32004 24286
rect 31388 23716 31444 23726
rect 31388 23378 31444 23660
rect 31388 23326 31390 23378
rect 31442 23326 31444 23378
rect 31388 23314 31444 23326
rect 31724 23380 31780 23390
rect 31164 23268 31220 23278
rect 31500 23268 31556 23278
rect 31164 23266 31332 23268
rect 31164 23214 31166 23266
rect 31218 23214 31332 23266
rect 31164 23212 31332 23214
rect 31164 23202 31220 23212
rect 31164 22932 31220 22942
rect 31164 22370 31220 22876
rect 31164 22318 31166 22370
rect 31218 22318 31220 22370
rect 31164 22306 31220 22318
rect 31276 22708 31332 23212
rect 31164 21252 31220 21262
rect 31276 21252 31332 22652
rect 31500 22484 31556 23212
rect 31612 23266 31668 23278
rect 31612 23214 31614 23266
rect 31666 23214 31668 23266
rect 31612 22932 31668 23214
rect 31724 23266 31780 23324
rect 31724 23214 31726 23266
rect 31778 23214 31780 23266
rect 31724 23202 31780 23214
rect 31612 22866 31668 22876
rect 31836 23044 31892 23054
rect 31500 22428 31668 22484
rect 31388 22260 31444 22270
rect 31388 22166 31444 22204
rect 31500 22258 31556 22270
rect 31500 22206 31502 22258
rect 31554 22206 31556 22258
rect 31500 21588 31556 22206
rect 31612 22036 31668 22428
rect 31612 21810 31668 21980
rect 31612 21758 31614 21810
rect 31666 21758 31668 21810
rect 31612 21746 31668 21758
rect 31500 21522 31556 21532
rect 31220 21196 31332 21252
rect 31164 21186 31220 21196
rect 31836 20802 31892 22988
rect 31948 22484 32004 24220
rect 32060 23938 32116 23950
rect 32060 23886 32062 23938
rect 32114 23886 32116 23938
rect 32060 23828 32116 23886
rect 32060 22932 32116 23772
rect 32172 23378 32228 24668
rect 32396 24724 32452 24734
rect 33180 24724 33236 24734
rect 32396 24722 33236 24724
rect 32396 24670 32398 24722
rect 32450 24670 33182 24722
rect 33234 24670 33236 24722
rect 32396 24668 33236 24670
rect 32396 24658 32452 24668
rect 32508 24162 32564 24668
rect 33180 24658 33236 24668
rect 33404 24724 33460 24734
rect 33404 24630 33460 24668
rect 32508 24110 32510 24162
rect 32562 24110 32564 24162
rect 32508 24098 32564 24110
rect 33516 24052 33572 25452
rect 33404 23996 33572 24052
rect 33628 24948 33684 24958
rect 33628 24050 33684 24892
rect 33628 23998 33630 24050
rect 33682 23998 33684 24050
rect 32396 23940 32452 23950
rect 32396 23846 32452 23884
rect 32956 23940 33012 23950
rect 32956 23846 33012 23884
rect 33068 23828 33124 23838
rect 33068 23734 33124 23772
rect 32172 23326 32174 23378
rect 32226 23326 32228 23378
rect 32172 23314 32228 23326
rect 32284 23716 32340 23726
rect 32284 23380 32340 23660
rect 33292 23492 33348 23502
rect 32396 23380 32452 23390
rect 32284 23378 32452 23380
rect 32284 23326 32398 23378
rect 32450 23326 32452 23378
rect 32284 23324 32452 23326
rect 32060 22866 32116 22876
rect 31948 22418 32004 22428
rect 32060 22258 32116 22270
rect 32060 22206 32062 22258
rect 32114 22206 32116 22258
rect 31948 22148 32004 22158
rect 32060 22148 32116 22206
rect 32004 22092 32116 22148
rect 32284 22146 32340 23324
rect 32396 23314 32452 23324
rect 33292 23378 33348 23436
rect 33292 23326 33294 23378
rect 33346 23326 33348 23378
rect 33292 23314 33348 23326
rect 32508 23156 32564 23166
rect 32956 23156 33012 23166
rect 32508 23154 32788 23156
rect 32508 23102 32510 23154
rect 32562 23102 32788 23154
rect 32508 23100 32788 23102
rect 32508 23090 32564 23100
rect 32508 22484 32564 22494
rect 32284 22094 32286 22146
rect 32338 22094 32340 22146
rect 31948 22082 32004 22092
rect 32284 22082 32340 22094
rect 32396 22372 32452 22382
rect 32396 21810 32452 22316
rect 32508 22260 32564 22428
rect 32620 22260 32676 22270
rect 32508 22258 32676 22260
rect 32508 22206 32622 22258
rect 32674 22206 32676 22258
rect 32508 22204 32676 22206
rect 32620 22148 32676 22204
rect 32620 22082 32676 22092
rect 32396 21758 32398 21810
rect 32450 21758 32452 21810
rect 32396 21746 32452 21758
rect 32508 21812 32564 21822
rect 31948 21588 32004 21598
rect 31948 21494 32004 21532
rect 32172 21586 32228 21598
rect 32172 21534 32174 21586
rect 32226 21534 32228 21586
rect 32060 21476 32116 21486
rect 32060 20914 32116 21420
rect 32172 21140 32228 21534
rect 32508 21586 32564 21756
rect 32508 21534 32510 21586
rect 32562 21534 32564 21586
rect 32508 21476 32564 21534
rect 32508 21410 32564 21420
rect 32620 21588 32676 21598
rect 32732 21588 32788 23100
rect 32844 23154 33012 23156
rect 32844 23102 32958 23154
rect 33010 23102 33012 23154
rect 32844 23100 33012 23102
rect 32844 22370 32900 23100
rect 32956 23090 33012 23100
rect 33180 22932 33236 22942
rect 32844 22318 32846 22370
rect 32898 22318 32900 22370
rect 32844 21812 32900 22318
rect 32844 21746 32900 21756
rect 32956 22930 33236 22932
rect 32956 22878 33182 22930
rect 33234 22878 33236 22930
rect 32956 22876 33236 22878
rect 32844 21588 32900 21598
rect 32732 21532 32844 21588
rect 32956 21588 33012 22876
rect 33180 22866 33236 22876
rect 33292 22708 33348 22718
rect 33404 22708 33460 23996
rect 33628 23986 33684 23998
rect 33740 23492 33796 25564
rect 34076 25508 34132 26236
rect 34188 26226 34244 26236
rect 33852 25452 34132 25508
rect 34188 25506 34244 25518
rect 34188 25454 34190 25506
rect 34242 25454 34244 25506
rect 33852 25172 33908 25452
rect 33852 25106 33908 25116
rect 34076 25060 34132 25070
rect 34076 24834 34132 25004
rect 34076 24782 34078 24834
rect 34130 24782 34132 24834
rect 34076 24770 34132 24782
rect 34076 23938 34132 23950
rect 34076 23886 34078 23938
rect 34130 23886 34132 23938
rect 33852 23492 33908 23502
rect 34076 23492 34132 23886
rect 34188 23548 34244 25454
rect 34412 25284 34468 26684
rect 34524 26516 34580 26526
rect 34524 26422 34580 26460
rect 34860 26404 34916 26414
rect 34860 26310 34916 26348
rect 34972 26292 35028 26302
rect 34972 25618 35028 26236
rect 34972 25566 34974 25618
rect 35026 25566 35028 25618
rect 34412 24610 34468 25228
rect 34860 25508 34916 25518
rect 34860 24722 34916 25452
rect 34972 25396 35028 25566
rect 34972 25330 35028 25340
rect 34860 24670 34862 24722
rect 34914 24670 34916 24722
rect 34860 24658 34916 24670
rect 34412 24558 34414 24610
rect 34466 24558 34468 24610
rect 34188 23492 34356 23548
rect 33740 23436 33852 23492
rect 33908 23436 34020 23492
rect 33852 23426 33908 23436
rect 33348 22652 33460 22708
rect 33516 23380 33572 23390
rect 33516 23266 33572 23324
rect 33964 23378 34020 23436
rect 34076 23426 34132 23436
rect 33964 23326 33966 23378
rect 34018 23326 34020 23378
rect 33964 23314 34020 23326
rect 33516 23214 33518 23266
rect 33570 23214 33572 23266
rect 33292 22642 33348 22652
rect 33404 22372 33460 22382
rect 33404 22278 33460 22316
rect 33292 22258 33348 22270
rect 33292 22206 33294 22258
rect 33346 22206 33348 22258
rect 33292 21924 33348 22206
rect 33292 21868 33460 21924
rect 33068 21588 33124 21598
rect 32956 21586 33124 21588
rect 32956 21534 33070 21586
rect 33122 21534 33124 21586
rect 32956 21532 33124 21534
rect 32172 21074 32228 21084
rect 32060 20862 32062 20914
rect 32114 20862 32116 20914
rect 32060 20850 32116 20862
rect 32620 20914 32676 21532
rect 32844 21522 32900 21532
rect 33068 21522 33124 21532
rect 33404 21586 33460 21868
rect 33516 21812 33572 23214
rect 34300 23156 34356 23492
rect 34300 23062 34356 23100
rect 34412 22932 34468 24558
rect 34636 23714 34692 23726
rect 34636 23662 34638 23714
rect 34690 23662 34692 23714
rect 34636 23380 34692 23662
rect 34636 23314 34692 23324
rect 34860 23268 34916 23278
rect 34860 23174 34916 23212
rect 34300 22876 34468 22932
rect 33964 22370 34020 22382
rect 33964 22318 33966 22370
rect 34018 22318 34020 22370
rect 33964 22260 34020 22318
rect 33516 21746 33572 21756
rect 33628 22204 33964 22260
rect 33628 21810 33684 22204
rect 33964 22194 34020 22204
rect 33628 21758 33630 21810
rect 33682 21758 33684 21810
rect 33628 21746 33684 21758
rect 33740 21924 33796 21934
rect 33404 21534 33406 21586
rect 33458 21534 33460 21586
rect 33404 21522 33460 21534
rect 33628 21588 33684 21598
rect 33628 21474 33684 21532
rect 33628 21422 33630 21474
rect 33682 21422 33684 21474
rect 33628 21410 33684 21422
rect 32620 20862 32622 20914
rect 32674 20862 32676 20914
rect 32620 20850 32676 20862
rect 33180 21252 33236 21262
rect 33740 21252 33796 21868
rect 33852 21812 33908 21822
rect 33852 21718 33908 21756
rect 31836 20750 31838 20802
rect 31890 20750 31892 20802
rect 31836 20738 31892 20750
rect 32732 20804 32788 20814
rect 32732 20710 32788 20748
rect 33180 20802 33236 21196
rect 33180 20750 33182 20802
rect 33234 20750 33236 20802
rect 33180 20738 33236 20750
rect 33516 21196 33796 21252
rect 33516 20804 33572 21196
rect 33516 20710 33572 20748
rect 33852 21140 33908 21150
rect 33852 20914 33908 21084
rect 33852 20862 33854 20914
rect 33906 20862 33908 20914
rect 31052 20626 31108 20636
rect 32172 20692 32228 20702
rect 32172 20598 32228 20636
rect 33852 20692 33908 20862
rect 33852 20626 33908 20636
rect 32508 20580 32564 20590
rect 31052 20244 31108 20254
rect 30940 20242 31108 20244
rect 30940 20190 31054 20242
rect 31106 20190 31108 20242
rect 30940 20188 31108 20190
rect 31052 20178 31108 20188
rect 31388 20244 31444 20254
rect 31388 20130 31444 20188
rect 31388 20078 31390 20130
rect 31442 20078 31444 20130
rect 31388 20066 31444 20078
rect 32508 20132 32564 20524
rect 32508 20066 32564 20076
rect 31948 20020 32004 20030
rect 31836 19964 31948 20020
rect 30940 19404 31444 19460
rect 30940 18562 30996 19404
rect 31388 19348 31444 19404
rect 31500 19348 31556 19358
rect 31388 19346 31556 19348
rect 31388 19294 31502 19346
rect 31554 19294 31556 19346
rect 31388 19292 31556 19294
rect 31836 19348 31892 19964
rect 31948 19954 32004 19964
rect 33180 20020 33236 20030
rect 33180 19926 33236 19964
rect 32508 19906 32564 19918
rect 32508 19854 32510 19906
rect 32562 19854 32564 19906
rect 31948 19794 32004 19806
rect 31948 19742 31950 19794
rect 32002 19742 32004 19794
rect 31948 19572 32004 19742
rect 32284 19796 32340 19806
rect 32284 19702 32340 19740
rect 32508 19684 32564 19854
rect 33068 19796 33124 19806
rect 32732 19684 32788 19694
rect 32508 19628 32732 19684
rect 32732 19618 32788 19628
rect 31948 19506 32004 19516
rect 32844 19572 32900 19582
rect 32732 19460 32788 19470
rect 32732 19366 32788 19404
rect 31948 19348 32004 19358
rect 31836 19346 32004 19348
rect 31836 19294 31950 19346
rect 32002 19294 32004 19346
rect 31836 19292 32004 19294
rect 31276 19236 31332 19246
rect 30940 18510 30942 18562
rect 30994 18510 30996 18562
rect 30940 18498 30996 18510
rect 31052 19234 31332 19236
rect 31052 19182 31278 19234
rect 31330 19182 31332 19234
rect 31052 19180 31332 19182
rect 31052 18562 31108 19180
rect 31276 19170 31332 19180
rect 31052 18510 31054 18562
rect 31106 18510 31108 18562
rect 31052 17892 31108 18510
rect 31500 18562 31556 19292
rect 31948 19282 32004 19292
rect 32844 19346 32900 19516
rect 33068 19460 33124 19740
rect 33068 19394 33124 19404
rect 34076 19348 34132 19358
rect 32844 19294 32846 19346
rect 32898 19294 32900 19346
rect 32844 19282 32900 19294
rect 33852 19346 34132 19348
rect 33852 19294 34078 19346
rect 34130 19294 34132 19346
rect 33852 19292 34132 19294
rect 33068 19236 33124 19246
rect 33068 19142 33124 19180
rect 33852 19234 33908 19292
rect 34076 19282 34132 19292
rect 33852 19182 33854 19234
rect 33906 19182 33908 19234
rect 33852 19170 33908 19182
rect 33180 19124 33236 19134
rect 32284 18676 32340 18686
rect 31500 18510 31502 18562
rect 31554 18510 31556 18562
rect 31500 18498 31556 18510
rect 32172 18620 32284 18676
rect 31276 18452 31332 18462
rect 31276 18450 31444 18452
rect 31276 18398 31278 18450
rect 31330 18398 31444 18450
rect 31276 18396 31444 18398
rect 31276 18386 31332 18396
rect 30828 17614 30830 17666
rect 30882 17614 30884 17666
rect 30604 17556 30660 17566
rect 30604 17554 30772 17556
rect 30604 17502 30606 17554
rect 30658 17502 30772 17554
rect 30604 17500 30772 17502
rect 30604 17490 30660 17500
rect 30380 17164 30548 17220
rect 30604 17220 30660 17230
rect 30268 17108 30324 17118
rect 30156 17106 30324 17108
rect 30156 17054 30270 17106
rect 30322 17054 30324 17106
rect 30156 17052 30324 17054
rect 30268 17042 30324 17052
rect 29036 16994 29428 16996
rect 29036 16942 29038 16994
rect 29090 16942 29428 16994
rect 29036 16940 29428 16942
rect 29036 16930 29092 16940
rect 29484 16884 29540 16894
rect 29372 16436 29428 16446
rect 29372 16212 29428 16380
rect 28700 15540 28756 15550
rect 28812 15540 28868 16156
rect 28700 15538 28868 15540
rect 28700 15486 28702 15538
rect 28754 15486 28868 15538
rect 28700 15484 28868 15486
rect 28924 16210 29428 16212
rect 28924 16158 29374 16210
rect 29426 16158 29428 16210
rect 28924 16156 29428 16158
rect 28924 15538 28980 16156
rect 29372 16146 29428 16156
rect 28924 15486 28926 15538
rect 28978 15486 28980 15538
rect 28700 15474 28756 15484
rect 28924 15474 28980 15486
rect 28476 15262 28478 15314
rect 28530 15262 28532 15314
rect 28252 14478 28254 14530
rect 28306 14478 28308 14530
rect 28252 14466 28308 14478
rect 28476 14420 28532 15262
rect 29372 15316 29428 15326
rect 29372 15222 29428 15260
rect 29484 15148 29540 16828
rect 29932 16772 29988 16782
rect 30380 16772 30436 17164
rect 30492 16996 30548 17006
rect 30492 16902 30548 16940
rect 30604 16994 30660 17164
rect 30604 16942 30606 16994
rect 30658 16942 30660 16994
rect 30604 16930 30660 16942
rect 30716 16884 30772 17500
rect 30828 17332 30884 17614
rect 30828 17266 30884 17276
rect 30940 17836 31108 17892
rect 31276 18228 31332 18238
rect 30716 16818 30772 16828
rect 30380 16716 30548 16772
rect 29932 16678 29988 16716
rect 30044 16324 30100 16334
rect 29708 16100 29764 16110
rect 29708 16006 29764 16044
rect 30044 16098 30100 16268
rect 30044 16046 30046 16098
rect 30098 16046 30100 16098
rect 30044 16034 30100 16046
rect 30380 16100 30436 16110
rect 29820 15876 29876 15914
rect 29820 15810 29876 15820
rect 29825 15708 30089 15718
rect 29881 15652 29929 15708
rect 29985 15652 30033 15708
rect 29825 15642 30089 15652
rect 29596 15428 29652 15438
rect 29596 15314 29652 15372
rect 30268 15428 30324 15438
rect 30380 15428 30436 16044
rect 30268 15426 30436 15428
rect 30268 15374 30270 15426
rect 30322 15374 30436 15426
rect 30268 15372 30436 15374
rect 30268 15362 30324 15372
rect 29596 15262 29598 15314
rect 29650 15262 29652 15314
rect 29596 15250 29652 15262
rect 28588 15090 28644 15102
rect 28588 15038 28590 15090
rect 28642 15038 28644 15090
rect 28588 14868 28644 15038
rect 28588 14802 28644 14812
rect 29036 15092 29540 15148
rect 28476 14354 28532 14364
rect 28252 14308 28308 14318
rect 28252 12402 28308 14252
rect 28252 12350 28254 12402
rect 28306 12350 28308 12402
rect 28252 12338 28308 12350
rect 28364 14306 28420 14318
rect 28364 14254 28366 14306
rect 28418 14254 28420 14306
rect 28252 12180 28308 12190
rect 28252 12086 28308 12124
rect 28364 12068 28420 14254
rect 28588 14308 28644 14318
rect 28588 13746 28644 14252
rect 28588 13694 28590 13746
rect 28642 13694 28644 13746
rect 28588 13682 28644 13694
rect 29036 12740 29092 15092
rect 29372 14530 29428 14542
rect 29372 14478 29374 14530
rect 29426 14478 29428 14530
rect 29148 14418 29204 14430
rect 29148 14366 29150 14418
rect 29202 14366 29204 14418
rect 29148 13972 29204 14366
rect 29148 13906 29204 13916
rect 29260 14306 29316 14318
rect 29260 14254 29262 14306
rect 29314 14254 29316 14306
rect 29148 12964 29204 12974
rect 29260 12964 29316 14254
rect 29372 13860 29428 14478
rect 30492 14532 30548 16716
rect 30716 16212 30772 16222
rect 30940 16212 30996 17836
rect 31276 17666 31332 18172
rect 31276 17614 31278 17666
rect 31330 17614 31332 17666
rect 31276 17602 31332 17614
rect 31388 17668 31444 18396
rect 32172 18450 32228 18620
rect 32172 18398 32174 18450
rect 32226 18398 32228 18450
rect 32172 18386 32228 18398
rect 32284 17778 32340 18620
rect 32396 18452 32452 18462
rect 32396 18358 32452 18396
rect 33068 18452 33124 18462
rect 33068 18358 33124 18396
rect 33180 18450 33236 19068
rect 34188 18788 34244 18798
rect 33292 18676 33348 18686
rect 33964 18676 34020 18686
rect 34188 18676 34244 18732
rect 33292 18582 33348 18620
rect 33404 18674 34020 18676
rect 33404 18622 33966 18674
rect 34018 18622 34020 18674
rect 33404 18620 34020 18622
rect 33180 18398 33182 18450
rect 33234 18398 33236 18450
rect 33180 18386 33236 18398
rect 33404 18228 33460 18620
rect 33964 18610 34020 18620
rect 34076 18674 34244 18676
rect 34076 18622 34190 18674
rect 34242 18622 34244 18674
rect 34076 18620 34244 18622
rect 33628 18452 33684 18462
rect 33852 18452 33908 18462
rect 33628 18450 33908 18452
rect 33628 18398 33630 18450
rect 33682 18398 33854 18450
rect 33906 18398 33908 18450
rect 33628 18396 33908 18398
rect 33628 18386 33684 18396
rect 33852 18386 33908 18396
rect 32284 17726 32286 17778
rect 32338 17726 32340 17778
rect 32284 17714 32340 17726
rect 33068 18172 33460 18228
rect 31612 17668 31668 17678
rect 31388 17666 31668 17668
rect 31388 17614 31614 17666
rect 31666 17614 31668 17666
rect 31388 17612 31668 17614
rect 31612 17602 31668 17612
rect 32732 17668 32788 17678
rect 31052 17444 31108 17454
rect 31052 17350 31108 17388
rect 31500 17442 31556 17454
rect 31500 17390 31502 17442
rect 31554 17390 31556 17442
rect 31388 17332 31444 17342
rect 31388 17106 31444 17276
rect 31388 17054 31390 17106
rect 31442 17054 31444 17106
rect 31388 17042 31444 17054
rect 31500 16324 31556 17390
rect 31724 17332 31780 17342
rect 31724 16996 31780 17276
rect 32172 17220 32228 17230
rect 32172 17106 32228 17164
rect 32172 17054 32174 17106
rect 32226 17054 32228 17106
rect 32172 17042 32228 17054
rect 31724 16902 31780 16940
rect 32396 16884 32452 16894
rect 31500 16258 31556 16268
rect 32284 16772 32340 16782
rect 31276 16212 31332 16222
rect 30940 16210 31332 16212
rect 30940 16158 31278 16210
rect 31330 16158 31332 16210
rect 30940 16156 31332 16158
rect 30716 15538 30772 16156
rect 31276 16146 31332 16156
rect 30716 15486 30718 15538
rect 30770 15486 30772 15538
rect 30716 15428 30772 15486
rect 30716 15362 30772 15372
rect 30828 16098 30884 16110
rect 30828 16046 30830 16098
rect 30882 16046 30884 16098
rect 30828 15876 30884 16046
rect 32284 16098 32340 16716
rect 32284 16046 32286 16098
rect 32338 16046 32340 16098
rect 32284 16034 32340 16046
rect 31724 15988 31780 15998
rect 31724 15894 31780 15932
rect 32060 15988 32116 15998
rect 32060 15894 32116 15932
rect 30828 15148 30884 15820
rect 31948 15876 32004 15886
rect 31948 15782 32004 15820
rect 32284 15652 32340 15662
rect 32284 15540 32340 15596
rect 32060 15484 32340 15540
rect 31276 15428 31332 15438
rect 31276 15148 31332 15372
rect 30828 15092 31108 15148
rect 31276 15092 31892 15148
rect 30492 14466 30548 14476
rect 29708 14418 29764 14430
rect 29708 14366 29710 14418
rect 29762 14366 29764 14418
rect 29372 13794 29428 13804
rect 29484 13858 29540 13870
rect 29484 13806 29486 13858
rect 29538 13806 29540 13858
rect 29148 12962 29316 12964
rect 29148 12910 29150 12962
rect 29202 12910 29316 12962
rect 29148 12908 29316 12910
rect 29372 12964 29428 12974
rect 29484 12964 29540 13806
rect 29708 13636 29764 14366
rect 30268 14418 30324 14430
rect 30268 14366 30270 14418
rect 30322 14366 30324 14418
rect 29932 14308 29988 14346
rect 29932 14242 29988 14252
rect 30156 14306 30212 14318
rect 30156 14254 30158 14306
rect 30210 14254 30212 14306
rect 29825 14140 30089 14150
rect 29881 14084 29929 14140
rect 29985 14084 30033 14140
rect 29825 14074 30089 14084
rect 30156 13860 30212 14254
rect 30268 13972 30324 14366
rect 30268 13906 30324 13916
rect 30716 13972 30772 13982
rect 30716 13878 30772 13916
rect 30156 13794 30212 13804
rect 30940 13860 30996 13870
rect 30492 13746 30548 13758
rect 30492 13694 30494 13746
rect 30546 13694 30548 13746
rect 30044 13636 30100 13646
rect 30492 13636 30548 13694
rect 29708 13634 30548 13636
rect 29708 13582 30046 13634
rect 30098 13582 30548 13634
rect 29708 13580 30548 13582
rect 30044 13570 30100 13580
rect 30380 13412 30436 13422
rect 30268 13356 30380 13412
rect 30156 13188 30212 13198
rect 29932 12964 29988 12974
rect 29372 12962 29988 12964
rect 29372 12910 29374 12962
rect 29426 12910 29934 12962
rect 29986 12910 29988 12962
rect 29372 12908 29988 12910
rect 29148 12898 29204 12908
rect 29372 12898 29428 12908
rect 29932 12898 29988 12908
rect 30156 12850 30212 13132
rect 30268 12964 30324 13356
rect 30380 13346 30436 13356
rect 30268 12962 30436 12964
rect 30268 12910 30270 12962
rect 30322 12910 30436 12962
rect 30268 12908 30436 12910
rect 30268 12898 30324 12908
rect 30156 12798 30158 12850
rect 30210 12798 30212 12850
rect 30156 12786 30212 12798
rect 29260 12740 29316 12750
rect 29036 12738 29316 12740
rect 29036 12686 29262 12738
rect 29314 12686 29316 12738
rect 29036 12684 29316 12686
rect 29260 12674 29316 12684
rect 29596 12740 29652 12750
rect 29596 12646 29652 12684
rect 29372 12628 29428 12638
rect 28924 12404 28980 12414
rect 28924 12310 28980 12348
rect 28364 12002 28420 12012
rect 28476 12178 28532 12190
rect 28476 12126 28478 12178
rect 28530 12126 28532 12178
rect 28476 11620 28532 12126
rect 28588 11620 28644 11630
rect 28476 11564 28588 11620
rect 28588 11554 28644 11564
rect 28140 10612 28196 11340
rect 28476 11284 28532 11294
rect 28140 10500 28196 10556
rect 28364 11172 28420 11182
rect 28252 10500 28308 10510
rect 28140 10498 28308 10500
rect 28140 10446 28254 10498
rect 28306 10446 28308 10498
rect 28140 10444 28308 10446
rect 28252 10434 28308 10444
rect 28364 10164 28420 11116
rect 28476 10276 28532 11228
rect 29372 10836 29428 12572
rect 29825 12572 30089 12582
rect 29881 12516 29929 12572
rect 29985 12516 30033 12572
rect 29825 12506 30089 12516
rect 29932 12292 29988 12302
rect 29932 12290 30324 12292
rect 29932 12238 29934 12290
rect 29986 12238 30324 12290
rect 29932 12236 30324 12238
rect 29932 12226 29988 12236
rect 29484 12180 29540 12190
rect 29484 11172 29540 12124
rect 29820 11620 29876 11630
rect 29596 11508 29652 11518
rect 29596 11394 29652 11452
rect 29596 11342 29598 11394
rect 29650 11342 29652 11394
rect 29596 11330 29652 11342
rect 29820 11394 29876 11564
rect 30268 11618 30324 12236
rect 30380 11732 30436 12908
rect 30492 12516 30548 13580
rect 30940 13636 30996 13804
rect 30940 13570 30996 13580
rect 30604 13522 30660 13534
rect 30604 13470 30606 13522
rect 30658 13470 30660 13522
rect 30604 12740 30660 13470
rect 31052 13074 31108 15092
rect 31724 14418 31780 14430
rect 31724 14366 31726 14418
rect 31778 14366 31780 14418
rect 31612 14308 31668 14318
rect 31500 13860 31556 13870
rect 31388 13858 31556 13860
rect 31388 13806 31502 13858
rect 31554 13806 31556 13858
rect 31388 13804 31556 13806
rect 31388 13188 31444 13804
rect 31500 13794 31556 13804
rect 31612 13746 31668 14252
rect 31612 13694 31614 13746
rect 31666 13694 31668 13746
rect 31500 13524 31556 13534
rect 31500 13430 31556 13468
rect 31388 13122 31444 13132
rect 31052 13022 31054 13074
rect 31106 13022 31108 13074
rect 31052 13010 31108 13022
rect 31164 12964 31220 12974
rect 31220 12908 31332 12964
rect 31164 12870 31220 12908
rect 30940 12852 30996 12862
rect 30940 12758 30996 12796
rect 30604 12674 30660 12684
rect 30716 12738 30772 12750
rect 30716 12686 30718 12738
rect 30770 12686 30772 12738
rect 30492 12460 30660 12516
rect 30380 11676 30548 11732
rect 30268 11566 30270 11618
rect 30322 11566 30324 11618
rect 30268 11554 30324 11566
rect 29820 11342 29822 11394
rect 29874 11342 29876 11394
rect 29820 11330 29876 11342
rect 30380 11508 30436 11518
rect 29708 11284 29764 11294
rect 29708 11190 29764 11228
rect 29484 11060 29540 11116
rect 30380 11060 30436 11452
rect 29484 11004 29652 11060
rect 29372 10770 29428 10780
rect 28812 10610 28868 10622
rect 28812 10558 28814 10610
rect 28866 10558 28868 10610
rect 28700 10388 28756 10398
rect 28476 10210 28532 10220
rect 28588 10386 28756 10388
rect 28588 10334 28702 10386
rect 28754 10334 28756 10386
rect 28588 10332 28756 10334
rect 28364 10098 28420 10108
rect 27580 9212 27860 9268
rect 27804 9156 27860 9212
rect 28028 9202 28084 9212
rect 28252 9826 28308 9838
rect 28252 9774 28254 9826
rect 28306 9774 28308 9826
rect 27692 9042 27748 9054
rect 27692 8990 27694 9042
rect 27746 8990 27748 9042
rect 27580 8932 27636 8942
rect 27580 8820 27636 8876
rect 27356 8818 27636 8820
rect 27356 8766 27358 8818
rect 27410 8766 27636 8818
rect 27356 8764 27636 8766
rect 27356 8754 27412 8764
rect 27020 7700 27076 7710
rect 26684 6962 26740 6972
rect 26796 7474 26852 7486
rect 26796 7422 26798 7474
rect 26850 7422 26852 7474
rect 26572 5854 26574 5906
rect 26626 5854 26628 5906
rect 26572 5842 26628 5854
rect 26684 6690 26740 6702
rect 26684 6638 26686 6690
rect 26738 6638 26740 6690
rect 26684 6356 26740 6638
rect 26348 5630 26350 5682
rect 26402 5630 26404 5682
rect 26348 5348 26404 5630
rect 26348 5282 26404 5292
rect 26236 4286 26238 4338
rect 26290 4286 26292 4338
rect 26236 4274 26292 4286
rect 26572 5012 26628 5022
rect 26572 4338 26628 4956
rect 26572 4286 26574 4338
rect 26626 4286 26628 4338
rect 26572 4228 26628 4286
rect 26572 4162 26628 4172
rect 26684 4226 26740 6300
rect 26796 5346 26852 7422
rect 27020 7474 27076 7644
rect 27020 7422 27022 7474
rect 27074 7422 27076 7474
rect 27020 7410 27076 7422
rect 27244 6130 27300 8204
rect 27580 8258 27636 8764
rect 27692 8596 27748 8990
rect 27804 8708 27860 9100
rect 28028 9044 28084 9054
rect 28252 9044 28308 9774
rect 28588 9044 28644 10332
rect 28700 10322 28756 10332
rect 28812 9268 28868 10558
rect 29596 10050 29652 11004
rect 29825 11004 30089 11014
rect 29881 10948 29929 11004
rect 29985 10948 30033 11004
rect 30380 10994 30436 11004
rect 29825 10938 30089 10948
rect 29596 9998 29598 10050
rect 29650 9998 29652 10050
rect 29596 9986 29652 9998
rect 29708 10612 29764 10622
rect 29708 9826 29764 10556
rect 29820 10498 29876 10510
rect 29820 10446 29822 10498
rect 29874 10446 29876 10498
rect 29820 10276 29876 10446
rect 29820 9938 29876 10220
rect 29820 9886 29822 9938
rect 29874 9886 29876 9938
rect 29820 9874 29876 9886
rect 29708 9774 29710 9826
rect 29762 9774 29764 9826
rect 29708 9762 29764 9774
rect 28812 9202 28868 9212
rect 29372 9604 29428 9614
rect 29372 9266 29428 9548
rect 29825 9436 30089 9446
rect 29881 9380 29929 9436
rect 29985 9380 30033 9436
rect 30492 9380 30548 11676
rect 29825 9370 30089 9380
rect 30380 9324 30548 9380
rect 29372 9214 29374 9266
rect 29426 9214 29428 9266
rect 29372 9202 29428 9214
rect 30044 9268 30100 9278
rect 28028 9042 28196 9044
rect 28028 8990 28030 9042
rect 28082 8990 28196 9042
rect 28028 8988 28196 8990
rect 28252 9042 28644 9044
rect 28252 8990 28590 9042
rect 28642 8990 28644 9042
rect 28252 8988 28644 8990
rect 28028 8978 28084 8988
rect 27804 8642 27860 8652
rect 27916 8930 27972 8942
rect 27916 8878 27918 8930
rect 27970 8878 27972 8930
rect 27692 8530 27748 8540
rect 27580 8206 27582 8258
rect 27634 8206 27636 8258
rect 27580 8194 27636 8206
rect 27804 8484 27860 8494
rect 27916 8484 27972 8878
rect 28140 8484 28196 8988
rect 27916 8428 28084 8484
rect 27804 8260 27860 8428
rect 27916 8260 27972 8270
rect 27804 8258 27972 8260
rect 27804 8206 27918 8258
rect 27970 8206 27972 8258
rect 27804 8204 27972 8206
rect 27692 7924 27748 7934
rect 27356 6692 27412 6702
rect 27356 6578 27412 6636
rect 27356 6526 27358 6578
rect 27410 6526 27412 6578
rect 27356 6514 27412 6526
rect 27244 6078 27246 6130
rect 27298 6078 27300 6130
rect 27244 6066 27300 6078
rect 27580 6468 27636 6478
rect 27468 5908 27524 5918
rect 27468 5572 27524 5852
rect 27468 5506 27524 5516
rect 26796 5294 26798 5346
rect 26850 5294 26852 5346
rect 26796 5282 26852 5294
rect 27580 5122 27636 6412
rect 27580 5070 27582 5122
rect 27634 5070 27636 5122
rect 27580 5058 27636 5070
rect 27132 4452 27188 4462
rect 27132 4358 27188 4396
rect 26684 4174 26686 4226
rect 26738 4174 26740 4226
rect 26684 4162 26740 4174
rect 27580 4228 27636 4238
rect 27580 4134 27636 4172
rect 27692 4116 27748 7868
rect 27804 7586 27860 8204
rect 27916 8194 27972 8204
rect 28028 7700 28084 8428
rect 28140 8418 28196 8428
rect 28252 8708 28308 8718
rect 28028 7634 28084 7644
rect 27804 7534 27806 7586
rect 27858 7534 27860 7586
rect 27804 7522 27860 7534
rect 28252 7364 28308 8652
rect 28476 8596 28532 8606
rect 28476 8146 28532 8540
rect 28476 8094 28478 8146
rect 28530 8094 28532 8146
rect 28364 8034 28420 8046
rect 28364 7982 28366 8034
rect 28418 7982 28420 8034
rect 28364 7474 28420 7982
rect 28364 7422 28366 7474
rect 28418 7422 28420 7474
rect 28364 7410 28420 7422
rect 28028 7308 28308 7364
rect 28028 6690 28084 7308
rect 28476 7252 28532 8094
rect 28252 7196 28532 7252
rect 28588 7924 28644 8988
rect 29932 9156 29988 9166
rect 29932 9042 29988 9100
rect 29932 8990 29934 9042
rect 29986 8990 29988 9042
rect 29932 8978 29988 8990
rect 29036 8932 29092 8942
rect 29036 8838 29092 8876
rect 29596 8370 29652 8382
rect 29596 8318 29598 8370
rect 29650 8318 29652 8370
rect 29596 8260 29652 8318
rect 29148 8034 29204 8046
rect 29148 7982 29150 8034
rect 29202 7982 29204 8034
rect 29148 7924 29204 7982
rect 28588 7868 29204 7924
rect 28252 6914 28308 7196
rect 28588 7028 28644 7868
rect 28700 7700 28756 7710
rect 28700 7474 28756 7644
rect 28700 7422 28702 7474
rect 28754 7422 28756 7474
rect 28700 7410 28756 7422
rect 28812 7586 28868 7598
rect 28812 7534 28814 7586
rect 28866 7534 28868 7586
rect 28252 6862 28254 6914
rect 28306 6862 28308 6914
rect 28252 6850 28308 6862
rect 28476 6972 28644 7028
rect 28028 6638 28030 6690
rect 28082 6638 28084 6690
rect 28028 6626 28084 6638
rect 28476 6578 28532 6972
rect 28476 6526 28478 6578
rect 28530 6526 28532 6578
rect 28476 6514 28532 6526
rect 28588 6802 28644 6814
rect 28588 6750 28590 6802
rect 28642 6750 28644 6802
rect 28588 6132 28644 6750
rect 28700 6132 28756 6142
rect 28588 6076 28700 6132
rect 28700 6066 28756 6076
rect 27804 6020 27860 6030
rect 27804 5926 27860 5964
rect 28812 6018 28868 7534
rect 29148 7362 29204 7374
rect 29148 7310 29150 7362
rect 29202 7310 29204 7362
rect 29148 6916 29204 7310
rect 29596 7364 29652 8204
rect 30044 8258 30100 9212
rect 30268 8818 30324 8830
rect 30268 8766 30270 8818
rect 30322 8766 30324 8818
rect 30268 8596 30324 8766
rect 30268 8530 30324 8540
rect 30044 8206 30046 8258
rect 30098 8206 30100 8258
rect 30044 8194 30100 8206
rect 30380 8260 30436 9324
rect 30492 9154 30548 9166
rect 30492 9102 30494 9154
rect 30546 9102 30548 9154
rect 30492 9044 30548 9102
rect 30492 8978 30548 8988
rect 30604 8930 30660 12460
rect 30716 12180 30772 12686
rect 31276 12290 31332 12908
rect 31276 12238 31278 12290
rect 31330 12238 31332 12290
rect 31276 12226 31332 12238
rect 30716 12114 30772 12124
rect 30940 12178 30996 12190
rect 30940 12126 30942 12178
rect 30994 12126 30996 12178
rect 30940 11508 30996 12126
rect 31388 12180 31444 12190
rect 31388 12086 31444 12124
rect 30940 11442 30996 11452
rect 31052 12066 31108 12078
rect 31052 12014 31054 12066
rect 31106 12014 31108 12066
rect 31052 11506 31108 12014
rect 31052 11454 31054 11506
rect 31106 11454 31108 11506
rect 31052 11442 31108 11454
rect 31500 11620 31556 11630
rect 31164 11396 31220 11406
rect 31164 11302 31220 11340
rect 31500 11394 31556 11564
rect 31500 11342 31502 11394
rect 31554 11342 31556 11394
rect 31500 11330 31556 11342
rect 30716 11284 30772 11294
rect 30772 11228 30884 11284
rect 30716 11190 30772 11228
rect 30828 10498 30884 11228
rect 30940 11172 30996 11182
rect 30940 11078 30996 11116
rect 31276 10836 31332 10846
rect 31612 10836 31668 13694
rect 31724 13412 31780 14366
rect 31724 13346 31780 13356
rect 31836 12628 31892 15092
rect 32060 14418 32116 15484
rect 32284 15316 32340 15326
rect 32284 15222 32340 15260
rect 32060 14366 32062 14418
rect 32114 14366 32116 14418
rect 32060 14354 32116 14366
rect 32396 14308 32452 16828
rect 32620 15986 32676 15998
rect 32620 15934 32622 15986
rect 32674 15934 32676 15986
rect 32508 15876 32564 15886
rect 32508 15782 32564 15820
rect 32620 15652 32676 15934
rect 32620 15586 32676 15596
rect 32732 15148 32788 17612
rect 33068 17444 33124 18172
rect 33740 18116 33796 18126
rect 33740 17780 33796 18060
rect 33180 17668 33236 17678
rect 33180 17666 33684 17668
rect 33180 17614 33182 17666
rect 33234 17614 33684 17666
rect 33180 17612 33684 17614
rect 33180 17602 33236 17612
rect 33068 17106 33124 17388
rect 33068 17054 33070 17106
rect 33122 17054 33124 17106
rect 33068 17042 33124 17054
rect 33180 17108 33236 17118
rect 33180 16100 33236 17052
rect 33628 17106 33684 17612
rect 33628 17054 33630 17106
rect 33682 17054 33684 17106
rect 33628 17042 33684 17054
rect 33740 17108 33796 17724
rect 33852 18004 33908 18014
rect 33852 17556 33908 17948
rect 33964 17780 34020 17790
rect 34076 17780 34132 18620
rect 34188 18610 34244 18620
rect 34300 17892 34356 22876
rect 34748 22596 34804 22606
rect 34748 22482 34804 22540
rect 34748 22430 34750 22482
rect 34802 22430 34804 22482
rect 34748 22418 34804 22430
rect 34524 22372 34580 22382
rect 34412 21924 34468 21934
rect 34412 21810 34468 21868
rect 34412 21758 34414 21810
rect 34466 21758 34468 21810
rect 34412 21746 34468 21758
rect 34524 21700 34580 22316
rect 35084 21812 35140 33964
rect 36204 33926 36260 33964
rect 35532 33908 35588 33918
rect 35420 33570 35476 33582
rect 35420 33518 35422 33570
rect 35474 33518 35476 33570
rect 35420 33460 35476 33518
rect 35420 33394 35476 33404
rect 35532 33348 35588 33852
rect 36428 33684 36484 34638
rect 36540 34692 36596 34702
rect 36540 34354 36596 34636
rect 36540 34302 36542 34354
rect 36594 34302 36596 34354
rect 36540 34290 36596 34302
rect 36764 34356 36820 34748
rect 37100 34738 37156 34748
rect 37324 34802 37380 34814
rect 37324 34750 37326 34802
rect 37378 34750 37380 34802
rect 36764 34262 36820 34300
rect 36876 34130 36932 34142
rect 36876 34078 36878 34130
rect 36930 34078 36932 34130
rect 36876 34020 36932 34078
rect 36876 33954 36932 33964
rect 37324 34020 37380 34750
rect 37324 33954 37380 33964
rect 37548 34690 37604 34702
rect 37548 34638 37550 34690
rect 37602 34638 37604 34690
rect 36979 33740 37243 33750
rect 37035 33684 37083 33740
rect 37139 33684 37187 33740
rect 36979 33674 37243 33684
rect 36428 33618 36484 33628
rect 35532 33254 35588 33292
rect 36428 33348 36484 33358
rect 35420 33236 35476 33246
rect 35420 33142 35476 33180
rect 36428 33122 36484 33292
rect 37100 33348 37156 33358
rect 37100 33254 37156 33292
rect 37436 33348 37492 33358
rect 36428 33070 36430 33122
rect 36482 33070 36484 33122
rect 36316 32676 36372 32686
rect 36316 32582 36372 32620
rect 36428 32116 36484 33070
rect 36988 33012 37044 33022
rect 36316 32060 36484 32116
rect 36540 32674 36596 32686
rect 36540 32622 36542 32674
rect 36594 32622 36596 32674
rect 35532 31780 35588 31790
rect 35532 31686 35588 31724
rect 35980 31778 36036 31790
rect 35980 31726 35982 31778
rect 36034 31726 36036 31778
rect 35980 31668 36036 31726
rect 36316 31668 36372 32060
rect 36428 31892 36484 31902
rect 36428 31798 36484 31836
rect 36540 31668 36596 32622
rect 36988 32674 37044 32956
rect 36988 32622 36990 32674
rect 37042 32622 37044 32674
rect 36988 32610 37044 32622
rect 36316 31612 36484 31668
rect 35980 31602 36036 31612
rect 35196 31106 35252 31118
rect 35196 31054 35198 31106
rect 35250 31054 35252 31106
rect 35196 30772 35252 31054
rect 36316 31108 36372 31118
rect 36316 31014 36372 31052
rect 36092 30884 36148 30894
rect 35196 30706 35252 30716
rect 35980 30882 36148 30884
rect 35980 30830 36094 30882
rect 36146 30830 36148 30882
rect 35980 30828 36148 30830
rect 35980 30324 36036 30828
rect 36092 30818 36148 30828
rect 35532 30100 35588 30110
rect 35532 29650 35588 30044
rect 35532 29598 35534 29650
rect 35586 29598 35588 29650
rect 35532 29586 35588 29598
rect 35420 29538 35476 29550
rect 35420 29486 35422 29538
rect 35474 29486 35476 29538
rect 35420 29428 35476 29486
rect 35980 29428 36036 30268
rect 35420 29362 35476 29372
rect 35532 29372 36036 29428
rect 36204 29652 36260 29662
rect 35308 29316 35364 29326
rect 35308 27858 35364 29260
rect 35420 28196 35476 28206
rect 35420 28082 35476 28140
rect 35420 28030 35422 28082
rect 35474 28030 35476 28082
rect 35420 28018 35476 28030
rect 35308 27806 35310 27858
rect 35362 27806 35364 27858
rect 35308 27794 35364 27806
rect 35532 27188 35588 29372
rect 36092 29316 36148 29326
rect 35644 29314 36148 29316
rect 35644 29262 36094 29314
rect 36146 29262 36148 29314
rect 35644 29260 36148 29262
rect 35644 29202 35700 29260
rect 35644 29150 35646 29202
rect 35698 29150 35700 29202
rect 35644 29138 35700 29150
rect 35868 28756 35924 28766
rect 35756 28420 35812 28430
rect 35756 28326 35812 28364
rect 35756 27972 35812 27982
rect 35644 27860 35700 27870
rect 35644 27766 35700 27804
rect 35644 27188 35700 27198
rect 35532 27186 35700 27188
rect 35532 27134 35646 27186
rect 35698 27134 35700 27186
rect 35532 27132 35700 27134
rect 35644 27122 35700 27132
rect 35756 26964 35812 27916
rect 35756 26514 35812 26908
rect 35756 26462 35758 26514
rect 35810 26462 35812 26514
rect 35756 26450 35812 26462
rect 35308 26404 35364 26414
rect 35308 26310 35364 26348
rect 35868 25732 35924 28700
rect 35980 28642 36036 29260
rect 36092 29250 36148 29260
rect 35980 28590 35982 28642
rect 36034 28590 36036 28642
rect 35980 28578 36036 28590
rect 36204 28420 36260 29596
rect 36428 28980 36484 31612
rect 36540 31602 36596 31612
rect 36652 32562 36708 32574
rect 36652 32510 36654 32562
rect 36706 32510 36708 32562
rect 36652 31556 36708 32510
rect 37436 32562 37492 33292
rect 37548 33236 37604 34638
rect 37660 33346 37716 35308
rect 38780 35252 38836 39200
rect 41020 36932 41076 39200
rect 41020 36866 41076 36876
rect 42252 36932 42308 36942
rect 41916 36820 41972 36830
rect 40796 36708 40852 36718
rect 40796 36482 40852 36652
rect 40796 36430 40798 36482
rect 40850 36430 40852 36482
rect 40796 36418 40852 36430
rect 41356 36708 41412 36718
rect 41356 36482 41412 36652
rect 41916 36594 41972 36764
rect 41916 36542 41918 36594
rect 41970 36542 41972 36594
rect 41916 36530 41972 36542
rect 41356 36430 41358 36482
rect 41410 36430 41412 36482
rect 41356 36418 41412 36430
rect 42252 36482 42308 36876
rect 43036 36932 43092 36942
rect 43036 36594 43092 36876
rect 43036 36542 43038 36594
rect 43090 36542 43092 36594
rect 43036 36530 43092 36542
rect 42252 36430 42254 36482
rect 42306 36430 42308 36482
rect 42252 36418 42308 36430
rect 39228 36370 39284 36382
rect 39228 36318 39230 36370
rect 39282 36318 39284 36370
rect 39228 35476 39284 36318
rect 39900 36372 39956 36382
rect 39900 36370 40068 36372
rect 39900 36318 39902 36370
rect 39954 36318 40068 36370
rect 39900 36316 40068 36318
rect 39900 36306 39956 36316
rect 39788 35812 39844 35822
rect 39228 35410 39284 35420
rect 39564 35810 39844 35812
rect 39564 35758 39790 35810
rect 39842 35758 39844 35810
rect 39564 35756 39844 35758
rect 38780 35186 38836 35196
rect 37884 34804 37940 34814
rect 37884 34710 37940 34748
rect 38780 34804 38836 34814
rect 37772 34690 37828 34702
rect 37772 34638 37774 34690
rect 37826 34638 37828 34690
rect 37772 34244 37828 34638
rect 38444 34690 38500 34702
rect 38444 34638 38446 34690
rect 38498 34638 38500 34690
rect 38444 34580 38500 34638
rect 38780 34580 38836 34748
rect 39564 34804 39620 35756
rect 39788 35746 39844 35756
rect 39900 35698 39956 35710
rect 39900 35646 39902 35698
rect 39954 35646 39956 35698
rect 39788 35588 39844 35598
rect 39900 35588 39956 35646
rect 39844 35532 39956 35588
rect 40012 35588 40068 36316
rect 42588 36258 42644 36270
rect 42588 36206 42590 36258
rect 42642 36206 42644 36258
rect 40908 35812 40964 35822
rect 40908 35718 40964 35756
rect 41132 35700 41188 35710
rect 41692 35700 41748 35710
rect 41132 35698 41748 35700
rect 41132 35646 41134 35698
rect 41186 35646 41694 35698
rect 41746 35646 41748 35698
rect 41132 35644 41748 35646
rect 40124 35588 40180 35598
rect 40012 35586 40180 35588
rect 40012 35534 40126 35586
rect 40178 35534 40180 35586
rect 40012 35532 40180 35534
rect 39788 35522 39844 35532
rect 39900 34916 39956 35532
rect 40012 34916 40068 34926
rect 39900 34914 40068 34916
rect 39900 34862 40014 34914
rect 40066 34862 40068 34914
rect 39900 34860 40068 34862
rect 40124 34916 40180 35532
rect 40236 35476 40292 35486
rect 40236 35382 40292 35420
rect 41020 35476 41076 35486
rect 40460 34916 40516 34926
rect 40124 34914 40516 34916
rect 40124 34862 40462 34914
rect 40514 34862 40516 34914
rect 40124 34860 40516 34862
rect 40012 34850 40068 34860
rect 40460 34850 40516 34860
rect 39564 34710 39620 34748
rect 41020 34802 41076 35420
rect 41132 35252 41188 35644
rect 41692 35634 41748 35644
rect 42252 35586 42308 35598
rect 42252 35534 42254 35586
rect 42306 35534 42308 35586
rect 41132 35186 41188 35196
rect 42140 35476 42196 35486
rect 41020 34750 41022 34802
rect 41074 34750 41076 34802
rect 41020 34738 41076 34750
rect 38444 34514 38500 34524
rect 38556 34524 38836 34580
rect 39004 34692 39060 34702
rect 37996 34244 38052 34254
rect 37772 34242 38052 34244
rect 37772 34190 37998 34242
rect 38050 34190 38052 34242
rect 37772 34188 38052 34190
rect 37996 33796 38052 34188
rect 37996 33730 38052 33740
rect 38220 34130 38276 34142
rect 38220 34078 38222 34130
rect 38274 34078 38276 34130
rect 37660 33294 37662 33346
rect 37714 33294 37716 33346
rect 37660 33282 37716 33294
rect 38220 33348 38276 34078
rect 38556 33458 38612 34524
rect 38556 33406 38558 33458
rect 38610 33406 38612 33458
rect 38556 33394 38612 33406
rect 39004 33458 39060 34636
rect 40012 34244 40068 34254
rect 40012 34150 40068 34188
rect 41580 34244 41636 34254
rect 39004 33406 39006 33458
rect 39058 33406 39060 33458
rect 39004 33394 39060 33406
rect 39116 34130 39172 34142
rect 39116 34078 39118 34130
rect 39170 34078 39172 34130
rect 38220 33282 38276 33292
rect 39116 33346 39172 34078
rect 39564 34132 39620 34142
rect 39564 34038 39620 34076
rect 40124 34132 40180 34142
rect 40124 34038 40180 34076
rect 41020 34132 41076 34142
rect 41020 34038 41076 34076
rect 41580 34130 41636 34188
rect 41580 34078 41582 34130
rect 41634 34078 41636 34130
rect 40908 34020 40964 34030
rect 40908 33926 40964 33964
rect 40012 33908 40068 33918
rect 40012 33814 40068 33852
rect 41244 33458 41300 33470
rect 41244 33406 41246 33458
rect 41298 33406 41300 33458
rect 39116 33294 39118 33346
rect 39170 33294 39172 33346
rect 37548 33170 37604 33180
rect 38780 32900 38836 32910
rect 38780 32788 38836 32844
rect 39116 32788 39172 33294
rect 39452 33348 39508 33358
rect 39452 33254 39508 33292
rect 40236 33348 40292 33358
rect 38780 32786 38948 32788
rect 38780 32734 38782 32786
rect 38834 32734 38948 32786
rect 38780 32732 38948 32734
rect 38780 32722 38836 32732
rect 38668 32676 38724 32686
rect 38668 32582 38724 32620
rect 37436 32510 37438 32562
rect 37490 32510 37492 32562
rect 36979 32172 37243 32182
rect 37035 32116 37083 32172
rect 37139 32116 37187 32172
rect 36979 32106 37243 32116
rect 37436 32002 37492 32510
rect 38444 32564 38500 32574
rect 38444 32470 38500 32508
rect 37772 32452 37828 32462
rect 37772 32358 37828 32396
rect 38668 32452 38724 32462
rect 37436 31950 37438 32002
rect 37490 31950 37492 32002
rect 37436 31938 37492 31950
rect 37884 32116 37940 32126
rect 37772 31892 37828 31902
rect 37772 31798 37828 31836
rect 37884 31778 37940 32060
rect 37884 31726 37886 31778
rect 37938 31726 37940 31778
rect 37884 31714 37940 31726
rect 36652 31490 36708 31500
rect 38108 31556 38164 31566
rect 37548 31220 37604 31230
rect 37324 31108 37380 31118
rect 36979 30604 37243 30614
rect 37035 30548 37083 30604
rect 37139 30548 37187 30604
rect 36979 30538 37243 30548
rect 36988 30100 37044 30110
rect 36988 30006 37044 30044
rect 37212 30098 37268 30110
rect 37212 30046 37214 30098
rect 37266 30046 37268 30098
rect 37100 29988 37156 29998
rect 36988 29540 37044 29550
rect 37100 29540 37156 29932
rect 36988 29538 37156 29540
rect 36988 29486 36990 29538
rect 37042 29486 37156 29538
rect 36988 29484 37156 29486
rect 36988 29474 37044 29484
rect 36428 28914 36484 28924
rect 36540 29428 36596 29438
rect 36540 28644 36596 29372
rect 37212 29316 37268 30046
rect 37324 29986 37380 31052
rect 37548 30994 37604 31164
rect 37548 30942 37550 30994
rect 37602 30942 37604 30994
rect 37548 30930 37604 30942
rect 37660 30210 37716 30222
rect 37660 30158 37662 30210
rect 37714 30158 37716 30210
rect 37660 30100 37716 30158
rect 37660 30034 37716 30044
rect 37324 29934 37326 29986
rect 37378 29934 37380 29986
rect 37324 29922 37380 29934
rect 37772 29652 37828 29662
rect 37772 29426 37828 29596
rect 37772 29374 37774 29426
rect 37826 29374 37828 29426
rect 37324 29316 37380 29326
rect 37212 29260 37324 29316
rect 37324 29222 37380 29260
rect 37772 29092 37828 29374
rect 36979 29036 37243 29046
rect 37035 28980 37083 29036
rect 37139 28980 37187 29036
rect 36979 28970 37243 28980
rect 37324 29036 37828 29092
rect 37100 28868 37156 28878
rect 36876 28644 36932 28654
rect 36540 28642 36932 28644
rect 36540 28590 36878 28642
rect 36930 28590 36932 28642
rect 36540 28588 36932 28590
rect 36876 28578 36932 28588
rect 36204 28326 36260 28364
rect 36316 28530 36372 28542
rect 36316 28478 36318 28530
rect 36370 28478 36372 28530
rect 36316 28084 36372 28478
rect 37100 28530 37156 28812
rect 37100 28478 37102 28530
rect 37154 28478 37156 28530
rect 37100 28466 37156 28478
rect 37212 28530 37268 28542
rect 37212 28478 37214 28530
rect 37266 28478 37268 28530
rect 37212 28420 37268 28478
rect 36372 28028 36820 28084
rect 36316 28018 36372 28028
rect 36316 27186 36372 27198
rect 36316 27134 36318 27186
rect 36370 27134 36372 27186
rect 35420 25676 35924 25732
rect 36092 27074 36148 27086
rect 36092 27022 36094 27074
rect 36146 27022 36148 27074
rect 36092 25732 36148 27022
rect 36204 26516 36260 26526
rect 36204 26422 36260 26460
rect 36316 26514 36372 27134
rect 36316 26462 36318 26514
rect 36370 26462 36372 26514
rect 36316 26450 36372 26462
rect 36764 26514 36820 28028
rect 37212 27972 37268 28364
rect 37212 27906 37268 27916
rect 37324 27970 37380 29036
rect 37324 27918 37326 27970
rect 37378 27918 37380 27970
rect 37324 27636 37380 27918
rect 37436 28866 37492 28878
rect 37436 28814 37438 28866
rect 37490 28814 37492 28866
rect 37436 27860 37492 28814
rect 37660 28868 37716 28878
rect 37660 28754 37716 28812
rect 37660 28702 37662 28754
rect 37714 28702 37716 28754
rect 37660 28690 37716 28702
rect 37436 27858 37716 27860
rect 37436 27806 37438 27858
rect 37490 27806 37716 27858
rect 37436 27804 37716 27806
rect 37436 27794 37492 27804
rect 37324 27580 37492 27636
rect 36979 27468 37243 27478
rect 37035 27412 37083 27468
rect 37139 27412 37187 27468
rect 36979 27402 37243 27412
rect 37100 27074 37156 27086
rect 37100 27022 37102 27074
rect 37154 27022 37156 27074
rect 37100 26908 37156 27022
rect 36764 26462 36766 26514
rect 36818 26462 36820 26514
rect 36764 26450 36820 26462
rect 36876 26852 37156 26908
rect 37324 27074 37380 27086
rect 37324 27022 37326 27074
rect 37378 27022 37380 27074
rect 36428 26068 36484 26078
rect 36876 26068 36932 26852
rect 37324 26516 37380 27022
rect 37324 26450 37380 26460
rect 37100 26292 37156 26302
rect 37100 26290 37380 26292
rect 37100 26238 37102 26290
rect 37154 26238 37380 26290
rect 37100 26236 37380 26238
rect 37100 26226 37156 26236
rect 35308 23940 35364 23950
rect 35196 23828 35252 23838
rect 35308 23828 35364 23884
rect 35196 23826 35364 23828
rect 35196 23774 35198 23826
rect 35250 23774 35364 23826
rect 35196 23772 35364 23774
rect 35196 23762 35252 23772
rect 35308 23266 35364 23278
rect 35308 23214 35310 23266
rect 35362 23214 35364 23266
rect 35196 23154 35252 23166
rect 35196 23102 35198 23154
rect 35250 23102 35252 23154
rect 35196 22820 35252 23102
rect 35196 22754 35252 22764
rect 35308 22932 35364 23214
rect 35308 22484 35364 22876
rect 35308 22418 35364 22428
rect 35308 22148 35364 22158
rect 35308 22054 35364 22092
rect 35420 21924 35476 25676
rect 36092 25666 36148 25676
rect 36316 26066 36932 26068
rect 36316 26014 36430 26066
rect 36482 26014 36932 26066
rect 36316 26012 36932 26014
rect 35644 25506 35700 25518
rect 35644 25454 35646 25506
rect 35698 25454 35700 25506
rect 35644 25172 35700 25454
rect 35868 25508 35924 25518
rect 35868 25394 35924 25452
rect 35868 25342 35870 25394
rect 35922 25342 35924 25394
rect 35868 25330 35924 25342
rect 35644 24164 35700 25116
rect 35980 25284 36036 25294
rect 35980 24722 36036 25228
rect 35980 24670 35982 24722
rect 36034 24670 36036 24722
rect 35980 24658 36036 24670
rect 36204 24612 36260 24622
rect 36204 24518 36260 24556
rect 36316 24610 36372 26012
rect 36428 26002 36484 26012
rect 36979 25900 37243 25910
rect 37035 25844 37083 25900
rect 37139 25844 37187 25900
rect 36979 25834 37243 25844
rect 36988 25732 37044 25742
rect 36988 25638 37044 25676
rect 37324 25732 37380 26236
rect 37324 25666 37380 25676
rect 37324 25396 37380 25406
rect 37324 25302 37380 25340
rect 36428 25282 36484 25294
rect 36428 25230 36430 25282
rect 36482 25230 36484 25282
rect 36428 25172 36484 25230
rect 37100 25284 37156 25294
rect 37100 25190 37156 25228
rect 36428 25106 36484 25116
rect 36764 24948 36820 24958
rect 36764 24834 36820 24892
rect 36764 24782 36766 24834
rect 36818 24782 36820 24834
rect 36764 24770 36820 24782
rect 36876 24834 36932 24846
rect 36876 24782 36878 24834
rect 36930 24782 36932 24834
rect 36316 24558 36318 24610
rect 36370 24558 36372 24610
rect 36316 24546 36372 24558
rect 36876 24500 36932 24782
rect 37100 24724 37156 24734
rect 37100 24630 37156 24668
rect 35644 24098 35700 24108
rect 36764 24444 36932 24500
rect 35532 24050 35588 24062
rect 35532 23998 35534 24050
rect 35586 23998 35588 24050
rect 35532 23380 35588 23998
rect 36092 24052 36148 24062
rect 35868 23938 35924 23950
rect 35868 23886 35870 23938
rect 35922 23886 35924 23938
rect 35868 23828 35924 23886
rect 35868 23762 35924 23772
rect 35868 23492 35924 23502
rect 35532 23378 35812 23380
rect 35532 23326 35534 23378
rect 35586 23326 35812 23378
rect 35532 23324 35812 23326
rect 35532 23314 35588 23324
rect 35756 23266 35812 23324
rect 35868 23378 35924 23436
rect 35868 23326 35870 23378
rect 35922 23326 35924 23378
rect 35868 23314 35924 23326
rect 35756 23214 35758 23266
rect 35810 23214 35812 23266
rect 35756 23202 35812 23214
rect 36092 23154 36148 23996
rect 36764 23266 36820 24444
rect 36979 24332 37243 24342
rect 37035 24276 37083 24332
rect 37139 24276 37187 24332
rect 36979 24266 37243 24276
rect 37100 23938 37156 23950
rect 37100 23886 37102 23938
rect 37154 23886 37156 23938
rect 37100 23828 37156 23886
rect 37100 23762 37156 23772
rect 37436 23548 37492 27580
rect 37548 25284 37604 25294
rect 37548 25190 37604 25228
rect 37548 24948 37604 24958
rect 37548 24052 37604 24892
rect 37548 23958 37604 23996
rect 36764 23214 36766 23266
rect 36818 23214 36820 23266
rect 36092 23102 36094 23154
rect 36146 23102 36148 23154
rect 36092 23090 36148 23102
rect 36428 23154 36484 23166
rect 36428 23102 36430 23154
rect 36482 23102 36484 23154
rect 36428 23044 36484 23102
rect 35644 22484 35700 22494
rect 35644 22390 35700 22428
rect 36204 22484 36260 22494
rect 36204 22370 36260 22428
rect 36204 22318 36206 22370
rect 36258 22318 36260 22370
rect 36204 22306 36260 22318
rect 36316 22260 36372 22270
rect 35756 22148 35812 22158
rect 35420 21868 35588 21924
rect 35084 21756 35252 21812
rect 34524 21634 34580 21644
rect 34636 21588 34692 21598
rect 35084 21588 35140 21598
rect 34636 21586 35140 21588
rect 34636 21534 34638 21586
rect 34690 21534 35086 21586
rect 35138 21534 35140 21586
rect 34636 21532 35140 21534
rect 34636 21028 34692 21532
rect 35084 21522 35140 21532
rect 34636 20962 34692 20972
rect 34972 20916 35028 20926
rect 34972 20822 35028 20860
rect 34412 20580 34468 20590
rect 34412 20578 34580 20580
rect 34412 20526 34414 20578
rect 34466 20526 34580 20578
rect 34412 20524 34580 20526
rect 34412 20514 34468 20524
rect 34524 20244 34580 20524
rect 34636 20244 34692 20254
rect 34524 20188 34636 20244
rect 34636 20178 34692 20188
rect 34412 20132 34468 20142
rect 35196 20132 35252 21756
rect 35420 21700 35476 21710
rect 35420 21606 35476 21644
rect 35420 21364 35476 21374
rect 35420 20692 35476 21308
rect 35420 20598 35476 20636
rect 34412 20130 34580 20132
rect 34412 20078 34414 20130
rect 34466 20078 34580 20130
rect 34412 20076 34580 20078
rect 34412 20066 34468 20076
rect 34412 19460 34468 19470
rect 34412 19366 34468 19404
rect 34524 19236 34580 20076
rect 35196 20066 35252 20076
rect 34300 17826 34356 17836
rect 34412 18450 34468 18462
rect 34412 18398 34414 18450
rect 34466 18398 34468 18450
rect 33964 17778 34132 17780
rect 33964 17726 33966 17778
rect 34018 17726 34132 17778
rect 33964 17724 34132 17726
rect 33964 17714 34020 17724
rect 34412 17668 34468 18398
rect 34524 17892 34580 19180
rect 34636 20018 34692 20030
rect 34636 19966 34638 20018
rect 34690 19966 34692 20018
rect 34636 19684 34692 19966
rect 35308 20020 35364 20030
rect 35308 19926 35364 19964
rect 34636 19236 34692 19628
rect 35308 19348 35364 19358
rect 34748 19236 34804 19246
rect 34636 19180 34748 19236
rect 34636 19122 34692 19180
rect 34748 19170 34804 19180
rect 35308 19234 35364 19292
rect 35532 19236 35588 21868
rect 35308 19182 35310 19234
rect 35362 19182 35364 19234
rect 34636 19070 34638 19122
rect 34690 19070 34692 19122
rect 34636 19058 34692 19070
rect 35308 18676 35364 19182
rect 35308 18610 35364 18620
rect 35420 19180 35588 19236
rect 35644 21252 35700 21262
rect 34860 18562 34916 18574
rect 34860 18510 34862 18562
rect 34914 18510 34916 18562
rect 34636 18452 34692 18462
rect 34636 18358 34692 18396
rect 34860 18116 34916 18510
rect 34972 18564 35028 18574
rect 34972 18562 35140 18564
rect 34972 18510 34974 18562
rect 35026 18510 35140 18562
rect 34972 18508 35140 18510
rect 34972 18498 35028 18508
rect 34860 18050 34916 18060
rect 34972 17892 35028 17902
rect 34524 17890 35028 17892
rect 34524 17838 34974 17890
rect 35026 17838 35028 17890
rect 34524 17836 35028 17838
rect 34972 17826 35028 17836
rect 35084 17780 35140 18508
rect 35420 18116 35476 19180
rect 35532 19010 35588 19022
rect 35532 18958 35534 19010
rect 35586 18958 35588 19010
rect 35532 18900 35588 18958
rect 35532 18834 35588 18844
rect 35644 18676 35700 21196
rect 35756 19572 35812 22092
rect 36092 21698 36148 21710
rect 36092 21646 36094 21698
rect 36146 21646 36148 21698
rect 36092 21252 36148 21646
rect 36092 21186 36148 21196
rect 36204 21586 36260 21598
rect 36204 21534 36206 21586
rect 36258 21534 36260 21586
rect 36092 20802 36148 20814
rect 36092 20750 36094 20802
rect 36146 20750 36148 20802
rect 36092 20356 36148 20750
rect 36204 20468 36260 21534
rect 36316 21474 36372 22204
rect 36428 22036 36484 22988
rect 36764 22484 36820 23214
rect 37212 23492 37492 23548
rect 37548 23716 37604 23726
rect 37212 23268 37268 23492
rect 37548 23378 37604 23660
rect 37548 23326 37550 23378
rect 37602 23326 37604 23378
rect 37548 23314 37604 23326
rect 37212 23212 37492 23268
rect 37212 23042 37268 23054
rect 37212 22990 37214 23042
rect 37266 22990 37268 23042
rect 37212 22932 37268 22990
rect 37212 22866 37268 22876
rect 37324 22820 37380 22830
rect 36979 22764 37243 22774
rect 37035 22708 37083 22764
rect 37139 22708 37187 22764
rect 36979 22698 37243 22708
rect 36764 22418 36820 22428
rect 36988 22596 37044 22606
rect 36988 22258 37044 22540
rect 37324 22370 37380 22764
rect 37324 22318 37326 22370
rect 37378 22318 37380 22370
rect 37324 22306 37380 22318
rect 36988 22206 36990 22258
rect 37042 22206 37044 22258
rect 36988 22194 37044 22206
rect 36428 21970 36484 21980
rect 36876 21698 36932 21710
rect 36876 21646 36878 21698
rect 36930 21646 36932 21698
rect 36764 21588 36820 21598
rect 36316 21422 36318 21474
rect 36370 21422 36372 21474
rect 36316 21410 36372 21422
rect 36428 21586 36820 21588
rect 36428 21534 36766 21586
rect 36818 21534 36820 21586
rect 36428 21532 36820 21534
rect 36428 21028 36484 21532
rect 36764 21522 36820 21532
rect 36876 21364 36932 21646
rect 37436 21700 37492 23212
rect 37660 22484 37716 27804
rect 37996 27188 38052 27198
rect 38108 27188 38164 31500
rect 38668 31106 38724 32396
rect 38780 32338 38836 32350
rect 38780 32286 38782 32338
rect 38834 32286 38836 32338
rect 38780 32116 38836 32286
rect 38780 32050 38836 32060
rect 38892 31892 38948 32732
rect 39116 32722 39172 32732
rect 40012 32900 40068 32910
rect 39340 32674 39396 32686
rect 39340 32622 39342 32674
rect 39394 32622 39396 32674
rect 39116 32564 39172 32574
rect 39116 32470 39172 32508
rect 39340 32116 39396 32622
rect 39340 32050 39396 32060
rect 39452 32562 39508 32574
rect 39452 32510 39454 32562
rect 39506 32510 39508 32562
rect 38780 31836 38948 31892
rect 39452 31892 39508 32510
rect 38780 31780 38836 31836
rect 39452 31826 39508 31836
rect 38780 31714 38836 31724
rect 39676 31780 39732 31790
rect 39676 31686 39732 31724
rect 38892 31668 38948 31678
rect 38892 31574 38948 31612
rect 39228 31554 39284 31566
rect 39228 31502 39230 31554
rect 39282 31502 39284 31554
rect 39228 31220 39284 31502
rect 39228 31154 39284 31164
rect 40012 31218 40068 32844
rect 40236 32450 40292 33292
rect 40572 33348 40628 33358
rect 41244 33348 41300 33406
rect 40572 33346 41188 33348
rect 40572 33294 40574 33346
rect 40626 33294 41188 33346
rect 40572 33292 41188 33294
rect 40572 33282 40628 33292
rect 40348 33236 40404 33246
rect 40348 33234 40516 33236
rect 40348 33182 40350 33234
rect 40402 33182 40516 33234
rect 40348 33180 40516 33182
rect 40348 33170 40404 33180
rect 40348 32564 40404 32574
rect 40460 32564 40516 33180
rect 40796 33124 40852 33134
rect 40796 33030 40852 33068
rect 40908 33124 40964 33134
rect 40908 33122 41076 33124
rect 40908 33070 40910 33122
rect 40962 33070 41076 33122
rect 40908 33068 41076 33070
rect 40908 33058 40964 33068
rect 40460 32508 40964 32564
rect 40348 32470 40404 32508
rect 40236 32398 40238 32450
rect 40290 32398 40292 32450
rect 40012 31166 40014 31218
rect 40066 31166 40068 31218
rect 40012 31154 40068 31166
rect 40124 31778 40180 31790
rect 40124 31726 40126 31778
rect 40178 31726 40180 31778
rect 40124 31220 40180 31726
rect 40124 31154 40180 31164
rect 38668 31054 38670 31106
rect 38722 31054 38724 31106
rect 38668 31042 38724 31054
rect 40236 30884 40292 32398
rect 40908 32450 40964 32508
rect 40908 32398 40910 32450
rect 40962 32398 40964 32450
rect 40908 32386 40964 32398
rect 40572 31780 40628 31790
rect 40572 31686 40628 31724
rect 41020 31778 41076 33068
rect 41020 31726 41022 31778
rect 41074 31726 41076 31778
rect 41020 31714 41076 31726
rect 41132 32452 41188 33292
rect 41244 33282 41300 33292
rect 41468 32564 41524 32574
rect 41468 32470 41524 32508
rect 41132 31666 41188 32396
rect 41132 31614 41134 31666
rect 41186 31614 41188 31666
rect 41132 31602 41188 31614
rect 41244 32340 41300 32350
rect 41244 31444 41300 32284
rect 41356 31780 41412 31790
rect 41580 31780 41636 34078
rect 41692 33234 41748 33246
rect 41692 33182 41694 33234
rect 41746 33182 41748 33234
rect 41692 33124 41748 33182
rect 41692 32228 41748 33068
rect 41916 32676 41972 32714
rect 41916 32610 41972 32620
rect 42028 32562 42084 32574
rect 42028 32510 42030 32562
rect 42082 32510 42084 32562
rect 41804 32452 41860 32462
rect 41804 32340 41860 32396
rect 41916 32340 41972 32350
rect 41804 32338 41972 32340
rect 41804 32286 41918 32338
rect 41970 32286 41972 32338
rect 41804 32284 41972 32286
rect 41916 32274 41972 32284
rect 42028 32340 42084 32510
rect 42028 32274 42084 32284
rect 41692 32172 41860 32228
rect 41804 31892 41860 32172
rect 42028 32116 42084 32126
rect 42028 31892 42084 32060
rect 41804 31826 41860 31836
rect 41916 31836 42084 31892
rect 41356 31778 41636 31780
rect 41356 31726 41358 31778
rect 41410 31726 41636 31778
rect 41356 31724 41636 31726
rect 41356 31714 41412 31724
rect 41020 31388 41300 31444
rect 41804 31668 41860 31678
rect 40908 31220 40964 31230
rect 40908 31126 40964 31164
rect 40124 30828 40292 30884
rect 40348 30994 40404 31006
rect 40348 30942 40350 30994
rect 40402 30942 40404 30994
rect 40348 30884 40404 30942
rect 39340 30660 39396 30670
rect 38556 30322 38612 30334
rect 38556 30270 38558 30322
rect 38610 30270 38612 30322
rect 38556 29540 38612 30270
rect 38780 30098 38836 30110
rect 38780 30046 38782 30098
rect 38834 30046 38836 30098
rect 38780 29652 38836 30046
rect 38780 29586 38836 29596
rect 38220 29484 38612 29540
rect 38220 29426 38276 29484
rect 38220 29374 38222 29426
rect 38274 29374 38276 29426
rect 38220 28866 38276 29374
rect 38220 28814 38222 28866
rect 38274 28814 38276 28866
rect 38220 28802 38276 28814
rect 38780 28642 38836 28654
rect 38780 28590 38782 28642
rect 38834 28590 38836 28642
rect 38220 28420 38276 28430
rect 38668 28420 38724 28430
rect 38276 28364 38388 28420
rect 38220 28326 38276 28364
rect 38220 27860 38276 27870
rect 38220 27766 38276 27804
rect 37996 27186 38164 27188
rect 37996 27134 37998 27186
rect 38050 27134 38164 27186
rect 37996 27132 38164 27134
rect 37996 27122 38052 27132
rect 38332 27076 38388 28364
rect 38668 28326 38724 28364
rect 38780 28084 38836 28590
rect 39340 28644 39396 30604
rect 40012 30212 40068 30222
rect 40012 30118 40068 30156
rect 39900 29426 39956 29438
rect 39900 29374 39902 29426
rect 39954 29374 39956 29426
rect 39340 28578 39396 28588
rect 39564 29314 39620 29326
rect 39564 29262 39566 29314
rect 39618 29262 39620 29314
rect 39564 28644 39620 29262
rect 39900 28756 39956 29374
rect 39900 28644 39956 28700
rect 39900 28588 40068 28644
rect 38780 28018 38836 28028
rect 39564 27970 39620 28588
rect 39676 28532 39732 28542
rect 39676 28530 39956 28532
rect 39676 28478 39678 28530
rect 39730 28478 39956 28530
rect 39676 28476 39956 28478
rect 39676 28466 39732 28476
rect 39900 28082 39956 28476
rect 39900 28030 39902 28082
rect 39954 28030 39956 28082
rect 39900 28018 39956 28030
rect 39564 27918 39566 27970
rect 39618 27918 39620 27970
rect 39564 27906 39620 27918
rect 40012 27748 40068 28588
rect 38332 27010 38388 27020
rect 39564 27746 40068 27748
rect 39564 27694 40014 27746
rect 40066 27694 40068 27746
rect 39564 27692 40068 27694
rect 38892 26850 38948 26862
rect 38892 26798 38894 26850
rect 38946 26798 38948 26850
rect 38332 26402 38388 26414
rect 38332 26350 38334 26402
rect 38386 26350 38388 26402
rect 38220 26290 38276 26302
rect 38220 26238 38222 26290
rect 38274 26238 38276 26290
rect 37996 26178 38052 26190
rect 37996 26126 37998 26178
rect 38050 26126 38052 26178
rect 37996 25956 38052 26126
rect 37884 25844 37940 25854
rect 37772 25508 37828 25518
rect 37772 25394 37828 25452
rect 37772 25342 37774 25394
rect 37826 25342 37828 25394
rect 37772 25330 37828 25342
rect 37884 25394 37940 25788
rect 37996 25732 38052 25900
rect 38220 25956 38276 26238
rect 38332 26292 38388 26350
rect 38332 26226 38388 26236
rect 38556 26292 38612 26302
rect 38556 26198 38612 26236
rect 38892 26180 38948 26798
rect 39116 26180 39172 26190
rect 38892 26178 39172 26180
rect 38892 26126 39118 26178
rect 39170 26126 39172 26178
rect 38892 26124 39172 26126
rect 38220 25890 38276 25900
rect 39116 25956 39172 26124
rect 37996 25676 39060 25732
rect 38220 25506 38276 25676
rect 38220 25454 38222 25506
rect 38274 25454 38276 25506
rect 38220 25442 38276 25454
rect 38332 25508 38388 25518
rect 37884 25342 37886 25394
rect 37938 25342 37940 25394
rect 37884 25330 37940 25342
rect 38332 25394 38388 25452
rect 38556 25508 38612 25518
rect 38556 25414 38612 25452
rect 38332 25342 38334 25394
rect 38386 25342 38388 25394
rect 38332 25330 38388 25342
rect 38780 25394 38836 25406
rect 38780 25342 38782 25394
rect 38834 25342 38836 25394
rect 38780 25060 38836 25342
rect 38444 25004 38836 25060
rect 38892 25282 38948 25294
rect 38892 25230 38894 25282
rect 38946 25230 38948 25282
rect 38108 24836 38164 24846
rect 38108 24742 38164 24780
rect 38444 24724 38500 25004
rect 38444 24630 38500 24668
rect 37996 24610 38052 24622
rect 37996 24558 37998 24610
rect 38050 24558 38052 24610
rect 37884 24276 37940 24286
rect 37772 23266 37828 23278
rect 37772 23214 37774 23266
rect 37826 23214 37828 23266
rect 37772 22820 37828 23214
rect 37884 23268 37940 24220
rect 37996 24052 38052 24558
rect 37996 23986 38052 23996
rect 38108 24612 38164 24622
rect 37884 23174 37940 23212
rect 37996 23716 38052 23726
rect 37772 22754 37828 22764
rect 37996 22708 38052 23660
rect 37996 22642 38052 22652
rect 37772 22596 37828 22606
rect 37772 22502 37828 22540
rect 37436 21634 37492 21644
rect 37548 22428 37716 22484
rect 37100 21588 37156 21598
rect 37100 21586 37380 21588
rect 37100 21534 37102 21586
rect 37154 21534 37380 21586
rect 37100 21532 37380 21534
rect 37100 21522 37156 21532
rect 36204 20402 36260 20412
rect 36316 20972 36484 21028
rect 36652 21308 36932 21364
rect 36316 20802 36372 20972
rect 36316 20750 36318 20802
rect 36370 20750 36372 20802
rect 36092 20290 36148 20300
rect 35980 20132 36036 20142
rect 36316 20132 36372 20750
rect 36428 20804 36484 20814
rect 36428 20710 36484 20748
rect 35980 20130 36372 20132
rect 35980 20078 35982 20130
rect 36034 20078 36372 20130
rect 35980 20076 36372 20078
rect 35980 20066 36036 20076
rect 36316 20020 36372 20076
rect 36652 20356 36708 21308
rect 36979 21196 37243 21206
rect 37035 21140 37083 21196
rect 37139 21140 37187 21196
rect 36979 21130 37243 21140
rect 37324 20802 37380 21532
rect 37436 21474 37492 21486
rect 37436 21422 37438 21474
rect 37490 21422 37492 21474
rect 37436 21364 37492 21422
rect 37436 21298 37492 21308
rect 37436 20916 37492 20926
rect 37436 20822 37492 20860
rect 37324 20750 37326 20802
rect 37378 20750 37380 20802
rect 37324 20738 37380 20750
rect 37548 20580 37604 22428
rect 38108 22372 38164 24556
rect 38220 24388 38276 24398
rect 38220 23380 38276 24332
rect 38220 22932 38276 23324
rect 38444 24052 38500 24062
rect 38332 23044 38388 23054
rect 38332 22950 38388 22988
rect 38220 22866 38276 22876
rect 38220 22596 38276 22606
rect 38444 22596 38500 23996
rect 38556 23940 38612 25004
rect 38892 24948 38948 25230
rect 38668 24892 38892 24948
rect 38668 24834 38724 24892
rect 38892 24882 38948 24892
rect 38668 24782 38670 24834
rect 38722 24782 38724 24834
rect 38668 24770 38724 24782
rect 38892 24724 38948 24734
rect 38780 24612 38836 24622
rect 38780 24518 38836 24556
rect 38556 23874 38612 23884
rect 38556 23492 38612 23502
rect 38556 23156 38612 23436
rect 38556 23090 38612 23100
rect 38780 23044 38836 23054
rect 38220 22594 38500 22596
rect 38220 22542 38222 22594
rect 38274 22542 38500 22594
rect 38220 22540 38500 22542
rect 38668 23042 38836 23044
rect 38668 22990 38782 23042
rect 38834 22990 38836 23042
rect 38668 22988 38836 22990
rect 38220 22530 38276 22540
rect 38332 22372 38388 22382
rect 38108 22370 38388 22372
rect 38108 22318 38334 22370
rect 38386 22318 38388 22370
rect 38108 22316 38388 22318
rect 37660 22260 37716 22270
rect 37884 22260 37940 22270
rect 37660 22166 37716 22204
rect 37772 22204 37884 22260
rect 37772 21810 37828 22204
rect 37884 22194 37940 22204
rect 38108 22260 38164 22316
rect 38332 22306 38388 22316
rect 38444 22372 38500 22382
rect 38108 22194 38164 22204
rect 38220 22148 38276 22158
rect 38444 22148 38500 22316
rect 38220 22146 38500 22148
rect 38220 22094 38222 22146
rect 38274 22094 38500 22146
rect 38220 22092 38500 22094
rect 38220 22082 38276 22092
rect 37772 21758 37774 21810
rect 37826 21758 37828 21810
rect 37772 21252 37828 21758
rect 38108 22036 38164 22046
rect 38108 21810 38164 21980
rect 38108 21758 38110 21810
rect 38162 21758 38164 21810
rect 38108 21746 38164 21758
rect 38444 21812 38500 21822
rect 37772 21186 37828 21196
rect 37996 21700 38052 21710
rect 37324 20524 37604 20580
rect 37660 21140 37716 21150
rect 36428 20020 36484 20030
rect 36316 20018 36484 20020
rect 36316 19966 36430 20018
rect 36482 19966 36484 20018
rect 36316 19964 36484 19966
rect 36428 19954 36484 19964
rect 36652 20018 36708 20300
rect 36652 19966 36654 20018
rect 36706 19966 36708 20018
rect 36204 19908 36260 19918
rect 35756 19516 36148 19572
rect 35980 19348 36036 19358
rect 35980 19254 36036 19292
rect 35756 19234 35812 19246
rect 35756 19182 35758 19234
rect 35810 19182 35812 19234
rect 35756 19124 35812 19182
rect 35756 19058 35812 19068
rect 36092 19124 36148 19516
rect 36204 19234 36260 19852
rect 36204 19182 36206 19234
rect 36258 19182 36260 19234
rect 36204 19170 36260 19182
rect 36092 19058 36148 19068
rect 36428 19122 36484 19134
rect 36428 19070 36430 19122
rect 36482 19070 36484 19122
rect 36428 18900 36484 19070
rect 36484 18844 36596 18900
rect 36428 18834 36484 18844
rect 36316 18676 36372 18686
rect 35644 18620 35812 18676
rect 34412 17602 34468 17612
rect 34748 17668 34804 17678
rect 35084 17668 35140 17724
rect 34748 17574 34804 17612
rect 34860 17612 35140 17668
rect 35196 18060 35476 18116
rect 35532 18338 35588 18350
rect 35532 18286 35534 18338
rect 35586 18286 35588 18338
rect 35532 18116 35588 18286
rect 35756 18116 35812 18620
rect 36316 18582 36372 18620
rect 36540 18564 36596 18844
rect 36652 18676 36708 19966
rect 36764 20468 36820 20478
rect 36764 19460 36820 20412
rect 37324 20130 37380 20524
rect 37324 20078 37326 20130
rect 37378 20078 37380 20130
rect 37324 20066 37380 20078
rect 37660 20018 37716 21084
rect 37996 20692 38052 21644
rect 38444 21698 38500 21756
rect 38444 21646 38446 21698
rect 38498 21646 38500 21698
rect 38444 21634 38500 21646
rect 38668 21700 38724 22988
rect 38780 22978 38836 22988
rect 38668 21634 38724 21644
rect 38780 22820 38836 22830
rect 38780 22482 38836 22764
rect 38780 22430 38782 22482
rect 38834 22430 38836 22482
rect 38108 20804 38164 20814
rect 38108 20710 38164 20748
rect 37996 20626 38052 20636
rect 38780 20356 38836 22430
rect 38556 20300 38836 20356
rect 37660 19966 37662 20018
rect 37714 19966 37716 20018
rect 37548 19908 37604 19918
rect 36979 19628 37243 19638
rect 37035 19572 37083 19628
rect 37139 19572 37187 19628
rect 36979 19562 37243 19572
rect 36764 19404 36932 19460
rect 36764 18676 36820 18686
rect 36652 18620 36764 18676
rect 36764 18610 36820 18620
rect 36540 18508 36708 18564
rect 36652 18452 36708 18508
rect 36764 18452 36820 18462
rect 36652 18450 36820 18452
rect 36652 18398 36766 18450
rect 36818 18398 36820 18450
rect 36652 18396 36820 18398
rect 36764 18386 36820 18396
rect 36876 18452 36932 19404
rect 37212 19236 37268 19246
rect 36876 18386 36932 18396
rect 36988 19234 37268 19236
rect 36988 19182 37214 19234
rect 37266 19182 37268 19234
rect 36988 19180 37268 19182
rect 35532 18060 35812 18116
rect 35868 18340 35924 18350
rect 35196 17668 35252 18060
rect 35868 18004 35924 18284
rect 36988 18228 37044 19180
rect 37212 19170 37268 19180
rect 37548 18788 37604 19852
rect 37660 19684 37716 19966
rect 37660 19618 37716 19628
rect 37884 20132 37940 20142
rect 37548 18722 37604 18732
rect 37660 19236 37716 19246
rect 37100 18620 37492 18676
rect 37100 18450 37156 18620
rect 37100 18398 37102 18450
rect 37154 18398 37156 18450
rect 37100 18386 37156 18398
rect 37324 18452 37380 18462
rect 37436 18452 37492 18620
rect 37548 18452 37604 18462
rect 37436 18450 37604 18452
rect 37436 18398 37550 18450
rect 37602 18398 37604 18450
rect 37436 18396 37604 18398
rect 37324 18358 37380 18396
rect 37548 18386 37604 18396
rect 35868 17938 35924 17948
rect 36764 18172 36988 18228
rect 37212 18338 37268 18350
rect 37212 18286 37214 18338
rect 37266 18286 37268 18338
rect 37212 18228 37268 18286
rect 37212 18172 37380 18228
rect 35308 17892 35364 17902
rect 35756 17892 35812 17902
rect 35308 17890 35812 17892
rect 35308 17838 35310 17890
rect 35362 17838 35758 17890
rect 35810 17838 35812 17890
rect 35308 17836 35812 17838
rect 35308 17826 35364 17836
rect 35756 17826 35812 17836
rect 35532 17668 35588 17678
rect 36316 17668 36372 17678
rect 35196 17612 35476 17668
rect 34188 17556 34244 17566
rect 33852 17500 34132 17556
rect 33740 17042 33796 17052
rect 33404 16996 33460 17006
rect 33404 16902 33460 16940
rect 33852 16996 33908 17006
rect 33852 16902 33908 16940
rect 33964 16884 34020 16894
rect 33964 16790 34020 16828
rect 34076 16660 34132 17500
rect 34188 17554 34356 17556
rect 34188 17502 34190 17554
rect 34242 17502 34356 17554
rect 34188 17500 34356 17502
rect 34188 17490 34244 17500
rect 34076 16594 34132 16604
rect 33180 16098 33796 16100
rect 33180 16046 33182 16098
rect 33234 16046 33796 16098
rect 33180 16044 33796 16046
rect 33180 16034 33236 16044
rect 32844 15988 32900 15998
rect 32844 15316 32900 15932
rect 32956 15876 33012 15886
rect 32956 15782 33012 15820
rect 33628 15874 33684 15886
rect 33628 15822 33630 15874
rect 33682 15822 33684 15874
rect 33404 15764 33460 15774
rect 32844 15250 32900 15260
rect 32956 15652 33012 15662
rect 32732 15092 32900 15148
rect 32508 14308 32564 14318
rect 32396 14252 32508 14308
rect 32508 14214 32564 14252
rect 32844 14084 32900 15092
rect 32956 14530 33012 15596
rect 32956 14478 32958 14530
rect 33010 14478 33012 14530
rect 32956 14466 33012 14478
rect 33404 15316 33460 15708
rect 33628 15652 33684 15822
rect 33628 15586 33684 15596
rect 33740 15538 33796 16044
rect 33740 15486 33742 15538
rect 33794 15486 33796 15538
rect 33740 15474 33796 15486
rect 33964 15874 34020 15886
rect 33964 15822 33966 15874
rect 34018 15822 34020 15874
rect 33404 14420 33460 15260
rect 33516 15428 33572 15438
rect 33516 14756 33572 15372
rect 33628 15314 33684 15326
rect 33628 15262 33630 15314
rect 33682 15262 33684 15314
rect 33628 14868 33684 15262
rect 33964 15316 34020 15822
rect 34300 15316 34356 17500
rect 34412 17444 34468 17454
rect 34412 17350 34468 17388
rect 34636 17442 34692 17454
rect 34636 17390 34638 17442
rect 34690 17390 34692 17442
rect 34636 16996 34692 17390
rect 34748 17108 34804 17118
rect 34748 17014 34804 17052
rect 34636 16930 34692 16940
rect 34412 16884 34468 16894
rect 34412 16210 34468 16828
rect 34412 16158 34414 16210
rect 34466 16158 34468 16210
rect 34412 16146 34468 16158
rect 34412 15372 34692 15428
rect 34412 15316 34468 15372
rect 34300 15314 34468 15316
rect 34300 15262 34414 15314
rect 34466 15262 34468 15314
rect 34300 15260 34468 15262
rect 33964 15250 34020 15260
rect 34412 15250 34468 15260
rect 34524 15202 34580 15214
rect 34524 15150 34526 15202
rect 34578 15150 34580 15202
rect 34524 15148 34580 15150
rect 33740 15092 34580 15148
rect 33740 15090 33796 15092
rect 33740 15038 33742 15090
rect 33794 15038 33796 15090
rect 33740 15026 33796 15038
rect 34636 14868 34692 15372
rect 33628 14812 33908 14868
rect 33516 14700 33684 14756
rect 33628 14642 33684 14700
rect 33628 14590 33630 14642
rect 33682 14590 33684 14642
rect 33628 14578 33684 14590
rect 33404 14364 33572 14420
rect 33068 14308 33124 14318
rect 33068 14214 33124 14252
rect 33292 14308 33348 14318
rect 33292 14306 33460 14308
rect 33292 14254 33294 14306
rect 33346 14254 33460 14306
rect 33292 14252 33460 14254
rect 33292 14242 33348 14252
rect 32844 14028 33236 14084
rect 33180 13970 33236 14028
rect 33180 13918 33182 13970
rect 33234 13918 33236 13970
rect 33180 13906 33236 13918
rect 31948 13860 32004 13870
rect 33068 13860 33124 13870
rect 31948 13858 33124 13860
rect 31948 13806 31950 13858
rect 32002 13806 33070 13858
rect 33122 13806 33124 13858
rect 31948 13804 33124 13806
rect 31948 13794 32004 13804
rect 33068 13794 33124 13804
rect 33292 13746 33348 13758
rect 33292 13694 33294 13746
rect 33346 13694 33348 13746
rect 32060 13636 32116 13646
rect 32284 13636 32340 13646
rect 32116 13580 32228 13636
rect 32060 13570 32116 13580
rect 31836 12562 31892 12572
rect 32060 12404 32116 12414
rect 31724 12402 32116 12404
rect 31724 12350 32062 12402
rect 32114 12350 32116 12402
rect 31724 12348 32116 12350
rect 31724 11282 31780 12348
rect 32060 12338 32116 12348
rect 31948 12178 32004 12190
rect 31948 12126 31950 12178
rect 32002 12126 32004 12178
rect 31948 11620 32004 12126
rect 32172 11956 32228 13580
rect 32284 13542 32340 13580
rect 32508 13636 32564 13646
rect 32396 13524 32452 13534
rect 32396 12850 32452 13468
rect 32508 12964 32564 13580
rect 33292 13524 33348 13694
rect 33404 13636 33460 14252
rect 33404 13570 33460 13580
rect 33292 13458 33348 13468
rect 32732 12964 32788 12974
rect 32508 12962 32788 12964
rect 32508 12910 32734 12962
rect 32786 12910 32788 12962
rect 32508 12908 32788 12910
rect 32732 12898 32788 12908
rect 32396 12798 32398 12850
rect 32450 12798 32452 12850
rect 32396 12786 32452 12798
rect 32284 12404 32340 12414
rect 33404 12404 33460 12414
rect 33516 12404 33572 14364
rect 33740 13972 33796 13982
rect 32284 12402 33348 12404
rect 32284 12350 32286 12402
rect 32338 12350 33348 12402
rect 32284 12348 33348 12350
rect 32284 12338 32340 12348
rect 33180 12178 33236 12190
rect 33180 12126 33182 12178
rect 33234 12126 33236 12178
rect 33180 12068 33236 12126
rect 33180 12002 33236 12012
rect 32172 11890 32228 11900
rect 33068 11956 33124 11966
rect 32508 11844 32564 11854
rect 32564 11788 32676 11844
rect 32508 11778 32564 11788
rect 31948 11564 32116 11620
rect 31836 11508 31892 11518
rect 31836 11396 31892 11452
rect 31948 11396 32004 11406
rect 31836 11394 32004 11396
rect 31836 11342 31950 11394
rect 32002 11342 32004 11394
rect 31836 11340 32004 11342
rect 31948 11330 32004 11340
rect 32060 11394 32116 11564
rect 32060 11342 32062 11394
rect 32114 11342 32116 11394
rect 31724 11230 31726 11282
rect 31778 11230 31780 11282
rect 31724 11060 31780 11230
rect 32060 11284 32116 11342
rect 32396 11508 32452 11518
rect 32396 11394 32452 11452
rect 32396 11342 32398 11394
rect 32450 11342 32452 11394
rect 32396 11330 32452 11342
rect 32060 11218 32116 11228
rect 31724 10994 31780 11004
rect 32508 11170 32564 11182
rect 32508 11118 32510 11170
rect 32562 11118 32564 11170
rect 32172 10836 32228 10846
rect 31612 10780 32004 10836
rect 31052 10722 31108 10734
rect 31052 10670 31054 10722
rect 31106 10670 31108 10722
rect 30828 10446 30830 10498
rect 30882 10446 30884 10498
rect 30828 10434 30884 10446
rect 30940 10610 30996 10622
rect 30940 10558 30942 10610
rect 30994 10558 30996 10610
rect 30604 8878 30606 8930
rect 30658 8878 30660 8930
rect 30604 8866 30660 8878
rect 30716 9826 30772 9838
rect 30716 9774 30718 9826
rect 30770 9774 30772 9826
rect 30716 8596 30772 9774
rect 30940 9826 30996 10558
rect 30940 9774 30942 9826
rect 30994 9774 30996 9826
rect 30940 9604 30996 9774
rect 30716 8530 30772 8540
rect 30828 9548 30940 9604
rect 30604 8372 30660 8382
rect 30828 8372 30884 9548
rect 30940 9538 30996 9548
rect 31052 9492 31108 10670
rect 31052 9426 31108 9436
rect 31164 10164 31220 10174
rect 31164 9266 31220 10108
rect 31164 9214 31166 9266
rect 31218 9214 31220 9266
rect 31164 9202 31220 9214
rect 31276 9266 31332 10780
rect 31500 10724 31556 10734
rect 31556 10668 31780 10724
rect 31500 10658 31556 10668
rect 31724 10610 31780 10668
rect 31724 10558 31726 10610
rect 31778 10558 31780 10610
rect 31724 10386 31780 10558
rect 31724 10334 31726 10386
rect 31778 10334 31780 10386
rect 31724 10322 31780 10334
rect 31724 9940 31780 9950
rect 31388 9716 31444 9726
rect 31388 9622 31444 9660
rect 31724 9714 31780 9884
rect 31724 9662 31726 9714
rect 31778 9662 31780 9714
rect 31724 9650 31780 9662
rect 31276 9214 31278 9266
rect 31330 9214 31332 9266
rect 31276 9202 31332 9214
rect 31724 9268 31780 9278
rect 30604 8370 30884 8372
rect 30604 8318 30606 8370
rect 30658 8318 30884 8370
rect 30604 8316 30884 8318
rect 30604 8306 30660 8316
rect 29825 7868 30089 7878
rect 29881 7812 29929 7868
rect 29985 7812 30033 7868
rect 29825 7802 30089 7812
rect 30380 7588 30436 8204
rect 30828 7698 30884 8316
rect 31052 9042 31108 9054
rect 31052 8990 31054 9042
rect 31106 8990 31108 9042
rect 31052 8484 31108 8990
rect 31724 9042 31780 9212
rect 31948 9156 32004 10780
rect 32172 10742 32228 10780
rect 32060 10386 32116 10398
rect 32060 10334 32062 10386
rect 32114 10334 32116 10386
rect 32060 10276 32116 10334
rect 32060 9826 32116 10220
rect 32508 9940 32564 11118
rect 32508 9874 32564 9884
rect 32620 11060 32676 11788
rect 32732 11284 32788 11294
rect 32732 11282 32900 11284
rect 32732 11230 32734 11282
rect 32786 11230 32900 11282
rect 32732 11228 32900 11230
rect 32732 11218 32788 11228
rect 32844 11172 32900 11228
rect 32844 11106 32900 11116
rect 32620 9940 32676 11004
rect 33068 10834 33124 11900
rect 33292 11394 33348 12348
rect 33404 12402 33572 12404
rect 33404 12350 33406 12402
rect 33458 12350 33572 12402
rect 33404 12348 33572 12350
rect 33404 12338 33460 12348
rect 33516 11732 33572 12348
rect 33628 13748 33684 13758
rect 33628 12962 33684 13692
rect 33740 13746 33796 13916
rect 33740 13694 33742 13746
rect 33794 13694 33796 13746
rect 33740 13682 33796 13694
rect 33628 12910 33630 12962
rect 33682 12910 33684 12962
rect 33628 12402 33684 12910
rect 33852 12516 33908 14812
rect 34300 14812 34692 14868
rect 34076 14308 34132 14318
rect 33964 13636 34020 13646
rect 33964 13542 34020 13580
rect 33964 12852 34020 12862
rect 33964 12738 34020 12796
rect 33964 12686 33966 12738
rect 34018 12686 34020 12738
rect 33964 12674 34020 12686
rect 33628 12350 33630 12402
rect 33682 12350 33684 12402
rect 33628 12338 33684 12350
rect 33740 12460 33908 12516
rect 33516 11676 33684 11732
rect 33516 11508 33572 11518
rect 33292 11342 33294 11394
rect 33346 11342 33348 11394
rect 33292 11330 33348 11342
rect 33404 11506 33572 11508
rect 33404 11454 33518 11506
rect 33570 11454 33572 11506
rect 33404 11452 33572 11454
rect 33404 11396 33460 11452
rect 33516 11442 33572 11452
rect 33628 11508 33684 11676
rect 33404 11330 33460 11340
rect 33068 10782 33070 10834
rect 33122 10782 33124 10834
rect 33068 10770 33124 10782
rect 33404 10612 33460 10622
rect 33404 10518 33460 10556
rect 33628 10386 33684 11452
rect 33740 10500 33796 12460
rect 33852 12290 33908 12302
rect 33852 12238 33854 12290
rect 33906 12238 33908 12290
rect 33852 11956 33908 12238
rect 33852 11890 33908 11900
rect 33964 12178 34020 12190
rect 33964 12126 33966 12178
rect 34018 12126 34020 12178
rect 33964 12068 34020 12126
rect 33964 11732 34020 12012
rect 33740 10434 33796 10444
rect 33852 11676 34020 11732
rect 34076 11732 34132 14252
rect 34188 13636 34244 13646
rect 34188 13542 34244 13580
rect 34300 11788 34356 14812
rect 34860 14756 34916 17612
rect 34972 17444 35028 17454
rect 34972 16210 35028 17388
rect 35084 17332 35140 17342
rect 35084 17108 35140 17276
rect 35084 17106 35252 17108
rect 35084 17054 35086 17106
rect 35138 17054 35252 17106
rect 35084 17052 35252 17054
rect 35084 17042 35140 17052
rect 35196 16212 35252 17052
rect 35308 16212 35364 16222
rect 34972 16158 34974 16210
rect 35026 16158 35028 16210
rect 34972 16146 35028 16158
rect 35084 16210 35364 16212
rect 35084 16158 35310 16210
rect 35362 16158 35364 16210
rect 35084 16156 35364 16158
rect 34524 14700 34916 14756
rect 34524 14084 34580 14700
rect 35084 14644 35140 16156
rect 35308 16146 35364 16156
rect 35420 15988 35476 17612
rect 35532 17574 35588 17612
rect 35756 17666 36372 17668
rect 35756 17614 36318 17666
rect 36370 17614 36372 17666
rect 35756 17612 36372 17614
rect 35644 17556 35700 17566
rect 35644 17106 35700 17500
rect 35644 17054 35646 17106
rect 35698 17054 35700 17106
rect 35644 17042 35700 17054
rect 35756 16100 35812 17612
rect 36316 17602 36372 17612
rect 35868 17442 35924 17454
rect 35868 17390 35870 17442
rect 35922 17390 35924 17442
rect 35868 17108 35924 17390
rect 35868 17042 35924 17052
rect 36092 17442 36148 17454
rect 36092 17390 36094 17442
rect 36146 17390 36148 17442
rect 35980 16994 36036 17006
rect 35980 16942 35982 16994
rect 36034 16942 36036 16994
rect 35308 15932 35476 15988
rect 35532 16044 35812 16100
rect 35868 16882 35924 16894
rect 35868 16830 35870 16882
rect 35922 16830 35924 16882
rect 35308 15652 35364 15932
rect 35196 15596 35364 15652
rect 35196 15204 35252 15596
rect 35308 15428 35364 15438
rect 35532 15428 35588 16044
rect 35868 15988 35924 16830
rect 35980 16660 36036 16942
rect 35980 16594 36036 16604
rect 36092 16212 36148 17390
rect 36204 16884 36260 16894
rect 36204 16790 36260 16828
rect 36428 16882 36484 16894
rect 36428 16830 36430 16882
rect 36482 16830 36484 16882
rect 36428 16772 36484 16830
rect 36652 16884 36708 16894
rect 36652 16790 36708 16828
rect 36316 16324 36372 16334
rect 36092 16146 36148 16156
rect 36204 16268 36316 16324
rect 36204 16098 36260 16268
rect 36316 16258 36372 16268
rect 36204 16046 36206 16098
rect 36258 16046 36260 16098
rect 36204 15988 36260 16046
rect 36428 16100 36484 16716
rect 36428 16034 36484 16044
rect 35756 15932 36260 15988
rect 36540 15988 36596 15998
rect 35756 15876 35812 15932
rect 36540 15894 36596 15932
rect 35308 15426 35588 15428
rect 35308 15374 35310 15426
rect 35362 15374 35588 15426
rect 35308 15372 35588 15374
rect 35308 15362 35364 15372
rect 35196 15148 35364 15204
rect 34860 14588 35140 14644
rect 34860 14418 34916 14588
rect 34860 14366 34862 14418
rect 34914 14366 34916 14418
rect 34860 14354 34916 14366
rect 34972 14420 35028 14430
rect 34972 14326 35028 14364
rect 34636 14308 34692 14318
rect 34636 14214 34692 14252
rect 34524 14028 34692 14084
rect 34412 13972 34468 13982
rect 34412 13636 34468 13916
rect 34524 13636 34580 13646
rect 34412 13634 34580 13636
rect 34412 13582 34526 13634
rect 34578 13582 34580 13634
rect 34412 13580 34580 13582
rect 34524 13570 34580 13580
rect 34412 12068 34468 12078
rect 34412 11974 34468 12012
rect 34300 11732 34468 11788
rect 33628 10334 33630 10386
rect 33682 10334 33684 10386
rect 33628 10322 33684 10334
rect 33180 10276 33236 10286
rect 33516 10276 33572 10286
rect 33236 10220 33460 10276
rect 33180 10210 33236 10220
rect 32620 9938 33124 9940
rect 32620 9886 32622 9938
rect 32674 9886 33124 9938
rect 32620 9884 33124 9886
rect 32060 9774 32062 9826
rect 32114 9774 32116 9826
rect 32060 9762 32116 9774
rect 32620 9380 32676 9884
rect 33068 9714 33124 9884
rect 33068 9662 33070 9714
rect 33122 9662 33124 9714
rect 33068 9650 33124 9662
rect 33180 9716 33236 9726
rect 33180 9714 33348 9716
rect 33180 9662 33182 9714
rect 33234 9662 33348 9714
rect 33180 9660 33348 9662
rect 33180 9650 33236 9660
rect 32284 9324 32676 9380
rect 32844 9602 32900 9614
rect 32844 9550 32846 9602
rect 32898 9550 32900 9602
rect 32172 9156 32228 9166
rect 31948 9100 32172 9156
rect 32172 9062 32228 9100
rect 31724 8990 31726 9042
rect 31778 8990 31780 9042
rect 31724 8978 31780 8990
rect 31500 8932 31556 8942
rect 32284 8932 32340 9324
rect 32844 9268 32900 9550
rect 32844 9202 32900 9212
rect 33180 9492 33236 9502
rect 30940 8036 30996 8046
rect 30940 7942 30996 7980
rect 30828 7646 30830 7698
rect 30882 7646 30884 7698
rect 30828 7634 30884 7646
rect 29596 7298 29652 7308
rect 29820 7474 29876 7486
rect 29820 7422 29822 7474
rect 29874 7422 29876 7474
rect 29148 6850 29204 6860
rect 29820 6692 29876 7422
rect 30380 7474 30436 7532
rect 30940 7588 30996 7598
rect 31052 7588 31108 8428
rect 31276 8596 31332 8606
rect 31276 8146 31332 8540
rect 31276 8094 31278 8146
rect 31330 8094 31332 8146
rect 31276 8082 31332 8094
rect 31276 7588 31332 7598
rect 31052 7586 31332 7588
rect 31052 7534 31278 7586
rect 31330 7534 31332 7586
rect 31052 7532 31332 7534
rect 30940 7494 30996 7532
rect 31276 7522 31332 7532
rect 30380 7422 30382 7474
rect 30434 7422 30436 7474
rect 30380 7410 30436 7422
rect 31388 7476 31444 7486
rect 31052 7364 31108 7374
rect 30828 7252 30884 7262
rect 30716 7250 30884 7252
rect 30716 7198 30830 7250
rect 30882 7198 30884 7250
rect 30716 7196 30884 7198
rect 30044 7028 30100 7038
rect 30100 6972 30212 7028
rect 30044 6962 30100 6972
rect 29820 6626 29876 6636
rect 29148 6580 29204 6590
rect 29148 6486 29204 6524
rect 29708 6468 29764 6478
rect 29708 6374 29764 6412
rect 29825 6300 30089 6310
rect 29881 6244 29929 6300
rect 29985 6244 30033 6300
rect 29825 6234 30089 6244
rect 28812 5966 28814 6018
rect 28866 5966 28868 6018
rect 28812 5684 28868 5966
rect 29708 6132 29764 6142
rect 28924 5908 28980 5918
rect 28924 5814 28980 5852
rect 29708 5906 29764 6076
rect 29708 5854 29710 5906
rect 29762 5854 29764 5906
rect 29708 5842 29764 5854
rect 28812 5628 29092 5684
rect 28588 5236 28644 5246
rect 28364 5124 28420 5134
rect 28364 5122 28532 5124
rect 28364 5070 28366 5122
rect 28418 5070 28532 5122
rect 28364 5068 28532 5070
rect 28364 5058 28420 5068
rect 28364 4788 28420 4798
rect 27804 4452 27860 4462
rect 27804 4338 27860 4396
rect 27804 4286 27806 4338
rect 27858 4286 27860 4338
rect 27804 4274 27860 4286
rect 27692 4050 27748 4060
rect 27916 4228 27972 4238
rect 27804 3668 27860 3678
rect 27916 3668 27972 4172
rect 27804 3666 27972 3668
rect 27804 3614 27806 3666
rect 27858 3614 27972 3666
rect 27804 3612 27972 3614
rect 27804 3602 27860 3612
rect 25900 2818 25956 2828
rect 27356 3556 27412 3566
rect 22316 1820 22484 1876
rect 22428 800 22484 1820
rect 27356 800 27412 3500
rect 28364 3554 28420 4732
rect 28476 4226 28532 5068
rect 28588 5010 28644 5180
rect 28588 4958 28590 5010
rect 28642 4958 28644 5010
rect 28588 4946 28644 4958
rect 28812 4564 28868 4574
rect 28812 4450 28868 4508
rect 28812 4398 28814 4450
rect 28866 4398 28868 4450
rect 28812 4386 28868 4398
rect 28476 4174 28478 4226
rect 28530 4174 28532 4226
rect 28476 3780 28532 4174
rect 28924 4338 28980 4350
rect 28924 4286 28926 4338
rect 28978 4286 28980 4338
rect 28476 3714 28532 3724
rect 28588 4116 28644 4126
rect 28588 3778 28644 4060
rect 28588 3726 28590 3778
rect 28642 3726 28644 3778
rect 28588 3714 28644 3726
rect 28924 3778 28980 4286
rect 28924 3726 28926 3778
rect 28978 3726 28980 3778
rect 28364 3502 28366 3554
rect 28418 3502 28420 3554
rect 28364 3490 28420 3502
rect 28924 3332 28980 3726
rect 29036 3780 29092 5628
rect 29708 5572 29764 5582
rect 29260 5460 29316 5470
rect 29260 5346 29316 5404
rect 29260 5294 29262 5346
rect 29314 5294 29316 5346
rect 29260 5282 29316 5294
rect 29596 5348 29652 5358
rect 29596 5254 29652 5292
rect 29372 5122 29428 5134
rect 29372 5070 29374 5122
rect 29426 5070 29428 5122
rect 29372 4788 29428 5070
rect 29372 4722 29428 4732
rect 29484 4450 29540 4462
rect 29484 4398 29486 4450
rect 29538 4398 29540 4450
rect 29484 4116 29540 4398
rect 29708 4116 29764 5516
rect 30156 5234 30212 6972
rect 30156 5182 30158 5234
rect 30210 5182 30212 5234
rect 30156 5170 30212 5182
rect 30380 6020 30436 6030
rect 29825 4732 30089 4742
rect 29881 4676 29929 4732
rect 29985 4676 30033 4732
rect 29825 4666 30089 4676
rect 30380 4564 30436 5964
rect 30604 6020 30660 6030
rect 30604 5346 30660 5964
rect 30604 5294 30606 5346
rect 30658 5294 30660 5346
rect 30604 5282 30660 5294
rect 30492 5012 30548 5022
rect 30492 5010 30660 5012
rect 30492 4958 30494 5010
rect 30546 4958 30660 5010
rect 30492 4956 30660 4958
rect 30492 4946 30548 4956
rect 30380 4498 30436 4508
rect 30604 4452 30660 4956
rect 30604 4358 30660 4396
rect 29820 4340 29876 4350
rect 30716 4340 30772 7196
rect 30828 7186 30884 7196
rect 31052 6690 31108 7308
rect 31052 6638 31054 6690
rect 31106 6638 31108 6690
rect 31052 6626 31108 6638
rect 31276 6692 31332 6702
rect 31388 6692 31444 7420
rect 31276 6690 31444 6692
rect 31276 6638 31278 6690
rect 31330 6638 31444 6690
rect 31276 6636 31444 6638
rect 30828 6580 30884 6590
rect 30828 6486 30884 6524
rect 31164 6578 31220 6590
rect 31164 6526 31166 6578
rect 31218 6526 31220 6578
rect 31164 6468 31220 6526
rect 31164 6402 31220 6412
rect 31052 5796 31108 5806
rect 31052 5702 31108 5740
rect 31276 5122 31332 6636
rect 31388 6356 31444 6366
rect 31388 5906 31444 6300
rect 31388 5854 31390 5906
rect 31442 5854 31444 5906
rect 31388 5842 31444 5854
rect 31276 5070 31278 5122
rect 31330 5070 31332 5122
rect 31276 5058 31332 5070
rect 31500 5122 31556 8876
rect 31948 8876 32340 8932
rect 32508 9042 32564 9054
rect 32508 8990 32510 9042
rect 32562 8990 32564 9042
rect 31948 8258 32004 8876
rect 31948 8206 31950 8258
rect 32002 8206 32004 8258
rect 31948 8194 32004 8206
rect 32060 8148 32116 8158
rect 31612 8036 31668 8046
rect 31612 7140 31668 7980
rect 32060 7140 32116 8092
rect 32172 8146 32228 8158
rect 32172 8094 32174 8146
rect 32226 8094 32228 8146
rect 32172 7700 32228 8094
rect 32508 7700 32564 8990
rect 33180 9042 33236 9436
rect 33180 8990 33182 9042
rect 33234 8990 33236 9042
rect 33180 8978 33236 8990
rect 32732 8258 32788 8270
rect 32732 8206 32734 8258
rect 32786 8206 32788 8258
rect 32732 8148 32788 8206
rect 33180 8260 33236 8270
rect 33180 8166 33236 8204
rect 32732 8082 32788 8092
rect 33292 7700 33348 9660
rect 33404 8372 33460 10220
rect 33516 9492 33572 10220
rect 33516 9426 33572 9436
rect 33628 9828 33684 9838
rect 33516 8484 33572 8494
rect 33628 8484 33684 9772
rect 33516 8482 33684 8484
rect 33516 8430 33518 8482
rect 33570 8430 33684 8482
rect 33516 8428 33684 8430
rect 33740 9042 33796 9054
rect 33740 8990 33742 9042
rect 33794 8990 33796 9042
rect 33740 8596 33796 8990
rect 33516 8418 33572 8428
rect 33740 8372 33796 8540
rect 33404 8306 33460 8316
rect 33628 8316 33796 8372
rect 33628 8036 33684 8316
rect 33852 8260 33908 11676
rect 34076 11666 34132 11676
rect 34412 11396 34468 11732
rect 34636 11508 34692 14028
rect 35084 13970 35140 14588
rect 35084 13918 35086 13970
rect 35138 13918 35140 13970
rect 35084 13906 35140 13918
rect 35196 14420 35252 14430
rect 34860 13074 34916 13086
rect 34860 13022 34862 13074
rect 34914 13022 34916 13074
rect 34860 12964 34916 13022
rect 34860 12898 34916 12908
rect 34972 12962 35028 12974
rect 34972 12910 34974 12962
rect 35026 12910 35028 12962
rect 34972 12852 35028 12910
rect 34972 12786 35028 12796
rect 34860 12628 34916 12638
rect 34916 12572 35028 12628
rect 34860 12562 34916 12572
rect 34860 12068 34916 12078
rect 34860 11974 34916 12012
rect 34972 11844 35028 12572
rect 34860 11788 35028 11844
rect 34636 11452 34804 11508
rect 34076 11340 34468 11396
rect 34524 11394 34580 11406
rect 34524 11342 34526 11394
rect 34578 11342 34580 11394
rect 33964 11282 34020 11294
rect 33964 11230 33966 11282
rect 34018 11230 34020 11282
rect 33964 10724 34020 11230
rect 34076 10724 34132 11340
rect 34300 11172 34356 11182
rect 34300 11078 34356 11116
rect 34524 11060 34580 11342
rect 34524 10994 34580 11004
rect 34076 10668 34244 10724
rect 33964 10658 34020 10668
rect 33964 10498 34020 10510
rect 33964 10446 33966 10498
rect 34018 10446 34020 10498
rect 33964 10386 34020 10446
rect 33964 10334 33966 10386
rect 34018 10334 34020 10386
rect 33964 10322 34020 10334
rect 34076 10388 34132 10398
rect 34076 9826 34132 10332
rect 34188 9938 34244 10668
rect 34300 10612 34356 10622
rect 34300 10518 34356 10556
rect 34188 9886 34190 9938
rect 34242 9886 34244 9938
rect 34188 9874 34244 9886
rect 34300 10052 34356 10062
rect 34076 9774 34078 9826
rect 34130 9774 34132 9826
rect 34076 9762 34132 9774
rect 34300 9826 34356 9996
rect 34300 9774 34302 9826
rect 34354 9774 34356 9826
rect 34300 9762 34356 9774
rect 34524 9044 34580 9054
rect 34524 9042 34692 9044
rect 34524 8990 34526 9042
rect 34578 8990 34692 9042
rect 34524 8988 34692 8990
rect 34524 8978 34580 8988
rect 34636 8932 34692 8988
rect 34748 8932 34804 11452
rect 34860 11396 34916 11788
rect 34860 10610 34916 11340
rect 35084 10612 35140 10622
rect 34860 10558 34862 10610
rect 34914 10558 34916 10610
rect 34860 10546 34916 10558
rect 34972 10610 35140 10612
rect 34972 10558 35086 10610
rect 35138 10558 35140 10610
rect 34972 10556 35140 10558
rect 34860 10052 34916 10062
rect 34972 10052 35028 10556
rect 35084 10546 35140 10556
rect 34916 9996 35028 10052
rect 35084 10388 35140 10398
rect 34860 9938 34916 9996
rect 34860 9886 34862 9938
rect 34914 9886 34916 9938
rect 34860 9874 34916 9886
rect 35084 9826 35140 10332
rect 35084 9774 35086 9826
rect 35138 9774 35140 9826
rect 35084 9762 35140 9774
rect 35196 9268 35252 14364
rect 35308 11172 35364 15148
rect 35532 14530 35588 15372
rect 35644 15874 35812 15876
rect 35644 15822 35758 15874
rect 35810 15822 35812 15874
rect 35644 15820 35812 15822
rect 35644 14980 35700 15820
rect 35756 15810 35812 15820
rect 36316 15874 36372 15886
rect 36316 15822 36318 15874
rect 36370 15822 36372 15874
rect 36316 15652 36372 15822
rect 36204 15596 36372 15652
rect 35644 14914 35700 14924
rect 35756 15540 35812 15550
rect 35756 15428 35812 15484
rect 35980 15428 36036 15438
rect 35756 15426 36036 15428
rect 35756 15374 35982 15426
rect 36034 15374 36036 15426
rect 35756 15372 36036 15374
rect 35532 14478 35534 14530
rect 35586 14478 35588 14530
rect 35532 14466 35588 14478
rect 35644 14642 35700 14654
rect 35644 14590 35646 14642
rect 35698 14590 35700 14642
rect 35644 14308 35700 14590
rect 35644 14242 35700 14252
rect 35420 14084 35476 14094
rect 35476 14028 35588 14084
rect 35420 14018 35476 14028
rect 35308 11106 35364 11116
rect 35420 13860 35476 13870
rect 35420 11060 35476 13804
rect 35420 10994 35476 11004
rect 35308 10722 35364 10734
rect 35308 10670 35310 10722
rect 35362 10670 35364 10722
rect 35308 9828 35364 10670
rect 35420 10610 35476 10622
rect 35420 10558 35422 10610
rect 35474 10558 35476 10610
rect 35420 10164 35476 10558
rect 35420 10098 35476 10108
rect 35308 9762 35364 9772
rect 34860 8932 34916 8942
rect 34748 8876 34860 8932
rect 33852 8194 33908 8204
rect 34300 8372 34356 8382
rect 33516 7700 33572 7710
rect 32172 7644 33460 7700
rect 32284 7476 32340 7486
rect 32284 7362 32340 7420
rect 32284 7310 32286 7362
rect 32338 7310 32340 7362
rect 32284 7298 32340 7310
rect 32732 7252 32788 7262
rect 32060 7084 32452 7140
rect 31612 7074 31668 7084
rect 31612 6578 31668 6590
rect 31612 6526 31614 6578
rect 31666 6526 31668 6578
rect 31612 5236 31668 6526
rect 31612 5170 31668 5180
rect 31724 6580 31780 6590
rect 31724 5236 31780 6524
rect 31948 6580 32004 6590
rect 32284 6580 32340 6590
rect 31948 6578 32340 6580
rect 31948 6526 31950 6578
rect 32002 6526 32286 6578
rect 32338 6526 32340 6578
rect 31948 6524 32340 6526
rect 31948 6514 32004 6524
rect 32284 6514 32340 6524
rect 32396 6578 32452 7084
rect 32620 6804 32676 6814
rect 32396 6526 32398 6578
rect 32450 6526 32452 6578
rect 32396 6514 32452 6526
rect 32508 6692 32564 6702
rect 32396 6130 32452 6142
rect 32396 6078 32398 6130
rect 32450 6078 32452 6130
rect 31836 6020 31892 6030
rect 31836 5926 31892 5964
rect 32284 5906 32340 5918
rect 32284 5854 32286 5906
rect 32338 5854 32340 5906
rect 31724 5234 32004 5236
rect 31724 5182 31726 5234
rect 31778 5182 32004 5234
rect 31724 5180 32004 5182
rect 31724 5170 31780 5180
rect 31500 5070 31502 5122
rect 31554 5070 31556 5122
rect 31500 5058 31556 5070
rect 30940 4340 30996 4350
rect 30716 4338 30996 4340
rect 30716 4286 30942 4338
rect 30994 4286 30996 4338
rect 30716 4284 30996 4286
rect 29820 4246 29876 4284
rect 30940 4274 30996 4284
rect 31948 4338 32004 5180
rect 32284 5122 32340 5854
rect 32396 5348 32452 6078
rect 32396 5282 32452 5292
rect 32284 5070 32286 5122
rect 32338 5070 32340 5122
rect 32284 5058 32340 5070
rect 32508 5122 32564 6636
rect 32620 6690 32676 6748
rect 32620 6638 32622 6690
rect 32674 6638 32676 6690
rect 32620 6626 32676 6638
rect 32620 5348 32676 5358
rect 32732 5348 32788 7196
rect 33180 7140 33236 7150
rect 32956 6692 33012 6702
rect 33012 6636 33124 6692
rect 32956 6626 33012 6636
rect 32844 6580 32900 6590
rect 32844 6486 32900 6524
rect 33068 6132 33124 6636
rect 33180 6356 33236 7084
rect 33292 6692 33348 6702
rect 33292 6578 33348 6636
rect 33292 6526 33294 6578
rect 33346 6526 33348 6578
rect 33292 6514 33348 6526
rect 33404 6690 33460 7644
rect 33516 7474 33572 7644
rect 33516 7422 33518 7474
rect 33570 7422 33572 7474
rect 33516 7410 33572 7422
rect 33404 6638 33406 6690
rect 33458 6638 33460 6690
rect 33404 6468 33460 6638
rect 33628 6692 33684 7980
rect 33740 8146 33796 8158
rect 33740 8094 33742 8146
rect 33794 8094 33796 8146
rect 33740 7476 33796 8094
rect 34188 8148 34244 8158
rect 34188 7586 34244 8092
rect 34188 7534 34190 7586
rect 34242 7534 34244 7586
rect 34188 7522 34244 7534
rect 33740 7382 33796 7420
rect 33852 7364 33908 7374
rect 33852 7270 33908 7308
rect 34300 7028 34356 8316
rect 34300 6916 34356 6972
rect 33628 6626 33684 6636
rect 33964 6860 34356 6916
rect 34524 7812 34580 7822
rect 34524 7698 34580 7756
rect 34524 7646 34526 7698
rect 34578 7646 34580 7698
rect 33964 6690 34020 6860
rect 33964 6638 33966 6690
rect 34018 6638 34020 6690
rect 33964 6626 34020 6638
rect 34300 6692 34356 6702
rect 34300 6598 34356 6636
rect 33404 6412 33572 6468
rect 33180 6300 33348 6356
rect 33180 6132 33236 6142
rect 33068 6130 33236 6132
rect 33068 6078 33182 6130
rect 33234 6078 33236 6130
rect 33068 6076 33236 6078
rect 33180 6066 33236 6076
rect 32956 5908 33012 5918
rect 32956 5814 33012 5852
rect 33292 5908 33348 6300
rect 33292 5906 33460 5908
rect 33292 5854 33294 5906
rect 33346 5854 33460 5906
rect 33292 5852 33460 5854
rect 33292 5842 33348 5852
rect 32620 5346 32788 5348
rect 32620 5294 32622 5346
rect 32674 5294 32788 5346
rect 32620 5292 32788 5294
rect 32620 5282 32676 5292
rect 32508 5070 32510 5122
rect 32562 5070 32564 5122
rect 32508 5058 32564 5070
rect 33068 5236 33124 5246
rect 33068 5122 33124 5180
rect 33068 5070 33070 5122
rect 33122 5070 33124 5122
rect 33068 5058 33124 5070
rect 31948 4286 31950 4338
rect 32002 4286 32004 4338
rect 31948 4274 32004 4286
rect 32396 4900 32452 4910
rect 29932 4228 29988 4238
rect 29932 4134 29988 4172
rect 29708 4060 29876 4116
rect 29484 4050 29540 4060
rect 29372 3780 29428 3790
rect 29036 3778 29428 3780
rect 29036 3726 29374 3778
rect 29426 3726 29428 3778
rect 29036 3724 29428 3726
rect 29372 3714 29428 3724
rect 29708 3780 29764 3790
rect 29820 3780 29876 4060
rect 29932 3780 29988 3790
rect 29820 3724 29932 3780
rect 29708 3686 29764 3724
rect 29932 3666 29988 3724
rect 29932 3614 29934 3666
rect 29986 3614 29988 3666
rect 29932 3602 29988 3614
rect 30604 3556 30660 3566
rect 30604 3462 30660 3500
rect 30940 3444 30996 3482
rect 30940 3378 30996 3388
rect 31276 3442 31332 3454
rect 31276 3390 31278 3442
rect 31330 3390 31332 3442
rect 28924 2324 28980 3276
rect 30268 3330 30324 3342
rect 30268 3278 30270 3330
rect 30322 3278 30324 3330
rect 29825 3164 30089 3174
rect 29881 3108 29929 3164
rect 29985 3108 30033 3164
rect 29825 3098 30089 3108
rect 30268 2996 30324 3278
rect 30268 2930 30324 2940
rect 31276 2436 31332 3390
rect 32396 3444 32452 4844
rect 32620 4898 32676 4910
rect 32620 4846 32622 4898
rect 32674 4846 32676 4898
rect 32620 4564 32676 4846
rect 32620 4498 32676 4508
rect 33292 4340 33348 4350
rect 32508 4228 32564 4238
rect 32508 4134 32564 4172
rect 33292 3668 33348 4284
rect 33292 3602 33348 3612
rect 33404 3666 33460 5852
rect 33516 5234 33572 6412
rect 34076 6466 34132 6478
rect 34076 6414 34078 6466
rect 34130 6414 34132 6466
rect 33964 6020 34020 6030
rect 34076 6020 34132 6414
rect 34188 6020 34244 6030
rect 34524 6020 34580 7646
rect 34076 6018 34244 6020
rect 34076 5966 34190 6018
rect 34242 5966 34244 6018
rect 34076 5964 34244 5966
rect 33964 5926 34020 5964
rect 33516 5182 33518 5234
rect 33570 5182 33572 5234
rect 33516 5170 33572 5182
rect 33852 5908 33908 5918
rect 33852 5124 33908 5852
rect 34076 5684 34132 5694
rect 33964 5124 34020 5134
rect 33852 5122 34020 5124
rect 33852 5070 33966 5122
rect 34018 5070 34020 5122
rect 33852 5068 34020 5070
rect 33964 5058 34020 5068
rect 33628 4900 33684 4910
rect 34076 4900 34132 5628
rect 34188 5124 34244 5964
rect 34412 5964 34524 6020
rect 34300 5906 34356 5918
rect 34300 5854 34302 5906
rect 34354 5854 34356 5906
rect 34300 5684 34356 5854
rect 34300 5618 34356 5628
rect 34188 5068 34356 5124
rect 34188 4900 34244 4910
rect 34076 4898 34244 4900
rect 34076 4846 34190 4898
rect 34242 4846 34244 4898
rect 34076 4844 34244 4846
rect 33628 4562 33684 4844
rect 34188 4834 34244 4844
rect 33628 4510 33630 4562
rect 33682 4510 33684 4562
rect 33628 4498 33684 4510
rect 34076 4564 34132 4574
rect 34076 4470 34132 4508
rect 33852 4452 33908 4462
rect 33852 4358 33908 4396
rect 34188 4340 34244 4350
rect 34300 4340 34356 5068
rect 34412 5122 34468 5964
rect 34524 5954 34580 5964
rect 34524 5236 34580 5246
rect 34524 5142 34580 5180
rect 34412 5070 34414 5122
rect 34466 5070 34468 5122
rect 34412 5058 34468 5070
rect 34524 4900 34580 4910
rect 34636 4900 34692 8876
rect 34860 8838 34916 8876
rect 34748 8372 34804 8382
rect 34748 8278 34804 8316
rect 35196 8146 35252 9212
rect 35532 9156 35588 14028
rect 35644 13972 35700 13982
rect 35756 13972 35812 15372
rect 35980 15362 36036 15372
rect 36204 14644 36260 15596
rect 36316 15428 36372 15438
rect 36764 15428 36820 18172
rect 36988 18162 37044 18172
rect 36979 18060 37243 18070
rect 37035 18004 37083 18060
rect 37139 18004 37187 18060
rect 36979 17994 37243 18004
rect 37100 17780 37156 17790
rect 37100 17686 37156 17724
rect 37324 17780 37380 18172
rect 37324 17714 37380 17724
rect 37548 18004 37604 18014
rect 37548 17666 37604 17948
rect 37548 17614 37550 17666
rect 37602 17614 37604 17666
rect 36876 16884 36932 16894
rect 36876 16790 36932 16828
rect 37100 16882 37156 16894
rect 37100 16830 37102 16882
rect 37154 16830 37156 16882
rect 37100 16660 37156 16830
rect 37436 16884 37492 16894
rect 37548 16884 37604 17614
rect 37436 16882 37604 16884
rect 37436 16830 37438 16882
rect 37490 16830 37604 16882
rect 37436 16828 37604 16830
rect 37436 16818 37492 16828
rect 37660 16660 37716 19180
rect 37772 19124 37828 19134
rect 37884 19124 37940 20076
rect 38220 20018 38276 20030
rect 38220 19966 38222 20018
rect 38274 19966 38276 20018
rect 38220 19796 38276 19966
rect 38444 20020 38500 20030
rect 38444 19926 38500 19964
rect 38556 19796 38612 20300
rect 38220 19740 38612 19796
rect 38556 19572 38612 19740
rect 38668 20130 38724 20142
rect 38668 20078 38670 20130
rect 38722 20078 38724 20130
rect 38668 19684 38724 20078
rect 38668 19618 38724 19628
rect 38780 20020 38836 20030
rect 38892 20020 38948 24668
rect 39004 24276 39060 25676
rect 39116 25620 39172 25900
rect 39340 26066 39396 26078
rect 39340 26014 39342 26066
rect 39394 26014 39396 26066
rect 39340 25732 39396 26014
rect 39340 25666 39396 25676
rect 39116 25554 39172 25564
rect 39452 25618 39508 25630
rect 39452 25566 39454 25618
rect 39506 25566 39508 25618
rect 39452 25508 39508 25566
rect 39452 25442 39508 25452
rect 39116 25282 39172 25294
rect 39116 25230 39118 25282
rect 39170 25230 39172 25282
rect 39116 24722 39172 25230
rect 39228 24836 39284 24874
rect 39228 24770 39284 24780
rect 39116 24670 39118 24722
rect 39170 24670 39172 24722
rect 39116 24658 39172 24670
rect 39564 24610 39620 27692
rect 40012 27682 40068 27692
rect 40012 27188 40068 27198
rect 40124 27188 40180 30828
rect 40348 30818 40404 30828
rect 40684 30324 40740 30334
rect 41020 30324 41076 31388
rect 41468 30884 41524 30894
rect 40684 30322 41076 30324
rect 40684 30270 40686 30322
rect 40738 30270 41076 30322
rect 40684 30268 41076 30270
rect 41244 30772 41300 30782
rect 40684 30258 40740 30268
rect 40348 29316 40404 29326
rect 40236 29314 40404 29316
rect 40236 29262 40350 29314
rect 40402 29262 40404 29314
rect 40236 29260 40404 29262
rect 40236 27972 40292 29260
rect 40348 29250 40404 29260
rect 41244 28980 41300 30716
rect 41468 30324 41524 30828
rect 41468 30258 41524 30268
rect 41244 28914 41300 28924
rect 40796 28756 40852 28766
rect 40796 28642 40852 28700
rect 40796 28590 40798 28642
rect 40850 28590 40852 28642
rect 40796 28578 40852 28590
rect 41580 28644 41636 28654
rect 41580 28550 41636 28588
rect 40684 28532 40740 28542
rect 40684 28438 40740 28476
rect 41244 28532 41300 28542
rect 41020 28084 41076 28094
rect 41020 27990 41076 28028
rect 40236 27906 40292 27916
rect 40908 27972 40964 27982
rect 40908 27878 40964 27916
rect 41244 27972 41300 28476
rect 41244 27858 41300 27916
rect 41244 27806 41246 27858
rect 41298 27806 41300 27858
rect 41244 27794 41300 27806
rect 39676 27132 39956 27188
rect 39676 27074 39732 27132
rect 39676 27022 39678 27074
rect 39730 27022 39732 27074
rect 39676 27010 39732 27022
rect 39788 26962 39844 26974
rect 39788 26910 39790 26962
rect 39842 26910 39844 26962
rect 39676 26516 39732 26526
rect 39788 26516 39844 26910
rect 39676 26514 39844 26516
rect 39676 26462 39678 26514
rect 39730 26462 39844 26514
rect 39676 26460 39844 26462
rect 39676 25506 39732 26460
rect 39900 26180 39956 27132
rect 40012 27186 40180 27188
rect 40012 27134 40014 27186
rect 40066 27134 40180 27186
rect 40012 27132 40180 27134
rect 40012 27122 40068 27132
rect 40124 26962 40180 26974
rect 40124 26910 40126 26962
rect 40178 26910 40180 26962
rect 40124 26908 40180 26910
rect 41804 26908 41860 31612
rect 40124 26852 40852 26908
rect 40796 26514 40852 26852
rect 40796 26462 40798 26514
rect 40850 26462 40852 26514
rect 40796 26450 40852 26462
rect 41580 26852 41860 26908
rect 40124 26404 40180 26414
rect 40012 26180 40068 26190
rect 39900 26178 40068 26180
rect 39900 26126 40014 26178
rect 40066 26126 40068 26178
rect 39900 26124 40068 26126
rect 40012 26114 40068 26124
rect 39676 25454 39678 25506
rect 39730 25454 39732 25506
rect 39676 25442 39732 25454
rect 40012 25508 40068 25518
rect 40124 25508 40180 26348
rect 41020 26404 41076 26414
rect 41020 26310 41076 26348
rect 40348 26292 40404 26302
rect 40348 26198 40404 26236
rect 41132 26292 41188 26302
rect 40068 25452 40180 25508
rect 41132 25506 41188 26236
rect 41132 25454 41134 25506
rect 41186 25454 41188 25506
rect 40012 25442 40068 25452
rect 41132 25442 41188 25454
rect 39564 24558 39566 24610
rect 39618 24558 39620 24610
rect 39564 24546 39620 24558
rect 39788 25396 39844 25406
rect 39116 24276 39172 24286
rect 39004 24220 39116 24276
rect 39116 24210 39172 24220
rect 39004 23828 39060 23838
rect 39004 23734 39060 23772
rect 39788 23716 39844 25340
rect 40572 25172 40628 25182
rect 40012 24722 40068 24734
rect 40012 24670 40014 24722
rect 40066 24670 40068 24722
rect 40012 24612 40068 24670
rect 40012 24546 40068 24556
rect 40572 24050 40628 25116
rect 40572 23998 40574 24050
rect 40626 23998 40628 24050
rect 40572 23986 40628 23998
rect 41244 24724 41300 24734
rect 39900 23940 39956 23950
rect 39900 23846 39956 23884
rect 41244 23938 41300 24668
rect 41244 23886 41246 23938
rect 41298 23886 41300 23938
rect 41244 23874 41300 23886
rect 39676 23604 39732 23614
rect 39564 23380 39620 23390
rect 39228 23154 39284 23166
rect 39228 23102 39230 23154
rect 39282 23102 39284 23154
rect 39228 22596 39284 23102
rect 39564 23156 39620 23324
rect 39676 23266 39732 23548
rect 39676 23214 39678 23266
rect 39730 23214 39732 23266
rect 39676 23202 39732 23214
rect 39564 23090 39620 23100
rect 39228 22260 39284 22540
rect 39676 22484 39732 22494
rect 39228 22194 39284 22204
rect 39452 22258 39508 22270
rect 39452 22206 39454 22258
rect 39506 22206 39508 22258
rect 39004 22148 39060 22158
rect 39004 20132 39060 22092
rect 39116 22146 39172 22158
rect 39116 22094 39118 22146
rect 39170 22094 39172 22146
rect 39116 21586 39172 22094
rect 39340 22146 39396 22158
rect 39340 22094 39342 22146
rect 39394 22094 39396 22146
rect 39340 21700 39396 22094
rect 39116 21534 39118 21586
rect 39170 21534 39172 21586
rect 39116 21522 39172 21534
rect 39228 21644 39396 21700
rect 39228 21588 39284 21644
rect 39228 21252 39284 21532
rect 39452 21588 39508 22206
rect 39676 21812 39732 22428
rect 39676 21746 39732 21756
rect 39788 21810 39844 23660
rect 40908 23826 40964 23838
rect 40908 23774 40910 23826
rect 40962 23774 40964 23826
rect 40908 23604 40964 23774
rect 41468 23826 41524 23838
rect 41468 23774 41470 23826
rect 41522 23774 41524 23826
rect 40908 23538 40964 23548
rect 41020 23714 41076 23726
rect 41020 23662 41022 23714
rect 41074 23662 41076 23714
rect 39900 23380 39956 23390
rect 39900 22482 39956 23324
rect 41020 23044 41076 23662
rect 41468 23492 41524 23774
rect 41244 23436 41524 23492
rect 41244 23044 41300 23436
rect 41020 22988 41300 23044
rect 40460 22932 40516 22942
rect 39900 22430 39902 22482
rect 39954 22430 39956 22482
rect 39900 22372 39956 22430
rect 39900 22306 39956 22316
rect 40236 22708 40292 22718
rect 40236 22148 40292 22652
rect 40236 22082 40292 22092
rect 40460 22258 40516 22876
rect 40460 22206 40462 22258
rect 40514 22206 40516 22258
rect 39788 21758 39790 21810
rect 39842 21758 39844 21810
rect 39788 21746 39844 21758
rect 40348 21700 40404 21710
rect 39452 21522 39508 21532
rect 40124 21588 40180 21598
rect 40124 21494 40180 21532
rect 39340 21476 39396 21486
rect 39340 21382 39396 21420
rect 39228 21196 39396 21252
rect 39228 20132 39284 20142
rect 39004 20130 39284 20132
rect 39004 20078 39230 20130
rect 39282 20078 39284 20130
rect 39004 20076 39284 20078
rect 38892 19964 39172 20020
rect 38556 19506 38612 19516
rect 37996 19348 38052 19358
rect 37996 19254 38052 19292
rect 37884 19068 38052 19124
rect 37772 18674 37828 19068
rect 37772 18622 37774 18674
rect 37826 18622 37828 18674
rect 37772 18610 37828 18622
rect 37884 18676 37940 18686
rect 37884 18562 37940 18620
rect 37884 18510 37886 18562
rect 37938 18510 37940 18562
rect 37884 18498 37940 18510
rect 37100 16604 37380 16660
rect 36979 16492 37243 16502
rect 37035 16436 37083 16492
rect 37139 16436 37187 16492
rect 36979 16426 37243 16436
rect 36988 16100 37044 16110
rect 36988 16006 37044 16044
rect 37212 15988 37268 15998
rect 37212 15894 37268 15932
rect 36316 15426 36820 15428
rect 36316 15374 36318 15426
rect 36370 15374 36820 15426
rect 36316 15372 36820 15374
rect 36316 15362 36372 15372
rect 36764 15314 36820 15372
rect 36764 15262 36766 15314
rect 36818 15262 36820 15314
rect 36764 15250 36820 15262
rect 36979 14924 37243 14934
rect 37035 14868 37083 14924
rect 37139 14868 37187 14924
rect 36979 14858 37243 14868
rect 37324 14756 37380 16604
rect 37436 16604 37716 16660
rect 37436 16100 37492 16604
rect 37660 16100 37716 16110
rect 37436 16044 37604 16100
rect 37436 15874 37492 15886
rect 37436 15822 37438 15874
rect 37490 15822 37492 15874
rect 37436 15426 37492 15822
rect 37436 15374 37438 15426
rect 37490 15374 37492 15426
rect 37436 15362 37492 15374
rect 37324 14690 37380 14700
rect 36204 14578 36260 14588
rect 37100 14532 37156 14542
rect 37100 14438 37156 14476
rect 35644 13970 35812 13972
rect 35644 13918 35646 13970
rect 35698 13918 35812 13970
rect 35644 13916 35812 13918
rect 36428 14418 36484 14430
rect 36428 14366 36430 14418
rect 36482 14366 36484 14418
rect 35644 13906 35700 13916
rect 36428 13860 36484 14366
rect 37548 14084 37604 16044
rect 37660 16098 37940 16100
rect 37660 16046 37662 16098
rect 37714 16046 37940 16098
rect 37660 16044 37940 16046
rect 37660 16034 37716 16044
rect 37884 15540 37940 16044
rect 37660 15484 37940 15540
rect 37660 14532 37716 15484
rect 37660 14466 37716 14476
rect 37324 14028 37604 14084
rect 37324 13970 37380 14028
rect 37324 13918 37326 13970
rect 37378 13918 37380 13970
rect 37324 13906 37380 13918
rect 36428 13766 36484 13804
rect 37436 13860 37492 13870
rect 36764 13746 36820 13758
rect 36764 13694 36766 13746
rect 36818 13694 36820 13746
rect 35644 12850 35700 12862
rect 35644 12798 35646 12850
rect 35698 12798 35700 12850
rect 35644 12180 35700 12798
rect 36764 12404 36820 13694
rect 37324 13746 37380 13758
rect 37324 13694 37326 13746
rect 37378 13694 37380 13746
rect 36979 13356 37243 13366
rect 37035 13300 37083 13356
rect 37139 13300 37187 13356
rect 36979 13290 37243 13300
rect 36764 12348 36932 12404
rect 36876 12292 36932 12348
rect 37324 12402 37380 13694
rect 37436 12962 37492 13804
rect 37436 12910 37438 12962
rect 37490 12910 37492 12962
rect 37436 12898 37492 12910
rect 37660 12964 37716 12974
rect 37324 12350 37326 12402
rect 37378 12350 37380 12402
rect 37324 12338 37380 12350
rect 36988 12292 37044 12302
rect 36876 12290 37044 12292
rect 36876 12238 36990 12290
rect 37042 12238 37044 12290
rect 36876 12236 37044 12238
rect 36988 12226 37044 12236
rect 35644 12114 35700 12124
rect 36316 12178 36372 12190
rect 36316 12126 36318 12178
rect 36370 12126 36372 12178
rect 36316 12068 36372 12126
rect 36764 12180 36820 12190
rect 36764 12086 36820 12124
rect 37660 12180 37716 12908
rect 37660 12086 37716 12124
rect 37884 12962 37940 12974
rect 37884 12910 37886 12962
rect 37938 12910 37940 12962
rect 35756 12012 36316 12068
rect 35756 11618 35812 12012
rect 36316 11974 36372 12012
rect 37884 12068 37940 12910
rect 37884 11974 37940 12012
rect 36979 11788 37243 11798
rect 37035 11732 37083 11788
rect 37139 11732 37187 11788
rect 36979 11722 37243 11732
rect 35756 11566 35758 11618
rect 35810 11566 35812 11618
rect 35756 11554 35812 11566
rect 35868 11508 35924 11518
rect 35868 11506 36484 11508
rect 35868 11454 35870 11506
rect 35922 11454 36484 11506
rect 35868 11452 36484 11454
rect 35868 11442 35924 11452
rect 35756 11394 35812 11406
rect 35756 11342 35758 11394
rect 35810 11342 35812 11394
rect 35756 11284 35812 11342
rect 35644 11228 35756 11284
rect 35644 10050 35700 11228
rect 35756 11218 35812 11228
rect 35756 11060 35812 11070
rect 35812 11004 35924 11060
rect 35756 10994 35812 11004
rect 35868 10836 35924 11004
rect 35868 10834 36260 10836
rect 35868 10782 35870 10834
rect 35922 10782 36260 10834
rect 35868 10780 36260 10782
rect 35868 10770 35924 10780
rect 35756 10610 35812 10622
rect 35756 10558 35758 10610
rect 35810 10558 35812 10610
rect 35756 10500 35812 10558
rect 35756 10434 35812 10444
rect 35868 10388 35924 10398
rect 35868 10294 35924 10332
rect 35644 9998 35646 10050
rect 35698 9998 35700 10050
rect 35644 9986 35700 9998
rect 35756 10052 35812 10062
rect 35756 9156 35812 9996
rect 35420 9100 35588 9156
rect 35644 9100 35812 9156
rect 36204 9938 36260 10780
rect 36428 10834 36484 11452
rect 37100 11506 37156 11518
rect 37100 11454 37102 11506
rect 37154 11454 37156 11506
rect 36540 11396 36596 11406
rect 36540 11394 36932 11396
rect 36540 11342 36542 11394
rect 36594 11342 36932 11394
rect 36540 11340 36932 11342
rect 36540 11330 36596 11340
rect 36428 10782 36430 10834
rect 36482 10782 36484 10834
rect 36428 10770 36484 10782
rect 36876 10834 36932 11340
rect 36876 10782 36878 10834
rect 36930 10782 36932 10834
rect 36876 10770 36932 10782
rect 36316 10724 36372 10734
rect 36316 10630 36372 10668
rect 37100 10722 37156 11454
rect 37996 11508 38052 19068
rect 38780 18676 38836 19964
rect 38836 18620 38948 18676
rect 38780 18582 38836 18620
rect 38332 18452 38388 18462
rect 38332 18338 38388 18396
rect 38332 18286 38334 18338
rect 38386 18286 38388 18338
rect 38108 17780 38164 17790
rect 38164 17724 38276 17780
rect 38108 17714 38164 17724
rect 38220 17666 38276 17724
rect 38220 17614 38222 17666
rect 38274 17614 38276 17666
rect 38220 17602 38276 17614
rect 38108 16884 38164 16894
rect 38108 16790 38164 16828
rect 38220 16324 38276 16334
rect 38108 16212 38164 16222
rect 38108 16118 38164 16156
rect 38220 16100 38276 16268
rect 38220 16034 38276 16044
rect 38332 15148 38388 18286
rect 38668 16996 38724 17006
rect 38724 16940 38836 16996
rect 38668 16930 38724 16940
rect 38444 15876 38500 15886
rect 38668 15876 38724 15886
rect 38444 15874 38612 15876
rect 38444 15822 38446 15874
rect 38498 15822 38612 15874
rect 38444 15820 38612 15822
rect 38444 15810 38500 15820
rect 38332 15092 38500 15148
rect 37996 11442 38052 11452
rect 37324 11284 37380 11294
rect 37324 11190 37380 11228
rect 37100 10670 37102 10722
rect 37154 10670 37156 10722
rect 36652 10612 36708 10622
rect 37100 10612 37156 10670
rect 37212 10724 37268 10734
rect 37212 10630 37268 10668
rect 36652 10610 37156 10612
rect 36652 10558 36654 10610
rect 36706 10558 37156 10610
rect 36652 10556 37156 10558
rect 36652 10546 36708 10556
rect 37100 10388 37156 10556
rect 37100 10332 37380 10388
rect 36979 10220 37243 10230
rect 37035 10164 37083 10220
rect 37139 10164 37187 10220
rect 36979 10154 37243 10164
rect 36204 9886 36206 9938
rect 36258 9886 36260 9938
rect 35420 8372 35476 9100
rect 35644 9044 35700 9100
rect 35532 8932 35588 8942
rect 35644 8932 35700 8988
rect 35532 8930 35700 8932
rect 35532 8878 35534 8930
rect 35586 8878 35700 8930
rect 35532 8876 35700 8878
rect 35756 8930 35812 8942
rect 35756 8878 35758 8930
rect 35810 8878 35812 8930
rect 35532 8866 35588 8876
rect 35756 8484 35812 8878
rect 35980 8820 36036 8830
rect 36204 8820 36260 9886
rect 37324 9154 37380 10332
rect 38332 9602 38388 9614
rect 38332 9550 38334 9602
rect 38386 9550 38388 9602
rect 38332 9380 38388 9550
rect 38332 9314 38388 9324
rect 37324 9102 37326 9154
rect 37378 9102 37380 9154
rect 37324 9090 37380 9102
rect 36316 9044 36372 9054
rect 36764 9044 36820 9054
rect 36316 9042 36820 9044
rect 36316 8990 36318 9042
rect 36370 8990 36766 9042
rect 36818 8990 36820 9042
rect 36316 8988 36820 8990
rect 36316 8978 36372 8988
rect 36764 8978 36820 8988
rect 37212 9042 37268 9054
rect 37212 8990 37214 9042
rect 37266 8990 37268 9042
rect 37212 8820 37268 8990
rect 38108 9042 38164 9054
rect 38108 8990 38110 9042
rect 38162 8990 38164 9042
rect 38108 8932 38164 8990
rect 38332 8932 38388 8942
rect 38108 8930 38388 8932
rect 38108 8878 38334 8930
rect 38386 8878 38388 8930
rect 38108 8876 38388 8878
rect 38332 8866 38388 8876
rect 36204 8764 36484 8820
rect 37212 8764 37380 8820
rect 35980 8726 36036 8764
rect 35980 8484 36036 8494
rect 35756 8482 36036 8484
rect 35756 8430 35982 8482
rect 36034 8430 36036 8482
rect 35756 8428 36036 8430
rect 35420 8306 35476 8316
rect 35980 8372 36036 8428
rect 35980 8306 36036 8316
rect 36092 8260 36148 8270
rect 36092 8166 36148 8204
rect 35980 8148 36036 8158
rect 35196 8094 35198 8146
rect 35250 8094 35252 8146
rect 35196 8082 35252 8094
rect 35868 8146 36036 8148
rect 35868 8094 35982 8146
rect 36034 8094 36036 8146
rect 35868 8092 36036 8094
rect 35532 8036 35588 8046
rect 35308 8034 35588 8036
rect 35308 7982 35534 8034
rect 35586 7982 35588 8034
rect 35308 7980 35588 7982
rect 35308 7700 35364 7980
rect 35532 7812 35588 7980
rect 35868 8036 35924 8092
rect 35980 8082 36036 8092
rect 35868 7970 35924 7980
rect 35980 7868 36372 7924
rect 35980 7812 36036 7868
rect 35532 7756 36036 7812
rect 35196 7644 35364 7700
rect 35420 7700 35476 7710
rect 36092 7700 36148 7710
rect 34972 7362 35028 7374
rect 34972 7310 34974 7362
rect 35026 7310 35028 7362
rect 34972 7140 35028 7310
rect 34972 7074 35028 7084
rect 34748 7028 34804 7038
rect 34748 6356 34804 6972
rect 35084 6804 35140 6814
rect 35084 6710 35140 6748
rect 34860 6692 34916 6702
rect 34916 6636 35028 6692
rect 34860 6598 34916 6636
rect 34748 6300 34916 6356
rect 34748 6132 34804 6142
rect 34748 6038 34804 6076
rect 34860 5572 34916 6300
rect 34972 5796 35028 6636
rect 35084 5796 35140 5806
rect 34972 5794 35140 5796
rect 34972 5742 35086 5794
rect 35138 5742 35140 5794
rect 34972 5740 35140 5742
rect 35084 5730 35140 5740
rect 35196 5684 35252 7644
rect 35420 7606 35476 7644
rect 35532 7698 36148 7700
rect 35532 7646 36094 7698
rect 36146 7646 36148 7698
rect 35532 7644 36148 7646
rect 35308 7474 35364 7486
rect 35308 7422 35310 7474
rect 35362 7422 35364 7474
rect 35308 6916 35364 7422
rect 35532 7474 35588 7644
rect 36092 7634 36148 7644
rect 36316 7698 36372 7868
rect 36316 7646 36318 7698
rect 36370 7646 36372 7698
rect 36316 7634 36372 7646
rect 36428 7812 36484 8764
rect 36979 8652 37243 8662
rect 37035 8596 37083 8652
rect 37139 8596 37187 8652
rect 36979 8586 37243 8596
rect 37212 8260 37268 8270
rect 36428 7586 36484 7756
rect 36428 7534 36430 7586
rect 36482 7534 36484 7586
rect 36428 7522 36484 7534
rect 36876 8148 36932 8158
rect 36876 7588 36932 8092
rect 37212 7700 37268 8204
rect 37324 8148 37380 8764
rect 37772 8372 37828 8382
rect 37772 8258 37828 8316
rect 37772 8206 37774 8258
rect 37826 8206 37828 8258
rect 37772 8194 37828 8206
rect 37436 8148 37492 8158
rect 37324 8146 37492 8148
rect 37324 8094 37438 8146
rect 37490 8094 37492 8146
rect 37324 8092 37492 8094
rect 37324 7700 37380 7710
rect 37212 7698 37380 7700
rect 37212 7646 37326 7698
rect 37378 7646 37380 7698
rect 37212 7644 37380 7646
rect 37324 7634 37380 7644
rect 36876 7494 36932 7532
rect 35532 7422 35534 7474
rect 35586 7422 35588 7474
rect 35420 6916 35476 6926
rect 35308 6914 35476 6916
rect 35308 6862 35422 6914
rect 35474 6862 35476 6914
rect 35308 6860 35476 6862
rect 35420 6850 35476 6860
rect 35532 5906 35588 7422
rect 35980 7476 36036 7486
rect 35980 7474 36260 7476
rect 35980 7422 35982 7474
rect 36034 7422 36260 7474
rect 35980 7420 36260 7422
rect 35980 7410 36036 7420
rect 36204 6916 36260 7420
rect 37436 7252 37492 8092
rect 37772 7812 37828 7822
rect 37772 7698 37828 7756
rect 37772 7646 37774 7698
rect 37826 7646 37828 7698
rect 37772 7634 37828 7646
rect 37436 7186 37492 7196
rect 38220 7476 38276 7486
rect 36979 7084 37243 7094
rect 37035 7028 37083 7084
rect 37139 7028 37187 7084
rect 36979 7018 37243 7028
rect 36316 6916 36372 6926
rect 36204 6914 36372 6916
rect 36204 6862 36318 6914
rect 36370 6862 36372 6914
rect 36204 6860 36372 6862
rect 36316 6850 36372 6860
rect 35980 6804 36036 6814
rect 35980 6710 36036 6748
rect 36540 6804 36596 6814
rect 35756 6692 35812 6702
rect 35756 6598 35812 6636
rect 35532 5854 35534 5906
rect 35586 5854 35588 5906
rect 35532 5842 35588 5854
rect 35644 6132 35700 6142
rect 35196 5618 35252 5628
rect 34860 5516 35140 5572
rect 35084 5234 35140 5516
rect 35084 5182 35086 5234
rect 35138 5182 35140 5234
rect 35084 5170 35140 5182
rect 35532 5236 35588 5246
rect 35644 5236 35700 6076
rect 36540 5906 36596 6748
rect 37548 6578 37604 6590
rect 37548 6526 37550 6578
rect 37602 6526 37604 6578
rect 37324 6020 37380 6030
rect 37324 5926 37380 5964
rect 36540 5854 36542 5906
rect 36594 5854 36596 5906
rect 36540 5842 36596 5854
rect 36979 5516 37243 5526
rect 37035 5460 37083 5516
rect 37139 5460 37187 5516
rect 36979 5450 37243 5460
rect 37100 5348 37156 5358
rect 35532 5234 35700 5236
rect 35532 5182 35534 5234
rect 35586 5182 35700 5234
rect 35532 5180 35700 5182
rect 35756 5236 35812 5246
rect 35532 5170 35588 5180
rect 35756 5142 35812 5180
rect 37100 5234 37156 5292
rect 37100 5182 37102 5234
rect 37154 5182 37156 5234
rect 34580 4844 34692 4900
rect 34972 5124 35028 5134
rect 34524 4806 34580 4844
rect 34244 4284 34356 4340
rect 34636 4564 34692 4574
rect 34972 4564 35028 5068
rect 36092 5012 36148 5022
rect 36092 4898 36148 4956
rect 36092 4846 36094 4898
rect 36146 4846 36148 4898
rect 36092 4834 36148 4846
rect 37100 4676 37156 5182
rect 37548 5012 37604 6526
rect 37660 6468 37716 6478
rect 38108 6468 38164 6478
rect 37660 6466 37828 6468
rect 37660 6414 37662 6466
rect 37714 6414 37828 6466
rect 37660 6412 37828 6414
rect 37660 6402 37716 6412
rect 37548 4918 37604 4956
rect 37100 4610 37156 4620
rect 35084 4564 35140 4574
rect 34972 4562 35140 4564
rect 34972 4510 35086 4562
rect 35138 4510 35140 4562
rect 34972 4508 35140 4510
rect 34188 4246 34244 4284
rect 34636 4226 34692 4508
rect 35084 4498 35140 4508
rect 37772 4452 37828 6412
rect 38108 6130 38164 6412
rect 38108 6078 38110 6130
rect 38162 6078 38164 6130
rect 38108 6066 38164 6078
rect 38220 6130 38276 7420
rect 38220 6078 38222 6130
rect 38274 6078 38276 6130
rect 38220 6066 38276 6078
rect 38332 5684 38388 5694
rect 38332 5590 38388 5628
rect 37772 4386 37828 4396
rect 38332 4676 38388 4686
rect 38220 4338 38276 4350
rect 38220 4286 38222 4338
rect 38274 4286 38276 4338
rect 37884 4228 37940 4238
rect 34636 4174 34638 4226
rect 34690 4174 34692 4226
rect 34636 4004 34692 4174
rect 37660 4226 37940 4228
rect 37660 4174 37886 4226
rect 37938 4174 37940 4226
rect 37660 4172 37940 4174
rect 37324 4116 37380 4126
rect 34636 3938 34692 3948
rect 36979 3948 37243 3958
rect 37035 3892 37083 3948
rect 37139 3892 37187 3948
rect 36979 3882 37243 3892
rect 33404 3614 33406 3666
rect 33458 3614 33460 3666
rect 33404 3602 33460 3614
rect 34636 3780 34692 3790
rect 34636 3666 34692 3724
rect 34636 3614 34638 3666
rect 34690 3614 34692 3666
rect 34636 3602 34692 3614
rect 35084 3556 35140 3566
rect 32508 3444 32564 3454
rect 32844 3444 32900 3482
rect 32396 3442 32564 3444
rect 32396 3390 32510 3442
rect 32562 3390 32564 3442
rect 32396 3388 32564 3390
rect 32508 3378 32564 3388
rect 32732 3388 32844 3444
rect 31276 2370 31332 2380
rect 28924 2258 28980 2268
rect 32732 2212 32788 3388
rect 32844 3378 32900 3388
rect 34188 3444 34244 3482
rect 35084 3462 35140 3500
rect 34188 3378 34244 3388
rect 37324 3442 37380 4060
rect 37324 3390 37326 3442
rect 37378 3390 37380 3442
rect 37324 3378 37380 3390
rect 37660 3554 37716 4172
rect 37884 4162 37940 4172
rect 38108 3780 38164 3790
rect 38220 3780 38276 4286
rect 38108 3778 38276 3780
rect 38108 3726 38110 3778
rect 38162 3726 38276 3778
rect 38108 3724 38276 3726
rect 38108 3714 38164 3724
rect 37660 3502 37662 3554
rect 37714 3502 37716 3554
rect 37660 3388 37716 3502
rect 38332 3554 38388 4620
rect 38332 3502 38334 3554
rect 38386 3502 38388 3554
rect 38332 3490 38388 3502
rect 33740 3332 33796 3342
rect 33740 3238 33796 3276
rect 37548 3332 37716 3388
rect 37548 2548 37604 3332
rect 32284 2156 32788 2212
rect 37212 2492 37604 2548
rect 32284 800 32340 2156
rect 37212 800 37268 2492
rect 38444 2212 38500 15092
rect 38556 14756 38612 15820
rect 38556 14690 38612 14700
rect 38668 14532 38724 15820
rect 38780 15204 38836 16940
rect 38892 16210 38948 18620
rect 38892 16158 38894 16210
rect 38946 16158 38948 16210
rect 38892 16100 38948 16158
rect 38892 16034 38948 16044
rect 38780 15148 38948 15204
rect 38668 14438 38724 14476
rect 38892 14756 38948 15148
rect 39116 14756 39172 19964
rect 39228 19908 39284 20076
rect 39228 19842 39284 19852
rect 39340 19684 39396 21196
rect 39452 20802 39508 20814
rect 39452 20750 39454 20802
rect 39506 20750 39508 20802
rect 39452 20692 39508 20750
rect 39452 20626 39508 20636
rect 40012 20690 40068 20702
rect 40012 20638 40014 20690
rect 40066 20638 40068 20690
rect 39676 20020 39732 20030
rect 39676 19926 39732 19964
rect 39340 19618 39396 19628
rect 39340 17780 39396 17790
rect 39340 14980 39396 17724
rect 39564 16884 39620 16894
rect 39564 15986 39620 16828
rect 39900 16100 39956 16110
rect 39900 16006 39956 16044
rect 39564 15934 39566 15986
rect 39618 15934 39620 15986
rect 39564 15922 39620 15934
rect 40012 15652 40068 20638
rect 40348 20690 40404 21644
rect 40460 20804 40516 22206
rect 40572 22148 40628 22158
rect 40684 22148 40740 22158
rect 40572 22146 40684 22148
rect 40572 22094 40574 22146
rect 40626 22094 40684 22146
rect 40572 22092 40684 22094
rect 40572 22082 40628 22092
rect 40572 20804 40628 20814
rect 40460 20802 40628 20804
rect 40460 20750 40574 20802
rect 40626 20750 40628 20802
rect 40460 20748 40628 20750
rect 40572 20738 40628 20748
rect 40348 20638 40350 20690
rect 40402 20638 40404 20690
rect 40124 19906 40180 19918
rect 40124 19854 40126 19906
rect 40178 19854 40180 19906
rect 40124 19572 40180 19854
rect 40348 19796 40404 20638
rect 40348 19730 40404 19740
rect 40460 20580 40516 20590
rect 40124 19506 40180 19516
rect 40124 19346 40180 19358
rect 40124 19294 40126 19346
rect 40178 19294 40180 19346
rect 40124 18228 40180 19294
rect 40460 19348 40516 20524
rect 40684 20244 40740 22092
rect 40796 22148 40852 22158
rect 40796 22146 41076 22148
rect 40796 22094 40798 22146
rect 40850 22094 41076 22146
rect 40796 22092 41076 22094
rect 40796 22082 40852 22092
rect 40908 21588 40964 21598
rect 40908 20690 40964 21532
rect 41020 21586 41076 22092
rect 41244 21810 41300 22988
rect 41468 23266 41524 23278
rect 41468 23214 41470 23266
rect 41522 23214 41524 23266
rect 41244 21758 41246 21810
rect 41298 21758 41300 21810
rect 41244 21746 41300 21758
rect 41356 22260 41412 22270
rect 41020 21534 41022 21586
rect 41074 21534 41076 21586
rect 41020 21522 41076 21534
rect 41356 21586 41412 22204
rect 41468 22148 41524 23214
rect 41580 23268 41636 26852
rect 41692 25620 41748 25630
rect 41916 25620 41972 31836
rect 41692 25618 41972 25620
rect 41692 25566 41694 25618
rect 41746 25566 41972 25618
rect 41692 25564 41972 25566
rect 42028 27074 42084 27086
rect 42028 27022 42030 27074
rect 42082 27022 42084 27074
rect 42028 26852 42084 27022
rect 41692 25554 41748 25564
rect 42028 25508 42084 26796
rect 41916 25452 42084 25508
rect 41916 25060 41972 25452
rect 42140 25284 42196 35420
rect 42252 34916 42308 35534
rect 42252 34850 42308 34860
rect 42588 34914 42644 36206
rect 42700 35812 42756 35822
rect 42700 35718 42756 35756
rect 43260 35308 43316 39200
rect 43932 36596 43988 36606
rect 43932 36502 43988 36540
rect 44132 36092 44396 36102
rect 44188 36036 44236 36092
rect 44292 36036 44340 36092
rect 44132 36026 44396 36036
rect 44716 35868 44996 35924
rect 44716 35810 44772 35868
rect 44716 35758 44718 35810
rect 44770 35758 44772 35810
rect 44716 35746 44772 35758
rect 43932 35700 43988 35710
rect 43932 35698 44100 35700
rect 43932 35646 43934 35698
rect 43986 35646 44100 35698
rect 43932 35644 44100 35646
rect 43932 35634 43988 35644
rect 42588 34862 42590 34914
rect 42642 34862 42644 34914
rect 42588 34850 42644 34862
rect 42812 35252 43316 35308
rect 43820 35586 43876 35598
rect 43820 35534 43822 35586
rect 43874 35534 43876 35586
rect 42700 34356 42756 34366
rect 42588 34354 42756 34356
rect 42588 34302 42702 34354
rect 42754 34302 42756 34354
rect 42588 34300 42756 34302
rect 42476 31778 42532 31790
rect 42476 31726 42478 31778
rect 42530 31726 42532 31778
rect 42476 30882 42532 31726
rect 42588 31668 42644 34300
rect 42700 34290 42756 34300
rect 42700 33346 42756 33358
rect 42700 33294 42702 33346
rect 42754 33294 42756 33346
rect 42700 32340 42756 33294
rect 42812 32786 42868 35196
rect 42924 34916 42980 34926
rect 42924 34822 42980 34860
rect 43820 34804 43876 35534
rect 44044 35028 44100 35644
rect 44828 35698 44884 35710
rect 44828 35646 44830 35698
rect 44882 35646 44884 35698
rect 44828 35588 44884 35646
rect 44828 35522 44884 35532
rect 43708 34244 43764 34254
rect 43820 34244 43876 34748
rect 43932 35026 44100 35028
rect 43932 34974 44046 35026
rect 44098 34974 44100 35026
rect 43932 34972 44100 34974
rect 43932 34356 43988 34972
rect 44044 34962 44100 34972
rect 44940 34802 44996 35868
rect 45500 34916 45556 39200
rect 45836 37380 45892 37390
rect 45612 35588 45668 35598
rect 45612 35494 45668 35532
rect 45500 34850 45556 34860
rect 45836 35026 45892 37324
rect 46732 36484 46788 36494
rect 46060 36372 46116 36382
rect 46060 36278 46116 36316
rect 46732 35924 46788 36428
rect 47740 36484 47796 39200
rect 47740 36418 47796 36428
rect 48860 36484 48916 36494
rect 49420 36484 49476 36494
rect 47404 36372 47460 36382
rect 47292 36370 47460 36372
rect 47292 36318 47406 36370
rect 47458 36318 47460 36370
rect 47292 36316 47460 36318
rect 46732 35858 46788 35868
rect 46844 36036 46900 36046
rect 45836 34974 45838 35026
rect 45890 34974 45892 35026
rect 44940 34750 44942 34802
rect 44994 34750 44996 34802
rect 44132 34524 44396 34534
rect 44188 34468 44236 34524
rect 44292 34468 44340 34524
rect 44132 34458 44396 34468
rect 43932 34300 44212 34356
rect 43708 34242 43876 34244
rect 43708 34190 43710 34242
rect 43762 34190 43876 34242
rect 43708 34188 43876 34190
rect 43708 34178 43764 34188
rect 44156 34130 44212 34300
rect 44940 34244 44996 34750
rect 45836 34692 45892 34974
rect 46060 35700 46116 35710
rect 46060 34914 46116 35644
rect 46396 35698 46452 35710
rect 46396 35646 46398 35698
rect 46450 35646 46452 35698
rect 46060 34862 46062 34914
rect 46114 34862 46116 34914
rect 46060 34850 46116 34862
rect 46284 35588 46340 35598
rect 45836 34626 45892 34636
rect 45164 34244 45220 34254
rect 44940 34242 45220 34244
rect 44940 34190 45166 34242
rect 45218 34190 45220 34242
rect 44940 34188 45220 34190
rect 45164 34178 45220 34188
rect 44156 34078 44158 34130
rect 44210 34078 44212 34130
rect 44156 34066 44212 34078
rect 46284 34130 46340 35532
rect 46284 34078 46286 34130
rect 46338 34078 46340 34130
rect 46284 34066 46340 34078
rect 43820 33796 43876 33806
rect 43820 33458 43876 33740
rect 45388 33460 45444 33470
rect 43820 33406 43822 33458
rect 43874 33406 43876 33458
rect 43820 33394 43876 33406
rect 45276 33458 45444 33460
rect 45276 33406 45390 33458
rect 45442 33406 45444 33458
rect 45276 33404 45444 33406
rect 43932 33348 43988 33358
rect 43932 33254 43988 33292
rect 44380 33348 44436 33358
rect 44380 33346 44660 33348
rect 44380 33294 44382 33346
rect 44434 33294 44660 33346
rect 44380 33292 44660 33294
rect 44380 33282 44436 33292
rect 43372 33236 43428 33246
rect 43708 33236 43764 33246
rect 43372 33234 43708 33236
rect 43372 33182 43374 33234
rect 43426 33182 43708 33234
rect 43372 33180 43708 33182
rect 43372 33170 43428 33180
rect 43708 33142 43764 33180
rect 44132 32956 44396 32966
rect 42812 32734 42814 32786
rect 42866 32734 42868 32786
rect 42812 32722 42868 32734
rect 43372 32900 43428 32910
rect 44188 32900 44236 32956
rect 44292 32900 44340 32956
rect 44132 32890 44396 32900
rect 43372 32562 43428 32844
rect 43932 32788 43988 32798
rect 43932 32694 43988 32732
rect 43372 32510 43374 32562
rect 43426 32510 43428 32562
rect 43372 32498 43428 32510
rect 43820 32674 43876 32686
rect 43820 32622 43822 32674
rect 43874 32622 43876 32674
rect 43820 32564 43876 32622
rect 43932 32564 43988 32574
rect 43820 32508 43932 32564
rect 43932 32498 43988 32508
rect 44044 32562 44100 32574
rect 44044 32510 44046 32562
rect 44098 32510 44100 32562
rect 43260 32452 43316 32462
rect 42700 32274 42756 32284
rect 43148 32450 43316 32452
rect 43148 32398 43262 32450
rect 43314 32398 43316 32450
rect 43148 32396 43316 32398
rect 42588 31602 42644 31612
rect 42700 31778 42756 31790
rect 42700 31726 42702 31778
rect 42754 31726 42756 31778
rect 42476 30830 42478 30882
rect 42530 30830 42532 30882
rect 42476 27970 42532 30830
rect 42588 30994 42644 31006
rect 42588 30942 42590 30994
rect 42642 30942 42644 30994
rect 42588 29988 42644 30942
rect 42588 29922 42644 29932
rect 42700 30996 42756 31726
rect 42476 27918 42478 27970
rect 42530 27918 42532 27970
rect 42364 27748 42420 27758
rect 42364 27654 42420 27692
rect 42476 27636 42532 27918
rect 42700 28754 42756 30940
rect 42924 31666 42980 31678
rect 42924 31614 42926 31666
rect 42978 31614 42980 31666
rect 42924 30324 42980 31614
rect 43148 31668 43204 32396
rect 43260 32386 43316 32396
rect 44044 32452 44100 32510
rect 44492 32452 44548 32462
rect 44044 32450 44548 32452
rect 44044 32398 44494 32450
rect 44546 32398 44548 32450
rect 44044 32396 44548 32398
rect 44044 32116 44100 32396
rect 44492 32386 44548 32396
rect 44044 32050 44100 32060
rect 43708 31892 43764 31902
rect 43708 31798 43764 31836
rect 44604 31780 44660 33292
rect 45164 33346 45220 33358
rect 45164 33294 45166 33346
rect 45218 33294 45220 33346
rect 45164 32788 45220 33294
rect 44940 32732 45164 32788
rect 44828 32564 44884 32574
rect 44716 31780 44772 31790
rect 44604 31778 44772 31780
rect 44604 31726 44718 31778
rect 44770 31726 44772 31778
rect 44604 31724 44772 31726
rect 44716 31714 44772 31724
rect 43036 30660 43092 30670
rect 43148 30660 43204 31612
rect 43596 31556 43652 31566
rect 43092 30604 43204 30660
rect 43260 31554 43652 31556
rect 43260 31502 43598 31554
rect 43650 31502 43652 31554
rect 43260 31500 43652 31502
rect 43036 30594 43092 30604
rect 43036 30324 43092 30334
rect 42924 30322 43092 30324
rect 42924 30270 43038 30322
rect 43090 30270 43092 30322
rect 42924 30268 43092 30270
rect 43036 30258 43092 30268
rect 42812 30100 42868 30110
rect 42812 30006 42868 30044
rect 43260 29988 43316 31500
rect 43596 31490 43652 31500
rect 43820 31554 43876 31566
rect 44044 31556 44100 31566
rect 43820 31502 43822 31554
rect 43874 31502 43876 31554
rect 43820 30436 43876 31502
rect 43932 31554 44100 31556
rect 43932 31502 44046 31554
rect 44098 31502 44100 31554
rect 43932 31500 44100 31502
rect 43932 31220 43988 31500
rect 44044 31490 44100 31500
rect 44132 31388 44396 31398
rect 44188 31332 44236 31388
rect 44292 31332 44340 31388
rect 44132 31322 44396 31332
rect 44828 31220 44884 32508
rect 44940 31666 44996 32732
rect 45164 32722 45220 32732
rect 45052 31780 45108 31790
rect 45276 31780 45332 33404
rect 45388 33394 45444 33404
rect 46284 33348 46340 33358
rect 46284 33254 46340 33292
rect 45836 33236 45892 33246
rect 46172 33236 46228 33246
rect 45836 33234 46228 33236
rect 45836 33182 45838 33234
rect 45890 33182 46174 33234
rect 46226 33182 46228 33234
rect 45836 33180 46228 33182
rect 45836 33170 45892 33180
rect 46172 33170 46228 33180
rect 46396 32788 46452 35646
rect 46844 35698 46900 35980
rect 46844 35646 46846 35698
rect 46898 35646 46900 35698
rect 46844 35634 46900 35646
rect 47292 35252 47348 36316
rect 47404 36306 47460 36316
rect 48300 36370 48356 36382
rect 48300 36318 48302 36370
rect 48354 36318 48356 36370
rect 47740 36260 47796 36270
rect 48300 36260 48356 36318
rect 47740 36258 47908 36260
rect 47740 36206 47742 36258
rect 47794 36206 47908 36258
rect 47740 36204 47908 36206
rect 47740 36194 47796 36204
rect 47628 35810 47684 35822
rect 47628 35758 47630 35810
rect 47682 35758 47684 35810
rect 47628 35364 47684 35758
rect 47628 35298 47684 35308
rect 47292 35186 47348 35196
rect 47516 35140 47572 35150
rect 47404 35084 47516 35140
rect 46844 34804 46900 34814
rect 46844 34710 46900 34748
rect 47068 34130 47124 34142
rect 47068 34078 47070 34130
rect 47122 34078 47124 34130
rect 46732 33460 46788 33470
rect 47068 33460 47124 34078
rect 46732 33458 47124 33460
rect 46732 33406 46734 33458
rect 46786 33406 47124 33458
rect 46732 33404 47124 33406
rect 46732 33348 46788 33404
rect 46732 33282 46788 33292
rect 47292 33236 47348 33246
rect 47292 33142 47348 33180
rect 46060 32732 46452 32788
rect 45388 32452 45444 32462
rect 45388 32358 45444 32396
rect 45724 32228 45780 32238
rect 45612 32004 45668 32014
rect 45500 31892 45556 31902
rect 45108 31724 45332 31780
rect 45388 31780 45444 31790
rect 45052 31686 45108 31724
rect 44940 31614 44942 31666
rect 44994 31614 44996 31666
rect 44940 31602 44996 31614
rect 43932 31164 44100 31220
rect 44828 31164 45332 31220
rect 43932 30996 43988 31006
rect 43932 30902 43988 30940
rect 43596 30380 43876 30436
rect 42924 29932 43316 29988
rect 43484 30210 43540 30222
rect 43484 30158 43486 30210
rect 43538 30158 43540 30210
rect 43484 29988 43540 30158
rect 42924 29650 42980 29932
rect 43484 29922 43540 29932
rect 42924 29598 42926 29650
rect 42978 29598 42980 29650
rect 42924 29586 42980 29598
rect 42812 29540 42868 29550
rect 42812 29446 42868 29484
rect 43596 29202 43652 30380
rect 44044 29988 44100 31164
rect 45164 30996 45220 31006
rect 44268 30994 45220 30996
rect 44268 30942 45166 30994
rect 45218 30942 45220 30994
rect 44268 30940 45220 30942
rect 44268 30210 44324 30940
rect 45164 30930 45220 30940
rect 44492 30772 44548 30782
rect 44492 30678 44548 30716
rect 44828 30436 44884 30446
rect 44268 30158 44270 30210
rect 44322 30158 44324 30210
rect 44268 30146 44324 30158
rect 44604 30324 44660 30334
rect 43596 29150 43598 29202
rect 43650 29150 43652 29202
rect 43596 29138 43652 29150
rect 43708 29932 44100 29988
rect 43596 28980 43652 28990
rect 42700 28702 42702 28754
rect 42754 28702 42756 28754
rect 42700 27858 42756 28702
rect 43372 28868 43428 28878
rect 43372 28754 43428 28812
rect 43372 28702 43374 28754
rect 43426 28702 43428 28754
rect 43372 28690 43428 28702
rect 42700 27806 42702 27858
rect 42754 27806 42756 27858
rect 42700 27794 42756 27806
rect 43372 27860 43428 27870
rect 43372 27766 43428 27804
rect 43372 27636 43428 27646
rect 42476 27580 42980 27636
rect 42924 27186 42980 27580
rect 42924 27134 42926 27186
rect 42978 27134 42980 27186
rect 42924 27122 42980 27134
rect 41916 24994 41972 25004
rect 42028 25228 42196 25284
rect 42252 27074 42308 27086
rect 42252 27022 42254 27074
rect 42306 27022 42308 27074
rect 42252 26964 42308 27022
rect 41916 24836 41972 24846
rect 41916 24164 41972 24780
rect 42028 24388 42084 25228
rect 42252 25172 42308 26908
rect 43260 27074 43316 27086
rect 43260 27022 43262 27074
rect 43314 27022 43316 27074
rect 43260 26964 43316 27022
rect 43260 26898 43316 26908
rect 42140 25116 42308 25172
rect 42476 25618 42532 25630
rect 42476 25566 42478 25618
rect 42530 25566 42532 25618
rect 42476 25172 42532 25566
rect 42140 24948 42196 25116
rect 42252 24948 42308 24958
rect 42140 24946 42308 24948
rect 42140 24894 42254 24946
rect 42306 24894 42308 24946
rect 42140 24892 42308 24894
rect 42252 24882 42308 24892
rect 42140 24722 42196 24734
rect 42140 24670 42142 24722
rect 42194 24670 42196 24722
rect 42140 24500 42196 24670
rect 42364 24724 42420 24734
rect 42476 24724 42532 25116
rect 42364 24722 42532 24724
rect 42364 24670 42366 24722
rect 42418 24670 42532 24722
rect 42364 24668 42532 24670
rect 42588 25506 42644 25518
rect 42588 25454 42590 25506
rect 42642 25454 42644 25506
rect 42588 24946 42644 25454
rect 43148 25508 43204 25518
rect 43372 25508 43428 27580
rect 43484 27074 43540 27086
rect 43484 27022 43486 27074
rect 43538 27022 43540 27074
rect 43484 26852 43540 27022
rect 43484 26786 43540 26796
rect 43596 25732 43652 28924
rect 43708 28866 43764 29932
rect 44132 29820 44396 29830
rect 44188 29764 44236 29820
rect 44292 29764 44340 29820
rect 44132 29754 44396 29764
rect 44156 29428 44212 29438
rect 44156 29334 44212 29372
rect 43708 28814 43710 28866
rect 43762 28814 43764 28866
rect 43708 28802 43764 28814
rect 43932 29314 43988 29326
rect 43932 29262 43934 29314
rect 43986 29262 43988 29314
rect 43932 28756 43988 29262
rect 44044 28980 44100 28990
rect 44044 28866 44100 28924
rect 44044 28814 44046 28866
rect 44098 28814 44100 28866
rect 44044 28802 44100 28814
rect 43596 25666 43652 25676
rect 43708 27858 43764 27870
rect 43708 27806 43710 27858
rect 43762 27806 43764 27858
rect 43596 25508 43652 25518
rect 43148 25506 43428 25508
rect 43148 25454 43150 25506
rect 43202 25454 43428 25506
rect 43148 25452 43428 25454
rect 43484 25452 43596 25508
rect 43148 25442 43204 25452
rect 42588 24894 42590 24946
rect 42642 24894 42644 24946
rect 42364 24658 42420 24668
rect 42588 24612 42644 24894
rect 42812 24836 42868 24846
rect 42812 24742 42868 24780
rect 42924 24724 42980 24734
rect 42924 24630 42980 24668
rect 42476 24556 42644 24612
rect 42476 24500 42532 24556
rect 42140 24444 42532 24500
rect 42028 24332 42196 24388
rect 42028 24164 42084 24174
rect 41916 24162 42084 24164
rect 41916 24110 42030 24162
rect 42082 24110 42084 24162
rect 41916 24108 42084 24110
rect 42028 24098 42084 24108
rect 41692 23938 41748 23950
rect 41692 23886 41694 23938
rect 41746 23886 41748 23938
rect 41692 23604 41748 23886
rect 41692 23538 41748 23548
rect 41580 23212 41860 23268
rect 41468 22082 41524 22092
rect 41580 23042 41636 23054
rect 41580 22990 41582 23042
rect 41634 22990 41636 23042
rect 41356 21534 41358 21586
rect 41410 21534 41412 21586
rect 41356 21522 41412 21534
rect 41580 21586 41636 22990
rect 41692 22932 41748 22942
rect 41692 22838 41748 22876
rect 41692 22370 41748 22382
rect 41692 22318 41694 22370
rect 41746 22318 41748 22370
rect 41692 22148 41748 22318
rect 41692 22082 41748 22092
rect 41580 21534 41582 21586
rect 41634 21534 41636 21586
rect 41580 21522 41636 21534
rect 41468 21028 41524 21038
rect 41244 20916 41300 20926
rect 41244 20804 41300 20860
rect 41468 20914 41524 20972
rect 41468 20862 41470 20914
rect 41522 20862 41524 20914
rect 41468 20850 41524 20862
rect 41244 20802 41412 20804
rect 41244 20750 41246 20802
rect 41298 20750 41412 20802
rect 41244 20748 41412 20750
rect 41244 20738 41300 20748
rect 40908 20638 40910 20690
rect 40962 20638 40964 20690
rect 40796 20580 40852 20590
rect 40796 20486 40852 20524
rect 40796 20244 40852 20254
rect 40684 20242 40852 20244
rect 40684 20190 40798 20242
rect 40850 20190 40852 20242
rect 40684 20188 40852 20190
rect 40796 20178 40852 20188
rect 40460 18450 40516 19292
rect 40684 19796 40740 19806
rect 40684 19346 40740 19740
rect 40684 19294 40686 19346
rect 40738 19294 40740 19346
rect 40684 19282 40740 19294
rect 40460 18398 40462 18450
rect 40514 18398 40516 18450
rect 40460 18386 40516 18398
rect 40796 18228 40852 18238
rect 40124 18162 40180 18172
rect 40684 18226 40852 18228
rect 40684 18174 40798 18226
rect 40850 18174 40852 18226
rect 40684 18172 40852 18174
rect 40348 17780 40404 17790
rect 40348 17686 40404 17724
rect 40236 16996 40292 17006
rect 40236 16770 40292 16940
rect 40236 16718 40238 16770
rect 40290 16718 40292 16770
rect 40236 16706 40292 16718
rect 40460 16100 40516 16110
rect 40460 16006 40516 16044
rect 39900 15596 40068 15652
rect 39564 15540 39620 15550
rect 39564 15202 39620 15484
rect 39564 15150 39566 15202
rect 39618 15150 39620 15202
rect 39564 15138 39620 15150
rect 39900 15148 39956 15596
rect 39340 14914 39396 14924
rect 39676 15092 39956 15148
rect 40012 15428 40068 15438
rect 39116 14700 39508 14756
rect 38892 14418 38948 14700
rect 39340 14532 39396 14542
rect 38892 14366 38894 14418
rect 38946 14366 38948 14418
rect 38892 14354 38948 14366
rect 39228 14420 39284 14430
rect 39228 14326 39284 14364
rect 39340 14418 39396 14476
rect 39340 14366 39342 14418
rect 39394 14366 39396 14418
rect 39340 14354 39396 14366
rect 38780 14308 38836 14318
rect 38668 14252 38780 14308
rect 38556 12964 38612 12974
rect 38556 12870 38612 12908
rect 38556 11394 38612 11406
rect 38556 11342 38558 11394
rect 38610 11342 38612 11394
rect 38556 10724 38612 11342
rect 38556 10658 38612 10668
rect 38668 10164 38724 14252
rect 38780 14242 38836 14252
rect 39340 13524 39396 13534
rect 39340 13074 39396 13468
rect 39340 13022 39342 13074
rect 39394 13022 39396 13074
rect 39340 13010 39396 13022
rect 39340 12290 39396 12302
rect 39340 12238 39342 12290
rect 39394 12238 39396 12290
rect 39228 12178 39284 12190
rect 39228 12126 39230 12178
rect 39282 12126 39284 12178
rect 39228 11844 39284 12126
rect 39340 12068 39396 12238
rect 39340 12002 39396 12012
rect 39228 11506 39284 11788
rect 39228 11454 39230 11506
rect 39282 11454 39284 11506
rect 39228 11442 39284 11454
rect 38780 11396 38836 11406
rect 38780 10612 38836 11340
rect 39340 10724 39396 10734
rect 39228 10668 39340 10724
rect 38892 10612 38948 10622
rect 38780 10556 38892 10612
rect 38892 10518 38948 10556
rect 39228 10610 39284 10668
rect 39340 10658 39396 10668
rect 39228 10558 39230 10610
rect 39282 10558 39284 10610
rect 38668 10052 38724 10108
rect 38556 9996 38724 10052
rect 38556 8148 38612 9996
rect 39228 9940 39284 10558
rect 39340 10500 39396 10510
rect 39452 10500 39508 14700
rect 39676 14532 39732 15092
rect 39676 14466 39732 14476
rect 40012 14530 40068 15372
rect 40684 15316 40740 18172
rect 40796 18162 40852 18172
rect 40908 16884 40964 20638
rect 41020 20130 41076 20142
rect 41020 20078 41022 20130
rect 41074 20078 41076 20130
rect 41020 19684 41076 20078
rect 41020 19618 41076 19628
rect 41132 20018 41188 20030
rect 41132 19966 41134 20018
rect 41186 19966 41188 20018
rect 41132 19460 41188 19966
rect 41356 20020 41412 20748
rect 41580 20690 41636 20702
rect 41804 20692 41860 23212
rect 41916 21028 41972 21038
rect 41916 20802 41972 20972
rect 41916 20750 41918 20802
rect 41970 20750 41972 20802
rect 41916 20738 41972 20750
rect 41580 20638 41582 20690
rect 41634 20638 41636 20690
rect 41580 20580 41636 20638
rect 41580 20514 41636 20524
rect 41692 20636 41860 20692
rect 42028 20692 42084 20702
rect 41356 19964 41524 20020
rect 41020 19404 41188 19460
rect 41020 18338 41076 19404
rect 41020 18286 41022 18338
rect 41074 18286 41076 18338
rect 41020 18226 41076 18286
rect 41020 18174 41022 18226
rect 41074 18174 41076 18226
rect 41020 18162 41076 18174
rect 41132 19234 41188 19246
rect 41132 19182 41134 19234
rect 41186 19182 41188 19234
rect 41132 17892 41188 19182
rect 41356 19012 41412 19022
rect 41356 18918 41412 18956
rect 41468 18674 41524 19964
rect 41468 18622 41470 18674
rect 41522 18622 41524 18674
rect 41468 18610 41524 18622
rect 40908 16818 40964 16828
rect 41020 17836 41132 17892
rect 40684 15250 40740 15260
rect 40796 16772 40852 16782
rect 40012 14478 40014 14530
rect 40066 14478 40068 14530
rect 40012 14466 40068 14478
rect 40236 14756 40292 14766
rect 39788 14418 39844 14430
rect 39788 14366 39790 14418
rect 39842 14366 39844 14418
rect 39564 14308 39620 14318
rect 39564 14306 39732 14308
rect 39564 14254 39566 14306
rect 39618 14254 39732 14306
rect 39564 14252 39732 14254
rect 39564 14242 39620 14252
rect 39676 13412 39732 14252
rect 39788 13860 39844 14366
rect 40236 14418 40292 14700
rect 40348 14532 40404 14542
rect 40348 14438 40404 14476
rect 40236 14366 40238 14418
rect 40290 14366 40292 14418
rect 40236 14354 40292 14366
rect 40796 14418 40852 16716
rect 40908 16548 40964 16558
rect 41020 16548 41076 17836
rect 41132 17826 41188 17836
rect 41468 17892 41524 17902
rect 41468 17778 41524 17836
rect 41468 17726 41470 17778
rect 41522 17726 41524 17778
rect 41468 17714 41524 17726
rect 41244 16996 41300 17006
rect 41244 16902 41300 16940
rect 41132 16884 41188 16894
rect 41132 16790 41188 16828
rect 41468 16882 41524 16894
rect 41468 16830 41470 16882
rect 41522 16830 41524 16882
rect 41468 16772 41524 16830
rect 41468 16706 41524 16716
rect 41020 16492 41636 16548
rect 40908 16212 40964 16492
rect 40908 15988 40964 16156
rect 41020 15988 41076 15998
rect 40908 15986 41076 15988
rect 40908 15934 41022 15986
rect 41074 15934 41076 15986
rect 40908 15932 41076 15934
rect 41020 15922 41076 15932
rect 41356 15874 41412 15886
rect 41356 15822 41358 15874
rect 41410 15822 41412 15874
rect 40908 15652 40964 15662
rect 40908 15426 40964 15596
rect 41020 15540 41076 15550
rect 41020 15446 41076 15484
rect 40908 15374 40910 15426
rect 40962 15374 40964 15426
rect 40908 15362 40964 15374
rect 41356 15428 41412 15822
rect 41468 15428 41524 15438
rect 41356 15426 41524 15428
rect 41356 15374 41470 15426
rect 41522 15374 41524 15426
rect 41356 15372 41524 15374
rect 41244 15316 41300 15326
rect 41244 15222 41300 15260
rect 40796 14366 40798 14418
rect 40850 14366 40852 14418
rect 40796 14354 40852 14366
rect 40908 14530 40964 14542
rect 40908 14478 40910 14530
rect 40962 14478 40964 14530
rect 40908 14084 40964 14478
rect 41132 14532 41188 14542
rect 41188 14476 41300 14532
rect 41132 14438 41188 14476
rect 40348 14028 40964 14084
rect 40348 13970 40404 14028
rect 40348 13918 40350 13970
rect 40402 13918 40404 13970
rect 40348 13906 40404 13918
rect 39788 13804 40180 13860
rect 39788 13636 39844 13646
rect 39788 13542 39844 13580
rect 40012 13524 40068 13534
rect 40012 13430 40068 13468
rect 40124 13412 40180 13804
rect 41244 13858 41300 14476
rect 41244 13806 41246 13858
rect 41298 13806 41300 13858
rect 41244 13794 41300 13806
rect 41132 13636 41188 13646
rect 41356 13636 41412 15372
rect 41468 15362 41524 15372
rect 39676 13356 39956 13412
rect 40124 13356 40404 13412
rect 39900 13074 39956 13356
rect 40236 13188 40292 13198
rect 39900 13022 39902 13074
rect 39954 13022 39956 13074
rect 39900 13010 39956 13022
rect 40124 13186 40292 13188
rect 40124 13134 40238 13186
rect 40290 13134 40292 13186
rect 40124 13132 40292 13134
rect 40012 12852 40068 12862
rect 40012 12402 40068 12796
rect 40012 12350 40014 12402
rect 40066 12350 40068 12402
rect 40012 12338 40068 12350
rect 39564 12292 39620 12302
rect 40124 12292 40180 13132
rect 40236 13122 40292 13132
rect 39564 12290 39732 12292
rect 39564 12238 39566 12290
rect 39618 12238 39732 12290
rect 39564 12236 39732 12238
rect 39564 12226 39620 12236
rect 39676 12178 39732 12236
rect 40124 12198 40180 12236
rect 40236 12964 40292 12974
rect 40348 12964 40404 13356
rect 40236 12962 40404 12964
rect 40236 12910 40238 12962
rect 40290 12910 40404 12962
rect 40236 12908 40404 12910
rect 41132 13074 41188 13580
rect 41132 13022 41134 13074
rect 41186 13022 41188 13074
rect 39676 12126 39678 12178
rect 39730 12126 39732 12178
rect 39676 12114 39732 12126
rect 40236 11732 40292 12908
rect 41132 12852 41188 13022
rect 41132 12786 41188 12796
rect 41244 13580 41412 13636
rect 41132 12292 41188 12302
rect 40348 12180 40404 12190
rect 40348 12178 40964 12180
rect 40348 12126 40350 12178
rect 40402 12126 40964 12178
rect 40348 12124 40964 12126
rect 40348 12114 40404 12124
rect 39788 11676 40292 11732
rect 39564 11508 39620 11518
rect 39564 11414 39620 11452
rect 39564 10836 39620 10846
rect 39564 10722 39620 10780
rect 39564 10670 39566 10722
rect 39618 10670 39620 10722
rect 39564 10658 39620 10670
rect 39788 10500 39844 11676
rect 40908 11618 40964 12124
rect 41132 12178 41188 12236
rect 41132 12126 41134 12178
rect 41186 12126 41188 12178
rect 41132 12114 41188 12126
rect 40908 11566 40910 11618
rect 40962 11566 40964 11618
rect 40908 11554 40964 11566
rect 41020 12068 41076 12078
rect 39340 10498 39508 10500
rect 39340 10446 39342 10498
rect 39394 10446 39508 10498
rect 39340 10444 39508 10446
rect 39564 10444 39844 10500
rect 39900 11506 39956 11518
rect 39900 11454 39902 11506
rect 39954 11454 39956 11506
rect 39340 10434 39396 10444
rect 39452 10052 39508 10062
rect 39228 9938 39396 9940
rect 39228 9886 39230 9938
rect 39282 9886 39396 9938
rect 39228 9884 39396 9886
rect 39228 9874 39284 9884
rect 39004 9826 39060 9838
rect 39004 9774 39006 9826
rect 39058 9774 39060 9826
rect 39004 9380 39060 9774
rect 39004 9314 39060 9324
rect 39340 9266 39396 9884
rect 39340 9214 39342 9266
rect 39394 9214 39396 9266
rect 39340 9202 39396 9214
rect 39452 9156 39508 9996
rect 39452 9090 39508 9100
rect 38892 8930 38948 8942
rect 38892 8878 38894 8930
rect 38946 8878 38948 8930
rect 38668 8820 38724 8830
rect 38668 8258 38724 8764
rect 38668 8206 38670 8258
rect 38722 8206 38724 8258
rect 38668 8194 38724 8206
rect 38780 8484 38836 8494
rect 38556 8082 38612 8092
rect 38668 7924 38724 7934
rect 38668 7698 38724 7868
rect 38668 7646 38670 7698
rect 38722 7646 38724 7698
rect 38668 7476 38724 7646
rect 38780 7586 38836 8428
rect 38892 8372 38948 8878
rect 38892 8306 38948 8316
rect 39452 7700 39508 7710
rect 39564 7700 39620 10444
rect 39900 10052 39956 11454
rect 40236 11394 40292 11406
rect 40236 11342 40238 11394
rect 40290 11342 40292 11394
rect 40124 10610 40180 10622
rect 40124 10558 40126 10610
rect 40178 10558 40180 10610
rect 40012 10052 40068 10062
rect 39676 10050 40068 10052
rect 39676 9998 40014 10050
rect 40066 9998 40068 10050
rect 39676 9996 40068 9998
rect 39676 9938 39732 9996
rect 40012 9986 40068 9996
rect 39676 9886 39678 9938
rect 39730 9886 39732 9938
rect 39676 9874 39732 9886
rect 40124 9938 40180 10558
rect 40124 9886 40126 9938
rect 40178 9886 40180 9938
rect 40124 9874 40180 9886
rect 40236 9828 40292 11342
rect 40908 11396 40964 11406
rect 41020 11396 41076 12012
rect 41244 11956 41300 13580
rect 41356 13412 41412 13422
rect 41356 13186 41412 13356
rect 41356 13134 41358 13186
rect 41410 13134 41412 13186
rect 41356 13122 41412 13134
rect 40908 11394 41076 11396
rect 40908 11342 40910 11394
rect 40962 11342 41076 11394
rect 40908 11340 41076 11342
rect 41132 11900 41300 11956
rect 40908 10836 40964 11340
rect 40572 10780 40964 10836
rect 40348 9828 40404 9838
rect 40236 9826 40404 9828
rect 40236 9774 40350 9826
rect 40402 9774 40404 9826
rect 40236 9772 40404 9774
rect 39900 9716 39956 9726
rect 39676 9604 39732 9614
rect 39676 9266 39732 9548
rect 39676 9214 39678 9266
rect 39730 9214 39732 9266
rect 39676 9202 39732 9214
rect 39508 7644 39620 7700
rect 39900 8484 39956 9660
rect 40348 9380 40404 9772
rect 40348 9314 40404 9324
rect 40012 9156 40068 9166
rect 40012 9062 40068 9100
rect 40572 8932 40628 10780
rect 40908 10612 40964 10622
rect 40908 10518 40964 10556
rect 41132 10500 41188 11900
rect 41244 11732 41300 11742
rect 41244 11618 41300 11676
rect 41244 11566 41246 11618
rect 41298 11566 41300 11618
rect 41244 11554 41300 11566
rect 41132 10406 41188 10444
rect 41468 10500 41524 10510
rect 41468 10406 41524 10444
rect 41580 10164 41636 16492
rect 41692 15148 41748 20636
rect 42028 20598 42084 20636
rect 42028 20018 42084 20030
rect 42028 19966 42030 20018
rect 42082 19966 42084 20018
rect 41804 19906 41860 19918
rect 41804 19854 41806 19906
rect 41858 19854 41860 19906
rect 41804 19236 41860 19854
rect 41804 18450 41860 19180
rect 41804 18398 41806 18450
rect 41858 18398 41860 18450
rect 41804 18386 41860 18398
rect 42028 19346 42084 19966
rect 42028 19294 42030 19346
rect 42082 19294 42084 19346
rect 42028 19012 42084 19294
rect 42028 18452 42084 18956
rect 42028 18358 42084 18396
rect 42028 17554 42084 17566
rect 42028 17502 42030 17554
rect 42082 17502 42084 17554
rect 42028 16884 42084 17502
rect 42028 16818 42084 16828
rect 42140 15876 42196 24332
rect 42700 23938 42756 23950
rect 42700 23886 42702 23938
rect 42754 23886 42756 23938
rect 42700 23716 42756 23886
rect 42700 23650 42756 23660
rect 42924 23714 42980 23726
rect 43484 23716 43540 25452
rect 43596 25442 43652 25452
rect 43708 24164 43764 27806
rect 43820 27860 43876 27870
rect 43820 27298 43876 27804
rect 43932 27748 43988 28700
rect 44268 28644 44324 28654
rect 44268 28550 44324 28588
rect 44132 28252 44396 28262
rect 44188 28196 44236 28252
rect 44292 28196 44340 28252
rect 44132 28186 44396 28196
rect 44268 27860 44324 27870
rect 44268 27766 44324 27804
rect 43932 27682 43988 27692
rect 43820 27246 43822 27298
rect 43874 27246 43876 27298
rect 43820 27234 43876 27246
rect 44604 26908 44660 30268
rect 44716 28868 44772 28878
rect 44716 28196 44772 28812
rect 44828 28420 44884 30380
rect 45164 29988 45220 29998
rect 45052 29986 45220 29988
rect 45052 29934 45166 29986
rect 45218 29934 45220 29986
rect 45052 29932 45220 29934
rect 44940 29652 44996 29662
rect 45052 29652 45108 29932
rect 45164 29922 45220 29932
rect 45276 29764 45332 31164
rect 45388 31218 45444 31724
rect 45388 31166 45390 31218
rect 45442 31166 45444 31218
rect 45388 31154 45444 31166
rect 45500 31106 45556 31836
rect 45612 31778 45668 31948
rect 45724 31890 45780 32172
rect 45724 31838 45726 31890
rect 45778 31838 45780 31890
rect 45724 31826 45780 31838
rect 45612 31726 45614 31778
rect 45666 31726 45668 31778
rect 45612 31714 45668 31726
rect 45500 31054 45502 31106
rect 45554 31054 45556 31106
rect 45500 30772 45556 31054
rect 45948 31108 46004 31118
rect 45948 31014 46004 31052
rect 45500 30706 45556 30716
rect 45836 30322 45892 30334
rect 45836 30270 45838 30322
rect 45890 30270 45892 30322
rect 44996 29596 45108 29652
rect 45164 29708 45332 29764
rect 45724 30212 45780 30222
rect 44940 29586 44996 29596
rect 44940 29314 44996 29326
rect 44940 29262 44942 29314
rect 44994 29262 44996 29314
rect 44940 28980 44996 29262
rect 44940 28866 44996 28924
rect 44940 28814 44942 28866
rect 44994 28814 44996 28866
rect 44940 28802 44996 28814
rect 45052 28530 45108 28542
rect 45052 28478 45054 28530
rect 45106 28478 45108 28530
rect 44828 28354 44884 28364
rect 44940 28418 44996 28430
rect 44940 28366 44942 28418
rect 44994 28366 44996 28418
rect 44940 28196 44996 28366
rect 44716 28140 44996 28196
rect 45052 27972 45108 28478
rect 44492 26852 44660 26908
rect 44716 27916 45108 27972
rect 44716 26908 44772 27916
rect 45052 27748 45108 27758
rect 44940 27186 44996 27198
rect 44940 27134 44942 27186
rect 44994 27134 44996 27186
rect 44940 27076 44996 27134
rect 44716 26852 44884 26908
rect 44132 26684 44396 26694
rect 44188 26628 44236 26684
rect 44292 26628 44340 26684
rect 44132 26618 44396 26628
rect 44492 26628 44548 26852
rect 44492 26572 44772 26628
rect 44492 26404 44548 26414
rect 44492 26310 44548 26348
rect 44604 26292 44660 26302
rect 44604 26198 44660 26236
rect 44492 26066 44548 26078
rect 44492 26014 44494 26066
rect 44546 26014 44548 26066
rect 43932 25732 43988 25742
rect 43932 25506 43988 25676
rect 43932 25454 43934 25506
rect 43986 25454 43988 25506
rect 43932 25442 43988 25454
rect 44492 25508 44548 26014
rect 44716 25508 44772 26572
rect 44492 25506 44772 25508
rect 44492 25454 44718 25506
rect 44770 25454 44772 25506
rect 44492 25452 44772 25454
rect 44716 25442 44772 25452
rect 44268 25396 44324 25406
rect 44268 25394 44660 25396
rect 44268 25342 44270 25394
rect 44322 25342 44660 25394
rect 44268 25340 44660 25342
rect 44268 25330 44324 25340
rect 44156 25284 44212 25294
rect 43932 25282 44212 25284
rect 43932 25230 44158 25282
rect 44210 25230 44212 25282
rect 43932 25228 44212 25230
rect 43932 24948 43988 25228
rect 44156 25218 44212 25228
rect 44132 25116 44396 25126
rect 44188 25060 44236 25116
rect 44292 25060 44340 25116
rect 44132 25050 44396 25060
rect 43932 24882 43988 24892
rect 44044 24834 44100 24846
rect 44044 24782 44046 24834
rect 44098 24782 44100 24834
rect 43932 24722 43988 24734
rect 43932 24670 43934 24722
rect 43986 24670 43988 24722
rect 43932 24388 43988 24670
rect 44044 24724 44100 24782
rect 44044 24658 44100 24668
rect 44268 24724 44324 24734
rect 44604 24724 44660 25340
rect 44268 24722 44660 24724
rect 44268 24670 44270 24722
rect 44322 24670 44606 24722
rect 44658 24670 44660 24722
rect 44268 24668 44660 24670
rect 44268 24658 44324 24668
rect 44604 24658 44660 24668
rect 43932 24322 43988 24332
rect 43596 24108 43764 24164
rect 43596 24052 43652 24108
rect 43596 23986 43652 23996
rect 43932 24052 43988 24062
rect 44828 24052 44884 26852
rect 43708 23940 43764 23950
rect 42924 23662 42926 23714
rect 42978 23662 42980 23714
rect 42812 23380 42868 23390
rect 42812 23286 42868 23324
rect 42924 23156 42980 23662
rect 43372 23660 43540 23716
rect 43596 23714 43652 23726
rect 43596 23662 43598 23714
rect 43650 23662 43652 23714
rect 43260 23380 43316 23390
rect 42980 23100 43204 23156
rect 42924 23090 42980 23100
rect 42588 22932 42644 22942
rect 42588 22370 42644 22876
rect 42588 22318 42590 22370
rect 42642 22318 42644 22370
rect 42588 22306 42644 22318
rect 42364 21586 42420 21598
rect 42364 21534 42366 21586
rect 42418 21534 42420 21586
rect 42364 20130 42420 21534
rect 42364 20078 42366 20130
rect 42418 20078 42420 20130
rect 42364 20020 42420 20078
rect 42364 19954 42420 19964
rect 42924 21588 42980 21598
rect 42924 20580 42980 21532
rect 43148 21364 43204 23100
rect 43260 23154 43316 23324
rect 43260 23102 43262 23154
rect 43314 23102 43316 23154
rect 43260 23090 43316 23102
rect 43260 22484 43316 22494
rect 43372 22484 43428 23660
rect 43484 23492 43540 23502
rect 43596 23492 43652 23662
rect 43540 23436 43652 23492
rect 43484 23378 43540 23436
rect 43484 23326 43486 23378
rect 43538 23326 43540 23378
rect 43484 23314 43540 23326
rect 43260 22482 43428 22484
rect 43260 22430 43262 22482
rect 43314 22430 43428 22482
rect 43260 22428 43428 22430
rect 43260 22418 43316 22428
rect 43708 21700 43764 23884
rect 43820 23492 43876 23502
rect 43820 23154 43876 23436
rect 43820 23102 43822 23154
rect 43874 23102 43876 23154
rect 43820 23090 43876 23102
rect 43820 21700 43876 21710
rect 43708 21698 43876 21700
rect 43708 21646 43822 21698
rect 43874 21646 43876 21698
rect 43708 21644 43876 21646
rect 43820 21634 43876 21644
rect 43148 21298 43204 21308
rect 42252 19234 42308 19246
rect 42252 19182 42254 19234
rect 42306 19182 42308 19234
rect 42252 18452 42308 19182
rect 42700 18676 42756 18686
rect 42700 18582 42756 18620
rect 42364 18452 42420 18462
rect 42252 18450 42420 18452
rect 42252 18398 42366 18450
rect 42418 18398 42420 18450
rect 42252 18396 42420 18398
rect 42364 17106 42420 18396
rect 42924 18340 42980 20524
rect 43932 20802 43988 23996
rect 44492 23996 44884 24052
rect 44132 23548 44396 23558
rect 44188 23492 44236 23548
rect 44292 23492 44340 23548
rect 44132 23482 44396 23492
rect 44044 22930 44100 22942
rect 44044 22878 44046 22930
rect 44098 22878 44100 22930
rect 44044 22484 44100 22878
rect 44380 22932 44436 22942
rect 44380 22838 44436 22876
rect 44044 22418 44100 22428
rect 44492 22484 44548 23996
rect 44940 23940 44996 27020
rect 45052 25396 45108 27692
rect 45164 25618 45220 29708
rect 45500 29652 45556 29662
rect 45276 29426 45332 29438
rect 45276 29374 45278 29426
rect 45330 29374 45332 29426
rect 45276 28644 45332 29374
rect 45276 28550 45332 28588
rect 45500 28532 45556 29596
rect 45724 29540 45780 30156
rect 45724 29446 45780 29484
rect 45724 28756 45780 28766
rect 45836 28756 45892 30270
rect 46060 29316 46116 32732
rect 46284 32562 46340 32574
rect 46284 32510 46286 32562
rect 46338 32510 46340 32562
rect 46172 31778 46228 31790
rect 46172 31726 46174 31778
rect 46226 31726 46228 31778
rect 46172 30996 46228 31726
rect 46284 31780 46340 32510
rect 46620 32562 46676 32574
rect 46620 32510 46622 32562
rect 46674 32510 46676 32562
rect 46620 31892 46676 32510
rect 46620 31826 46676 31836
rect 46732 32450 46788 32462
rect 46732 32398 46734 32450
rect 46786 32398 46788 32450
rect 46284 31714 46340 31724
rect 46396 30996 46452 31006
rect 46172 30994 46452 30996
rect 46172 30942 46398 30994
rect 46450 30942 46452 30994
rect 46172 30940 46452 30942
rect 46284 30098 46340 30110
rect 46284 30046 46286 30098
rect 46338 30046 46340 30098
rect 46284 29428 46340 30046
rect 46396 29652 46452 30940
rect 46732 30994 46788 32398
rect 47180 32450 47236 32462
rect 47180 32398 47182 32450
rect 47234 32398 47236 32450
rect 47180 32116 47236 32398
rect 47180 32050 47236 32060
rect 46956 32004 47012 32014
rect 46956 31910 47012 31948
rect 46844 31668 46900 31678
rect 47068 31668 47124 31678
rect 46900 31666 47124 31668
rect 46900 31614 47070 31666
rect 47122 31614 47124 31666
rect 46900 31612 47124 31614
rect 46844 31602 46900 31612
rect 47068 31602 47124 31612
rect 47404 31220 47460 35084
rect 47516 35074 47572 35084
rect 47628 34914 47684 34926
rect 47628 34862 47630 34914
rect 47682 34862 47684 34914
rect 47516 34130 47572 34142
rect 47516 34078 47518 34130
rect 47570 34078 47572 34130
rect 47516 33348 47572 34078
rect 47516 33282 47572 33292
rect 47628 33572 47684 34862
rect 47852 34914 47908 36204
rect 48300 36194 48356 36204
rect 48748 35812 48804 35822
rect 48748 35718 48804 35756
rect 47852 34862 47854 34914
rect 47906 34862 47908 34914
rect 47852 34850 47908 34862
rect 47964 35698 48020 35710
rect 47964 35646 47966 35698
rect 48018 35646 48020 35698
rect 47964 34916 48020 35646
rect 48860 35588 48916 36428
rect 49308 36482 49476 36484
rect 49308 36430 49422 36482
rect 49474 36430 49476 36482
rect 49308 36428 49476 36430
rect 49196 36372 49252 36382
rect 49196 36278 49252 36316
rect 49308 36148 49364 36428
rect 49420 36418 49476 36428
rect 49980 36372 50036 39200
rect 52108 37044 52164 37054
rect 51286 36876 51550 36886
rect 51342 36820 51390 36876
rect 51446 36820 51494 36876
rect 51286 36810 51550 36820
rect 49980 36306 50036 36316
rect 50540 36372 50596 36382
rect 50540 36278 50596 36316
rect 51660 36370 51716 36382
rect 51660 36318 51662 36370
rect 51714 36318 51716 36370
rect 48860 35522 48916 35532
rect 49084 35812 49140 35822
rect 47740 34132 47796 34142
rect 47740 34038 47796 34076
rect 47964 33908 48020 34860
rect 48972 35028 49028 35038
rect 48188 34692 48244 34702
rect 48188 34354 48244 34636
rect 48188 34302 48190 34354
rect 48242 34302 48244 34354
rect 48188 34290 48244 34302
rect 48860 34242 48916 34254
rect 48860 34190 48862 34242
rect 48914 34190 48916 34242
rect 48748 34132 48804 34142
rect 48748 34038 48804 34076
rect 48860 33908 48916 34190
rect 48972 34020 49028 34972
rect 49084 35026 49140 35756
rect 49196 35476 49252 35486
rect 49308 35476 49364 36092
rect 50204 36258 50260 36270
rect 50204 36206 50206 36258
rect 50258 36206 50260 36258
rect 50204 35700 50260 36206
rect 51436 35924 51492 35934
rect 51436 35830 51492 35868
rect 50204 35634 50260 35644
rect 50652 35810 50708 35822
rect 50652 35758 50654 35810
rect 50706 35758 50708 35810
rect 49252 35420 49364 35476
rect 49420 35476 49476 35486
rect 49196 35410 49252 35420
rect 49084 34974 49086 35026
rect 49138 34974 49140 35026
rect 49084 34962 49140 34974
rect 49420 34914 49476 35420
rect 50316 34916 50372 34926
rect 49420 34862 49422 34914
rect 49474 34862 49476 34914
rect 49420 34850 49476 34862
rect 50204 34914 50372 34916
rect 50204 34862 50318 34914
rect 50370 34862 50372 34914
rect 50204 34860 50372 34862
rect 49868 34804 49924 34814
rect 49868 34710 49924 34748
rect 49980 34468 50036 34478
rect 49084 34244 49140 34254
rect 49420 34244 49476 34254
rect 49084 34242 49476 34244
rect 49084 34190 49086 34242
rect 49138 34190 49422 34242
rect 49474 34190 49476 34242
rect 49084 34188 49476 34190
rect 49084 34178 49140 34188
rect 49420 34178 49476 34188
rect 49532 34132 49588 34142
rect 49532 34130 49812 34132
rect 49532 34078 49534 34130
rect 49586 34078 49812 34130
rect 49532 34076 49812 34078
rect 49532 34066 49588 34076
rect 48972 33964 49476 34020
rect 47964 33842 48020 33852
rect 48748 33852 48916 33908
rect 49420 33906 49476 33964
rect 49420 33854 49422 33906
rect 49474 33854 49476 33906
rect 47628 33124 47684 33516
rect 48188 33348 48244 33358
rect 48188 33254 48244 33292
rect 48748 33236 48804 33852
rect 49420 33842 49476 33854
rect 48860 33684 48916 33694
rect 48860 33458 48916 33628
rect 48860 33406 48862 33458
rect 48914 33406 48916 33458
rect 48860 33394 48916 33406
rect 49196 33348 49252 33358
rect 49196 33346 49476 33348
rect 49196 33294 49198 33346
rect 49250 33294 49476 33346
rect 49196 33292 49476 33294
rect 49196 33282 49252 33292
rect 48748 33170 48804 33180
rect 47628 33058 47684 33068
rect 48524 33124 48580 33134
rect 47852 32676 47908 32686
rect 47852 32674 48020 32676
rect 47852 32622 47854 32674
rect 47906 32622 48020 32674
rect 47852 32620 48020 32622
rect 47852 32610 47908 32620
rect 46732 30942 46734 30994
rect 46786 30942 46788 30994
rect 46732 30930 46788 30942
rect 47068 31164 47460 31220
rect 46396 29586 46452 29596
rect 46172 29316 46228 29326
rect 46116 29314 46228 29316
rect 46116 29262 46174 29314
rect 46226 29262 46228 29314
rect 46116 29260 46228 29262
rect 46060 29222 46116 29260
rect 46172 29250 46228 29260
rect 45780 28700 45892 28756
rect 45724 28690 45780 28700
rect 45388 28530 45556 28532
rect 45388 28478 45502 28530
rect 45554 28478 45556 28530
rect 45388 28476 45556 28478
rect 45276 28420 45332 28430
rect 45276 27524 45332 28364
rect 45276 27458 45332 27468
rect 45388 27300 45444 28476
rect 45500 28466 45556 28476
rect 45612 28530 45668 28542
rect 45612 28478 45614 28530
rect 45666 28478 45668 28530
rect 45500 28308 45556 28318
rect 45500 27860 45556 28252
rect 45500 27766 45556 27804
rect 45612 27300 45668 28478
rect 46284 28532 46340 29372
rect 46396 28756 46452 28766
rect 46396 28662 46452 28700
rect 46620 28532 46676 28542
rect 46284 28530 46676 28532
rect 46284 28478 46622 28530
rect 46674 28478 46676 28530
rect 46284 28476 46676 28478
rect 46284 28308 46340 28476
rect 46620 28466 46676 28476
rect 46284 28242 46340 28252
rect 45948 27860 46004 27870
rect 45948 27766 46004 27804
rect 46844 27858 46900 27870
rect 46844 27806 46846 27858
rect 46898 27806 46900 27858
rect 45276 27244 45444 27300
rect 45500 27244 45668 27300
rect 46620 27524 46676 27534
rect 46620 27298 46676 27468
rect 46620 27246 46622 27298
rect 46674 27246 46676 27298
rect 45276 26908 45332 27244
rect 45388 27076 45444 27086
rect 45500 27076 45556 27244
rect 46620 27234 46676 27246
rect 46844 27188 46900 27806
rect 46956 27746 47012 27758
rect 46956 27694 46958 27746
rect 47010 27694 47012 27746
rect 46956 27300 47012 27694
rect 46956 27206 47012 27244
rect 46844 27122 46900 27132
rect 45388 27074 45500 27076
rect 45388 27022 45390 27074
rect 45442 27022 45500 27074
rect 45388 27020 45500 27022
rect 45388 27010 45444 27020
rect 45500 27010 45556 27020
rect 46060 27074 46116 27086
rect 46060 27022 46062 27074
rect 46114 27022 46116 27074
rect 46060 26908 46116 27022
rect 46284 27076 46340 27086
rect 46284 26982 46340 27020
rect 45276 26852 46116 26908
rect 45388 26516 45444 26526
rect 45500 26516 45556 26852
rect 45388 26514 45556 26516
rect 45388 26462 45390 26514
rect 45442 26462 45556 26514
rect 45388 26460 45556 26462
rect 45388 26450 45444 26460
rect 46620 26404 46676 26414
rect 46620 26310 46676 26348
rect 45164 25566 45166 25618
rect 45218 25566 45220 25618
rect 45164 25554 45220 25566
rect 45948 26292 46004 26302
rect 45388 25508 45444 25518
rect 45388 25506 45556 25508
rect 45388 25454 45390 25506
rect 45442 25454 45556 25506
rect 45388 25452 45556 25454
rect 45388 25442 45444 25452
rect 45052 25340 45220 25396
rect 45052 24724 45108 24734
rect 45052 24630 45108 24668
rect 44492 22418 44548 22428
rect 44604 23884 44996 23940
rect 45052 24500 45108 24510
rect 45052 23940 45108 24444
rect 45164 24052 45220 25340
rect 45164 23986 45220 23996
rect 45276 24948 45332 24958
rect 45276 24050 45332 24892
rect 45500 24834 45556 25452
rect 45948 25396 46004 26236
rect 45500 24782 45502 24834
rect 45554 24782 45556 24834
rect 45500 24770 45556 24782
rect 45836 24948 45892 24958
rect 45836 24834 45892 24892
rect 45836 24782 45838 24834
rect 45890 24782 45892 24834
rect 45836 24770 45892 24782
rect 45276 23998 45278 24050
rect 45330 23998 45332 24050
rect 45276 23986 45332 23998
rect 45948 24500 46004 25340
rect 46060 26290 46116 26302
rect 46060 26238 46062 26290
rect 46114 26238 46116 26290
rect 46060 24724 46116 26238
rect 46508 26290 46564 26302
rect 46508 26238 46510 26290
rect 46562 26238 46564 26290
rect 46508 25844 46564 26238
rect 46956 26180 47012 26190
rect 46956 26086 47012 26124
rect 47068 26068 47124 31164
rect 47964 30994 48020 32620
rect 48076 32562 48132 32574
rect 48076 32510 48078 32562
rect 48130 32510 48132 32562
rect 48076 31666 48132 32510
rect 48188 31780 48244 31790
rect 48188 31686 48244 31724
rect 48076 31614 48078 31666
rect 48130 31614 48132 31666
rect 48076 31556 48132 31614
rect 48076 31500 48244 31556
rect 47964 30942 47966 30994
rect 48018 30942 48020 30994
rect 47964 30930 48020 30942
rect 48076 30884 48132 30894
rect 47180 30212 47236 30222
rect 47180 30118 47236 30156
rect 47964 29876 48020 29886
rect 47964 29650 48020 29820
rect 47964 29598 47966 29650
rect 48018 29598 48020 29650
rect 47964 29586 48020 29598
rect 48076 29650 48132 30828
rect 48188 30772 48244 31500
rect 48188 30706 48244 30716
rect 48524 30098 48580 33068
rect 49308 33122 49364 33134
rect 49308 33070 49310 33122
rect 49362 33070 49364 33122
rect 48748 32676 48804 32686
rect 48748 32582 48804 32620
rect 49308 32004 49364 33070
rect 49308 31938 49364 31948
rect 49420 32562 49476 33292
rect 49420 32510 49422 32562
rect 49474 32510 49476 32562
rect 49084 31892 49140 31902
rect 48860 31780 48916 31790
rect 48860 30882 48916 31724
rect 49084 31778 49140 31836
rect 49084 31726 49086 31778
rect 49138 31726 49140 31778
rect 49084 31714 49140 31726
rect 49420 31668 49476 32510
rect 49532 33346 49588 33358
rect 49532 33294 49534 33346
rect 49586 33294 49588 33346
rect 49532 32004 49588 33294
rect 49756 33346 49812 34076
rect 49756 33294 49758 33346
rect 49810 33294 49812 33346
rect 49756 33282 49812 33294
rect 49980 33234 50036 34412
rect 50092 34130 50148 34142
rect 50092 34078 50094 34130
rect 50146 34078 50148 34130
rect 50092 33572 50148 34078
rect 50092 33506 50148 33516
rect 50204 33684 50260 34860
rect 50316 34850 50372 34860
rect 50540 34914 50596 34926
rect 50540 34862 50542 34914
rect 50594 34862 50596 34914
rect 50540 34468 50596 34862
rect 50652 34692 50708 35758
rect 51660 35812 51716 36318
rect 51772 35812 51828 35822
rect 51660 35756 51772 35812
rect 51772 35718 51828 35756
rect 50876 35588 50932 35598
rect 50876 35494 50932 35532
rect 52108 35586 52164 36988
rect 52220 36484 52276 39200
rect 52220 36418 52276 36428
rect 52780 36482 52836 36494
rect 53116 36484 53172 36494
rect 52780 36430 52782 36482
rect 52834 36430 52836 36482
rect 52780 35924 52836 36430
rect 52108 35534 52110 35586
rect 52162 35534 52164 35586
rect 52108 35522 52164 35534
rect 52668 35868 52780 35924
rect 51286 35308 51550 35318
rect 51342 35252 51390 35308
rect 51446 35252 51494 35308
rect 51286 35242 51550 35252
rect 51212 35028 51268 35038
rect 51212 34934 51268 34972
rect 52668 35026 52724 35868
rect 52780 35858 52836 35868
rect 52892 36482 53172 36484
rect 52892 36430 53118 36482
rect 53170 36430 53172 36482
rect 52892 36428 53172 36430
rect 52780 35698 52836 35710
rect 52780 35646 52782 35698
rect 52834 35646 52836 35698
rect 52780 35588 52836 35646
rect 52780 35522 52836 35532
rect 52668 34974 52670 35026
rect 52722 34974 52724 35026
rect 52668 34962 52724 34974
rect 52892 35138 52948 36428
rect 53116 36418 53172 36428
rect 53788 36484 53844 36494
rect 53788 36390 53844 36428
rect 54460 36484 54516 39200
rect 56252 37268 56308 37278
rect 55020 36708 55076 36718
rect 55020 36594 55076 36652
rect 55020 36542 55022 36594
rect 55074 36542 55076 36594
rect 55020 36530 55076 36542
rect 54460 36418 54516 36428
rect 55468 36484 55524 36494
rect 55524 36428 55972 36484
rect 55468 36390 55524 36428
rect 53564 36258 53620 36270
rect 53564 36206 53566 36258
rect 53618 36206 53620 36258
rect 53564 36036 53620 36206
rect 54460 36260 54516 36270
rect 54460 36258 55188 36260
rect 54460 36206 54462 36258
rect 54514 36206 55188 36258
rect 54460 36204 55188 36206
rect 54460 36194 54516 36204
rect 54572 36092 54852 36148
rect 54572 36036 54628 36092
rect 53564 35970 53620 35980
rect 54460 35980 54628 36036
rect 53564 35700 53620 35710
rect 53452 35698 53620 35700
rect 53452 35646 53566 35698
rect 53618 35646 53620 35698
rect 53452 35644 53620 35646
rect 52892 35086 52894 35138
rect 52946 35086 52948 35138
rect 52892 35028 52948 35086
rect 53228 35140 53284 35150
rect 53452 35140 53508 35644
rect 53564 35634 53620 35644
rect 53228 35138 53508 35140
rect 53228 35086 53230 35138
rect 53282 35086 53508 35138
rect 53228 35084 53508 35086
rect 53228 35074 53284 35084
rect 52892 34962 52948 34972
rect 51548 34804 51604 34814
rect 54236 34804 54292 34814
rect 54460 34804 54516 35980
rect 54684 35924 54740 35934
rect 54684 35830 54740 35868
rect 54796 35922 54852 36092
rect 54796 35870 54798 35922
rect 54850 35870 54852 35922
rect 54796 35858 54852 35870
rect 54572 35698 54628 35710
rect 54572 35646 54574 35698
rect 54626 35646 54628 35698
rect 54572 35140 54628 35646
rect 54572 35084 54740 35140
rect 51548 34710 51604 34748
rect 53900 34802 54516 34804
rect 53900 34750 54238 34802
rect 54290 34750 54516 34802
rect 53900 34748 54516 34750
rect 54572 34914 54628 34926
rect 54572 34862 54574 34914
rect 54626 34862 54628 34914
rect 50652 34626 50708 34636
rect 50988 34692 51044 34702
rect 50540 34354 50596 34412
rect 50540 34302 50542 34354
rect 50594 34302 50596 34354
rect 50540 34290 50596 34302
rect 50428 34242 50484 34254
rect 50428 34190 50430 34242
rect 50482 34190 50484 34242
rect 50428 34132 50484 34190
rect 50540 34132 50596 34142
rect 50428 34076 50540 34132
rect 50540 34066 50596 34076
rect 50652 34132 50708 34142
rect 50652 34130 50820 34132
rect 50652 34078 50654 34130
rect 50706 34078 50820 34130
rect 50652 34076 50820 34078
rect 50652 34066 50708 34076
rect 50092 33348 50148 33358
rect 50204 33348 50260 33628
rect 50092 33346 50260 33348
rect 50092 33294 50094 33346
rect 50146 33294 50260 33346
rect 50092 33292 50260 33294
rect 50540 33796 50596 33806
rect 50092 33282 50148 33292
rect 49980 33182 49982 33234
rect 50034 33182 50036 33234
rect 49980 33170 50036 33182
rect 50428 33236 50484 33246
rect 50428 33142 50484 33180
rect 50540 32676 50596 33740
rect 50764 33570 50820 34076
rect 50988 33796 51044 34636
rect 51660 34692 51716 34702
rect 51660 34598 51716 34636
rect 51884 34690 51940 34702
rect 51884 34638 51886 34690
rect 51938 34638 51940 34690
rect 51884 34356 51940 34638
rect 51884 34290 51940 34300
rect 51548 34132 51604 34142
rect 51604 34076 51716 34132
rect 51548 34038 51604 34076
rect 50988 33730 51044 33740
rect 51100 34018 51156 34030
rect 51100 33966 51102 34018
rect 51154 33966 51156 34018
rect 50764 33518 50766 33570
rect 50818 33518 50820 33570
rect 50764 33506 50820 33518
rect 50764 33348 50820 33358
rect 51100 33348 51156 33966
rect 51286 33740 51550 33750
rect 51342 33684 51390 33740
rect 51446 33684 51494 33740
rect 51286 33674 51550 33684
rect 51212 33572 51268 33582
rect 51212 33478 51268 33516
rect 51548 33572 51604 33582
rect 50764 33346 51156 33348
rect 50764 33294 50766 33346
rect 50818 33294 51156 33346
rect 50764 33292 51156 33294
rect 50764 33282 50820 33292
rect 51100 33236 51156 33292
rect 51212 33236 51268 33246
rect 51100 33234 51268 33236
rect 51100 33182 51214 33234
rect 51266 33182 51268 33234
rect 51100 33180 51268 33182
rect 50540 32674 50708 32676
rect 50540 32622 50542 32674
rect 50594 32622 50708 32674
rect 50540 32620 50708 32622
rect 50540 32610 50596 32620
rect 49532 31938 49588 31948
rect 50204 32004 50260 32014
rect 50092 31668 50148 31678
rect 49420 31666 50148 31668
rect 49420 31614 50094 31666
rect 50146 31614 50148 31666
rect 49420 31612 50148 31614
rect 48860 30830 48862 30882
rect 48914 30830 48916 30882
rect 48860 30818 48916 30830
rect 49084 30994 49140 31006
rect 49084 30942 49086 30994
rect 49138 30942 49140 30994
rect 48524 30046 48526 30098
rect 48578 30046 48580 30098
rect 48524 30034 48580 30046
rect 48972 30322 49028 30334
rect 48972 30270 48974 30322
rect 49026 30270 49028 30322
rect 48972 29876 49028 30270
rect 48076 29598 48078 29650
rect 48130 29598 48132 29650
rect 48076 29586 48132 29598
rect 48860 29820 48972 29876
rect 48188 29204 48244 29214
rect 48188 29110 48244 29148
rect 48860 28756 48916 29820
rect 48972 29810 49028 29820
rect 48972 29652 49028 29662
rect 48972 29558 49028 29596
rect 48860 28700 49028 28756
rect 48188 28642 48244 28654
rect 48188 28590 48190 28642
rect 48242 28590 48244 28642
rect 48188 28084 48244 28590
rect 47292 28028 48244 28084
rect 47292 27970 47348 28028
rect 47292 27918 47294 27970
rect 47346 27918 47348 27970
rect 47292 27906 47348 27918
rect 48188 27970 48244 28028
rect 48188 27918 48190 27970
rect 48242 27918 48244 27970
rect 48188 27906 48244 27918
rect 47628 27860 47684 27870
rect 47404 27858 47684 27860
rect 47404 27806 47630 27858
rect 47682 27806 47684 27858
rect 47404 27804 47684 27806
rect 47292 27300 47348 27310
rect 47404 27300 47460 27804
rect 47628 27794 47684 27804
rect 47852 27860 47908 27870
rect 47852 27766 47908 27804
rect 48076 27860 48132 27870
rect 48076 27766 48132 27804
rect 48860 27748 48916 27758
rect 48300 27746 48916 27748
rect 48300 27694 48862 27746
rect 48914 27694 48916 27746
rect 48300 27692 48916 27694
rect 47292 27298 47460 27300
rect 47292 27246 47294 27298
rect 47346 27246 47460 27298
rect 47292 27244 47460 27246
rect 47516 27412 47572 27422
rect 47292 27234 47348 27244
rect 47180 27188 47236 27198
rect 47180 26962 47236 27132
rect 47180 26910 47182 26962
rect 47234 26910 47236 26962
rect 47180 26898 47236 26910
rect 47292 27076 47348 27086
rect 47068 26002 47124 26012
rect 47180 26068 47236 26078
rect 47292 26068 47348 27020
rect 47516 26908 47572 27356
rect 47740 27300 47796 27310
rect 47740 27206 47796 27244
rect 47852 27076 47908 27086
rect 47852 26982 47908 27020
rect 47740 26962 47796 26974
rect 47740 26910 47742 26962
rect 47794 26910 47796 26962
rect 47740 26908 47796 26910
rect 47516 26852 47796 26908
rect 47516 26628 47572 26638
rect 47516 26514 47572 26572
rect 47516 26462 47518 26514
rect 47570 26462 47572 26514
rect 47516 26450 47572 26462
rect 47180 26066 47348 26068
rect 47180 26014 47182 26066
rect 47234 26014 47348 26066
rect 47180 26012 47348 26014
rect 47180 26002 47236 26012
rect 46284 25788 47012 25844
rect 46172 25620 46228 25630
rect 46172 25526 46228 25564
rect 46060 24658 46116 24668
rect 46060 24500 46116 24510
rect 45948 24498 46116 24500
rect 45948 24446 46062 24498
rect 46114 24446 46116 24498
rect 45948 24444 46116 24446
rect 44380 22372 44436 22382
rect 44380 22278 44436 22316
rect 44132 21980 44396 21990
rect 44188 21924 44236 21980
rect 44292 21924 44340 21980
rect 44132 21914 44396 21924
rect 44380 21698 44436 21710
rect 44380 21646 44382 21698
rect 44434 21646 44436 21698
rect 43932 20750 43934 20802
rect 43986 20750 43988 20802
rect 43932 20132 43988 20750
rect 44156 21586 44212 21598
rect 44156 21534 44158 21586
rect 44210 21534 44212 21586
rect 44156 20690 44212 21534
rect 44380 20916 44436 21646
rect 44492 21588 44548 21598
rect 44492 21494 44548 21532
rect 44380 20850 44436 20860
rect 44156 20638 44158 20690
rect 44210 20638 44212 20690
rect 44156 20626 44212 20638
rect 44132 20412 44396 20422
rect 44188 20356 44236 20412
rect 44292 20356 44340 20412
rect 44132 20346 44396 20356
rect 43932 20066 43988 20076
rect 43260 20020 43316 20030
rect 43260 19908 43316 19964
rect 43820 20018 43876 20030
rect 43820 19966 43822 20018
rect 43874 19966 43876 20018
rect 43372 19908 43428 19918
rect 43260 19906 43428 19908
rect 43260 19854 43374 19906
rect 43426 19854 43428 19906
rect 43260 19852 43428 19854
rect 43372 19842 43428 19852
rect 42924 18274 42980 18284
rect 43260 19236 43316 19246
rect 43260 18340 43316 19180
rect 43820 18450 43876 19966
rect 44044 20020 44100 20030
rect 43932 19796 43988 19806
rect 43932 19458 43988 19740
rect 43932 19406 43934 19458
rect 43986 19406 43988 19458
rect 43932 19394 43988 19406
rect 44044 19236 44100 19964
rect 43820 18398 43822 18450
rect 43874 18398 43876 18450
rect 43820 18386 43876 18398
rect 43932 19180 44100 19236
rect 44492 20018 44548 20030
rect 44492 19966 44494 20018
rect 44546 19966 44548 20018
rect 43260 18274 43316 18284
rect 42924 17892 42980 17902
rect 42924 17780 42980 17836
rect 42364 17054 42366 17106
rect 42418 17054 42420 17106
rect 42364 17042 42420 17054
rect 42588 17724 42980 17780
rect 42252 16772 42308 16782
rect 42252 16100 42308 16716
rect 42364 16324 42420 16334
rect 42364 16230 42420 16268
rect 42476 16210 42532 16222
rect 42476 16158 42478 16210
rect 42530 16158 42532 16210
rect 42252 16098 42420 16100
rect 42252 16046 42254 16098
rect 42306 16046 42420 16098
rect 42252 16044 42420 16046
rect 42252 16034 42308 16044
rect 42028 15820 42196 15876
rect 41804 15428 41860 15438
rect 41804 15334 41860 15372
rect 41692 15092 41972 15148
rect 41804 14532 41860 14542
rect 41692 14530 41860 14532
rect 41692 14478 41806 14530
rect 41858 14478 41860 14530
rect 41692 14476 41860 14478
rect 41692 13186 41748 14476
rect 41804 14466 41860 14476
rect 41692 13134 41694 13186
rect 41746 13134 41748 13186
rect 41692 13122 41748 13134
rect 41916 13076 41972 15092
rect 41916 13010 41972 13020
rect 42028 11732 42084 15820
rect 42364 15538 42420 16044
rect 42364 15486 42366 15538
rect 42418 15486 42420 15538
rect 42364 15474 42420 15486
rect 42140 15316 42196 15326
rect 42476 15316 42532 16158
rect 42196 15260 42532 15316
rect 42140 15222 42196 15260
rect 42588 15148 42644 17724
rect 42924 17666 42980 17724
rect 42924 17614 42926 17666
rect 42978 17614 42980 17666
rect 42924 17602 42980 17614
rect 43148 17780 43204 17790
rect 43036 17220 43092 17230
rect 43036 16994 43092 17164
rect 43148 17108 43204 17724
rect 43932 17778 43988 19180
rect 44132 18844 44396 18854
rect 44188 18788 44236 18844
rect 44292 18788 44340 18844
rect 44132 18778 44396 18788
rect 44492 18676 44548 19966
rect 44492 18610 44548 18620
rect 44380 18452 44436 18462
rect 44604 18452 44660 23884
rect 44716 23716 44772 23726
rect 44716 23378 44772 23660
rect 44940 23714 44996 23726
rect 44940 23662 44942 23714
rect 44994 23662 44996 23714
rect 44716 23326 44718 23378
rect 44770 23326 44772 23378
rect 44716 23314 44772 23326
rect 44828 23492 44884 23502
rect 44940 23492 44996 23662
rect 44884 23436 44996 23492
rect 44828 22258 44884 23436
rect 44828 22206 44830 22258
rect 44882 22206 44884 22258
rect 44828 22194 44884 22206
rect 44828 21476 44884 21486
rect 44828 21382 44884 21420
rect 45052 21252 45108 23884
rect 45836 23940 45892 23950
rect 45724 23826 45780 23838
rect 45724 23774 45726 23826
rect 45778 23774 45780 23826
rect 45164 23716 45220 23726
rect 45388 23716 45444 23726
rect 45164 23714 45332 23716
rect 45164 23662 45166 23714
rect 45218 23662 45332 23714
rect 45164 23660 45332 23662
rect 45164 23650 45220 23660
rect 45276 23492 45332 23660
rect 45388 23714 45556 23716
rect 45388 23662 45390 23714
rect 45442 23662 45556 23714
rect 45388 23660 45556 23662
rect 45388 23650 45444 23660
rect 45500 23548 45556 23660
rect 45724 23604 45780 23774
rect 45836 23826 45892 23884
rect 45836 23774 45838 23826
rect 45890 23774 45892 23826
rect 45836 23762 45892 23774
rect 45948 23716 46004 24444
rect 46060 24434 46116 24444
rect 46284 24276 46340 25788
rect 46956 25730 47012 25788
rect 46956 25678 46958 25730
rect 47010 25678 47012 25730
rect 46956 25666 47012 25678
rect 47068 25620 47124 25630
rect 47068 25526 47124 25564
rect 46508 25396 46564 25406
rect 46508 25302 46564 25340
rect 47180 25284 47236 25294
rect 46956 25282 47236 25284
rect 46956 25230 47182 25282
rect 47234 25230 47236 25282
rect 46956 25228 47236 25230
rect 46620 24948 46676 24958
rect 46396 24724 46452 24734
rect 46396 24610 46452 24668
rect 46396 24558 46398 24610
rect 46450 24558 46452 24610
rect 46396 24546 46452 24558
rect 46060 24220 46340 24276
rect 46060 23938 46116 24220
rect 46508 24164 46564 24174
rect 46508 24050 46564 24108
rect 46508 23998 46510 24050
rect 46562 23998 46564 24050
rect 46508 23986 46564 23998
rect 46060 23886 46062 23938
rect 46114 23886 46116 23938
rect 46060 23874 46116 23886
rect 45948 23650 46004 23660
rect 45500 23492 45668 23548
rect 45724 23538 45780 23548
rect 45276 23426 45332 23436
rect 45276 23268 45332 23278
rect 45164 23154 45220 23166
rect 45164 23102 45166 23154
rect 45218 23102 45220 23154
rect 45164 22370 45220 23102
rect 45164 22318 45166 22370
rect 45218 22318 45220 22370
rect 45164 22260 45220 22318
rect 45164 21586 45220 22204
rect 45164 21534 45166 21586
rect 45218 21534 45220 21586
rect 45164 21522 45220 21534
rect 44828 21196 45108 21252
rect 44716 20132 44772 20142
rect 44716 19906 44772 20076
rect 44716 19854 44718 19906
rect 44770 19854 44772 19906
rect 44716 19842 44772 19854
rect 44828 19124 44884 21196
rect 44380 18358 44436 18396
rect 44492 18396 44660 18452
rect 44716 18450 44772 18462
rect 44716 18398 44718 18450
rect 44770 18398 44772 18450
rect 44156 18340 44212 18350
rect 44156 18246 44212 18284
rect 43932 17726 43934 17778
rect 43986 17726 43988 17778
rect 43932 17714 43988 17726
rect 43820 17668 43876 17678
rect 43148 17106 43652 17108
rect 43148 17054 43150 17106
rect 43202 17054 43652 17106
rect 43148 17052 43652 17054
rect 43148 17042 43204 17052
rect 43036 16942 43038 16994
rect 43090 16942 43092 16994
rect 43036 16930 43092 16942
rect 43596 16994 43652 17052
rect 43596 16942 43598 16994
rect 43650 16942 43652 16994
rect 43596 16930 43652 16942
rect 42700 16884 42756 16894
rect 42700 16790 42756 16828
rect 43372 16884 43428 16894
rect 43372 16882 43540 16884
rect 43372 16830 43374 16882
rect 43426 16830 43540 16882
rect 43372 16828 43540 16830
rect 43372 16818 43428 16828
rect 42924 16324 42980 16334
rect 42980 16268 43316 16324
rect 42924 15426 42980 16268
rect 43260 16210 43316 16268
rect 43260 16158 43262 16210
rect 43314 16158 43316 16210
rect 43260 16146 43316 16158
rect 43484 16100 43540 16828
rect 43372 16098 43540 16100
rect 43372 16046 43486 16098
rect 43538 16046 43540 16098
rect 43372 16044 43540 16046
rect 43372 15876 43428 16044
rect 43484 16034 43540 16044
rect 43820 15988 43876 17612
rect 44132 17276 44396 17286
rect 44188 17220 44236 17276
rect 44292 17220 44340 17276
rect 44132 17210 44396 17220
rect 43932 16994 43988 17006
rect 43932 16942 43934 16994
rect 43986 16942 43988 16994
rect 43932 16772 43988 16942
rect 43932 16706 43988 16716
rect 44156 16324 44212 16334
rect 44156 16210 44212 16268
rect 44156 16158 44158 16210
rect 44210 16158 44212 16210
rect 44156 16146 44212 16158
rect 43148 15820 43428 15876
rect 43708 15932 43876 15988
rect 43148 15538 43204 15820
rect 43148 15486 43150 15538
rect 43202 15486 43204 15538
rect 43148 15474 43204 15486
rect 43708 15538 43764 15932
rect 44132 15708 44396 15718
rect 44188 15652 44236 15708
rect 44292 15652 44340 15708
rect 44132 15642 44396 15652
rect 43708 15486 43710 15538
rect 43762 15486 43764 15538
rect 43708 15474 43764 15486
rect 44268 15540 44324 15550
rect 42924 15374 42926 15426
rect 42978 15374 42980 15426
rect 42924 15362 42980 15374
rect 43820 15426 43876 15438
rect 43820 15374 43822 15426
rect 43874 15374 43876 15426
rect 43260 15204 43316 15214
rect 43596 15204 43652 15214
rect 43260 15202 43652 15204
rect 43260 15150 43262 15202
rect 43314 15150 43598 15202
rect 43650 15150 43652 15202
rect 43260 15148 43652 15150
rect 42476 15092 42532 15102
rect 42588 15092 42756 15148
rect 43260 15138 43316 15148
rect 43596 15138 43652 15148
rect 43820 15204 43876 15374
rect 44268 15426 44324 15484
rect 44268 15374 44270 15426
rect 44322 15374 44324 15426
rect 44268 15362 44324 15374
rect 43820 15138 43876 15148
rect 42476 14998 42532 15036
rect 42476 13746 42532 13758
rect 42476 13694 42478 13746
rect 42530 13694 42532 13746
rect 42476 13524 42532 13694
rect 42476 13458 42532 13468
rect 42476 12178 42532 12190
rect 42476 12126 42478 12178
rect 42530 12126 42532 12178
rect 42476 11844 42532 12126
rect 42700 11954 42756 15092
rect 43932 14644 43988 14654
rect 43932 14418 43988 14588
rect 44268 14532 44324 14542
rect 44268 14438 44324 14476
rect 43932 14366 43934 14418
rect 43986 14366 43988 14418
rect 42700 11902 42702 11954
rect 42754 11902 42756 11954
rect 42700 11890 42756 11902
rect 42812 14196 42868 14206
rect 42476 11778 42532 11788
rect 42028 11666 42084 11676
rect 41804 11172 41860 11182
rect 41356 10108 41636 10164
rect 41692 11170 41860 11172
rect 41692 11118 41806 11170
rect 41858 11118 41860 11170
rect 41692 11116 41860 11118
rect 41692 10724 41748 11116
rect 41804 11106 41860 11116
rect 42140 11172 42196 11182
rect 42588 11172 42644 11182
rect 42140 11170 42644 11172
rect 42140 11118 42142 11170
rect 42194 11118 42590 11170
rect 42642 11118 42644 11170
rect 42140 11116 42644 11118
rect 41692 10164 41748 10668
rect 41804 10836 41860 10846
rect 42140 10836 42196 11116
rect 41860 10780 42196 10836
rect 41804 10610 41860 10780
rect 42588 10724 42644 11116
rect 42700 10724 42756 10734
rect 42588 10722 42756 10724
rect 42588 10670 42702 10722
rect 42754 10670 42756 10722
rect 42588 10668 42756 10670
rect 42700 10658 42756 10668
rect 41804 10558 41806 10610
rect 41858 10558 41860 10610
rect 41804 10546 41860 10558
rect 42252 10610 42308 10622
rect 42252 10558 42254 10610
rect 42306 10558 42308 10610
rect 42252 10388 42308 10558
rect 41692 10108 41972 10164
rect 41020 9828 41076 9838
rect 41020 9826 41188 9828
rect 41020 9774 41022 9826
rect 41074 9774 41188 9826
rect 41020 9772 41188 9774
rect 41020 9762 41076 9772
rect 40684 9716 40740 9726
rect 40684 9622 40740 9660
rect 39900 8370 39956 8428
rect 39900 8318 39902 8370
rect 39954 8318 39956 8370
rect 39452 7634 39508 7644
rect 38780 7534 38782 7586
rect 38834 7534 38836 7586
rect 38780 7522 38836 7534
rect 39340 7586 39396 7598
rect 39340 7534 39342 7586
rect 39394 7534 39396 7586
rect 38556 7420 38724 7476
rect 39116 7474 39172 7486
rect 39116 7422 39118 7474
rect 39170 7422 39172 7474
rect 38556 7028 38612 7420
rect 38668 7252 38724 7262
rect 39116 7252 39172 7422
rect 38668 7250 39172 7252
rect 38668 7198 38670 7250
rect 38722 7198 39172 7250
rect 38668 7196 39172 7198
rect 38668 7186 38724 7196
rect 38556 6972 38836 7028
rect 38780 6916 38836 6972
rect 38556 6692 38612 6702
rect 38780 6692 38836 6860
rect 39340 6804 39396 7534
rect 39004 6748 39396 6804
rect 39788 6914 39844 6926
rect 39788 6862 39790 6914
rect 39842 6862 39844 6914
rect 38892 6692 38948 6702
rect 38556 6690 38724 6692
rect 38556 6638 38558 6690
rect 38610 6638 38724 6690
rect 38556 6636 38724 6638
rect 38780 6690 38948 6692
rect 38780 6638 38894 6690
rect 38946 6638 38948 6690
rect 38780 6636 38948 6638
rect 38556 6626 38612 6636
rect 38668 6020 38724 6636
rect 38892 6626 38948 6636
rect 39004 6130 39060 6748
rect 39004 6078 39006 6130
rect 39058 6078 39060 6130
rect 39004 6066 39060 6078
rect 38668 5926 38724 5964
rect 39788 5908 39844 6862
rect 39900 6690 39956 8318
rect 40012 8876 40628 8932
rect 40796 9602 40852 9614
rect 40796 9550 40798 9602
rect 40850 9550 40852 9602
rect 40012 7698 40068 8876
rect 40236 8708 40292 8718
rect 40012 7646 40014 7698
rect 40066 7646 40068 7698
rect 40012 7634 40068 7646
rect 40124 8652 40236 8708
rect 40124 7474 40180 8652
rect 40236 8642 40292 8652
rect 40796 8708 40852 9550
rect 40908 9268 40964 9278
rect 40908 9174 40964 9212
rect 40796 8642 40852 8652
rect 41132 8484 41188 9772
rect 41244 9154 41300 9166
rect 41244 9102 41246 9154
rect 41298 9102 41300 9154
rect 41244 9044 41300 9102
rect 41244 8978 41300 8988
rect 41244 8484 41300 8494
rect 41132 8482 41300 8484
rect 41132 8430 41246 8482
rect 41298 8430 41300 8482
rect 41132 8428 41300 8430
rect 41244 8418 41300 8428
rect 40236 8146 40292 8158
rect 40236 8094 40238 8146
rect 40290 8094 40292 8146
rect 40236 7924 40292 8094
rect 40236 7858 40292 7868
rect 41132 7700 41188 7710
rect 41356 7700 41412 10108
rect 41804 9828 41860 9838
rect 41692 9716 41748 9726
rect 41692 9622 41748 9660
rect 41468 9604 41524 9614
rect 41468 9510 41524 9548
rect 41580 9602 41636 9614
rect 41580 9550 41582 9602
rect 41634 9550 41636 9602
rect 41580 8036 41636 9550
rect 41804 9154 41860 9772
rect 41804 9102 41806 9154
rect 41858 9102 41860 9154
rect 41804 8820 41860 9102
rect 41804 8754 41860 8764
rect 41580 7970 41636 7980
rect 41132 7698 41412 7700
rect 41132 7646 41134 7698
rect 41186 7646 41412 7698
rect 41132 7644 41412 7646
rect 41132 7634 41188 7644
rect 41580 7586 41636 7598
rect 41580 7534 41582 7586
rect 41634 7534 41636 7586
rect 40124 7422 40126 7474
rect 40178 7422 40180 7474
rect 40124 7410 40180 7422
rect 40908 7476 40964 7486
rect 40908 7382 40964 7420
rect 41468 7474 41524 7486
rect 41468 7422 41470 7474
rect 41522 7422 41524 7474
rect 39900 6638 39902 6690
rect 39954 6638 39956 6690
rect 39900 6626 39956 6638
rect 40796 6468 40852 6478
rect 40796 6374 40852 6412
rect 41468 6244 41524 7422
rect 41132 6188 41524 6244
rect 40236 5908 40292 5918
rect 39788 5906 39956 5908
rect 39788 5854 39790 5906
rect 39842 5854 39956 5906
rect 39788 5852 39956 5854
rect 39788 5842 39844 5852
rect 38556 5796 38612 5806
rect 38556 4900 38612 5740
rect 39116 5796 39172 5806
rect 38780 5124 38836 5134
rect 38780 5030 38836 5068
rect 38556 3666 38612 4844
rect 38892 4452 38948 4462
rect 38892 4358 38948 4396
rect 39116 4226 39172 5740
rect 39676 5684 39732 5694
rect 39228 5010 39284 5022
rect 39228 4958 39230 5010
rect 39282 4958 39284 5010
rect 39228 4788 39284 4958
rect 39676 5010 39732 5628
rect 39676 4958 39678 5010
rect 39730 4958 39732 5010
rect 39676 4946 39732 4958
rect 39900 5122 39956 5852
rect 40236 5814 40292 5852
rect 41020 5796 41076 5806
rect 41020 5702 41076 5740
rect 41132 5346 41188 6188
rect 41244 6020 41300 6030
rect 41580 6020 41636 7534
rect 41916 6916 41972 10108
rect 42140 9940 42196 9950
rect 42028 9714 42084 9726
rect 42028 9662 42030 9714
rect 42082 9662 42084 9714
rect 42028 9268 42084 9662
rect 42140 9714 42196 9884
rect 42140 9662 42142 9714
rect 42194 9662 42196 9714
rect 42140 9650 42196 9662
rect 42028 9202 42084 9212
rect 42252 9492 42308 10332
rect 42812 10276 42868 14140
rect 43484 13860 43540 13898
rect 43484 13794 43540 13804
rect 43484 13636 43540 13646
rect 42924 12068 42980 12078
rect 42924 10834 42980 12012
rect 43484 11506 43540 13580
rect 43932 13524 43988 14366
rect 44132 14140 44396 14150
rect 44188 14084 44236 14140
rect 44292 14084 44340 14140
rect 44132 14074 44396 14084
rect 43932 13458 43988 13468
rect 43596 13300 43652 13310
rect 43596 13074 43652 13244
rect 43596 13022 43598 13074
rect 43650 13022 43652 13074
rect 43596 13010 43652 13022
rect 44268 13300 44324 13310
rect 44492 13300 44548 18396
rect 44716 17892 44772 18398
rect 44716 17826 44772 17836
rect 44828 17554 44884 19068
rect 44828 17502 44830 17554
rect 44882 17502 44884 17554
rect 44828 17490 44884 17502
rect 44940 20690 44996 20702
rect 44940 20638 44942 20690
rect 44994 20638 44996 20690
rect 44940 20244 44996 20638
rect 44940 17220 44996 20188
rect 45164 19348 45220 19358
rect 45164 19254 45220 19292
rect 45164 18340 45220 18350
rect 45164 18246 45220 18284
rect 44716 17164 44996 17220
rect 45164 17442 45220 17454
rect 45164 17390 45166 17442
rect 45218 17390 45220 17442
rect 44604 15540 44660 15550
rect 44604 15446 44660 15484
rect 44716 15148 44772 17164
rect 45164 16772 45220 17390
rect 45276 17220 45332 23212
rect 45612 23268 45668 23492
rect 45612 23202 45668 23212
rect 46508 23268 46564 23278
rect 45388 23156 45444 23166
rect 45388 21700 45444 23100
rect 46060 23042 46116 23054
rect 46060 22990 46062 23042
rect 46114 22990 46116 23042
rect 46060 22484 46116 22990
rect 46396 22484 46452 22494
rect 46060 22428 46340 22484
rect 45500 22372 45556 22382
rect 45500 22278 45556 22316
rect 45724 22372 45780 22382
rect 45388 21644 45556 21700
rect 45388 21474 45444 21486
rect 45388 21422 45390 21474
rect 45442 21422 45444 21474
rect 45388 20132 45444 21422
rect 45388 20066 45444 20076
rect 45276 17106 45332 17164
rect 45276 17054 45278 17106
rect 45330 17054 45332 17106
rect 45276 17042 45332 17054
rect 45164 16706 45220 16716
rect 44940 16660 44996 16670
rect 44940 15316 44996 16604
rect 45276 16100 45332 16110
rect 45276 16006 45332 16044
rect 45500 15986 45556 21644
rect 45724 20692 45780 22316
rect 45836 22260 45892 22270
rect 46172 22260 46228 22270
rect 45892 22258 46228 22260
rect 45892 22206 46174 22258
rect 46226 22206 46228 22258
rect 45892 22204 46228 22206
rect 45836 22166 45892 22204
rect 46172 22194 46228 22204
rect 46284 22146 46340 22428
rect 46284 22094 46286 22146
rect 46338 22094 46340 22146
rect 46284 22036 46340 22094
rect 46060 21980 46340 22036
rect 46060 21700 46116 21980
rect 46396 21924 46452 22428
rect 46508 22370 46564 23212
rect 46508 22318 46510 22370
rect 46562 22318 46564 22370
rect 46508 22306 46564 22318
rect 46620 22260 46676 24892
rect 46956 24724 47012 25228
rect 47180 25218 47236 25228
rect 46956 24658 47012 24668
rect 47292 23940 47348 26012
rect 47740 25618 47796 26852
rect 48188 26964 48244 27002
rect 48188 26404 48244 26908
rect 47852 26348 48244 26404
rect 48300 26850 48356 27692
rect 48860 27682 48916 27692
rect 48412 27188 48468 27198
rect 48412 27076 48468 27132
rect 48524 27076 48580 27086
rect 48412 27074 48580 27076
rect 48412 27022 48526 27074
rect 48578 27022 48580 27074
rect 48412 27020 48580 27022
rect 48524 27010 48580 27020
rect 48972 26908 49028 28700
rect 49084 27298 49140 30942
rect 49420 30994 49476 31006
rect 49420 30942 49422 30994
rect 49474 30942 49476 30994
rect 49308 30884 49364 30894
rect 49308 30790 49364 30828
rect 49196 30212 49252 30222
rect 49196 29204 49252 30156
rect 49196 28866 49252 29148
rect 49196 28814 49198 28866
rect 49250 28814 49252 28866
rect 49196 28802 49252 28814
rect 49420 30098 49476 30942
rect 49420 30046 49422 30098
rect 49474 30046 49476 30098
rect 49308 28196 49364 28206
rect 49308 28082 49364 28140
rect 49308 28030 49310 28082
rect 49362 28030 49364 28082
rect 49308 28018 49364 28030
rect 49420 28084 49476 30046
rect 50092 29426 50148 31612
rect 50204 29538 50260 31948
rect 50652 31556 50708 32620
rect 50876 32450 50932 32462
rect 51212 32452 51268 33180
rect 51324 33236 51380 33246
rect 51324 33142 51380 33180
rect 51436 32452 51492 32462
rect 50876 32398 50878 32450
rect 50930 32398 50932 32450
rect 50876 32004 50932 32398
rect 50876 31938 50932 31948
rect 51100 32450 51492 32452
rect 51100 32398 51438 32450
rect 51490 32398 51492 32450
rect 51100 32396 51492 32398
rect 50876 31556 50932 31566
rect 50652 31554 50932 31556
rect 50652 31502 50878 31554
rect 50930 31502 50932 31554
rect 50652 31500 50932 31502
rect 50652 30436 50708 31500
rect 50876 31490 50932 31500
rect 50764 30772 50820 30782
rect 50764 30678 50820 30716
rect 50652 30370 50708 30380
rect 50428 30212 50484 30222
rect 50428 30118 50484 30156
rect 50204 29486 50206 29538
rect 50258 29486 50260 29538
rect 50204 29474 50260 29486
rect 50092 29374 50094 29426
rect 50146 29374 50148 29426
rect 50092 29362 50148 29374
rect 50316 29316 50372 29326
rect 49532 29204 49588 29214
rect 49588 29148 49700 29204
rect 49532 29138 49588 29148
rect 49532 28084 49588 28094
rect 49420 28082 49588 28084
rect 49420 28030 49534 28082
rect 49586 28030 49588 28082
rect 49420 28028 49588 28030
rect 49532 28018 49588 28028
rect 49196 27914 49252 27926
rect 49196 27862 49198 27914
rect 49250 27862 49252 27914
rect 49196 27412 49252 27862
rect 49196 27356 49588 27412
rect 49084 27246 49086 27298
rect 49138 27246 49140 27298
rect 49084 27234 49140 27246
rect 49532 27188 49588 27356
rect 49420 27132 49588 27188
rect 49308 27076 49364 27086
rect 48300 26798 48302 26850
rect 48354 26798 48356 26850
rect 47852 25956 47908 26348
rect 47964 26180 48020 26190
rect 48300 26180 48356 26798
rect 48020 26124 48356 26180
rect 48748 26852 49028 26908
rect 49196 27020 49308 27076
rect 49196 26962 49252 27020
rect 49308 27010 49364 27020
rect 49196 26910 49198 26962
rect 49250 26910 49252 26962
rect 49196 26898 49252 26910
rect 49420 26908 49476 27132
rect 49644 27076 49700 29148
rect 49980 28868 50036 28878
rect 49756 28754 49812 28766
rect 49756 28702 49758 28754
rect 49810 28702 49812 28754
rect 49756 28082 49812 28702
rect 49980 28642 50036 28812
rect 50316 28754 50372 29260
rect 50316 28702 50318 28754
rect 50370 28702 50372 28754
rect 50316 28690 50372 28702
rect 49980 28590 49982 28642
rect 50034 28590 50036 28642
rect 49980 28578 50036 28590
rect 49756 28030 49758 28082
rect 49810 28030 49812 28082
rect 49756 28018 49812 28030
rect 50540 27972 50596 27982
rect 50204 27858 50260 27870
rect 50204 27806 50206 27858
rect 50258 27806 50260 27858
rect 50204 27636 50260 27806
rect 50316 27860 50372 27870
rect 50316 27766 50372 27804
rect 50540 27858 50596 27916
rect 50764 27860 50820 27870
rect 50540 27806 50542 27858
rect 50594 27806 50596 27858
rect 50540 27794 50596 27806
rect 50652 27804 50764 27860
rect 50204 27570 50260 27580
rect 50652 27298 50708 27804
rect 50764 27794 50820 27804
rect 50876 27858 50932 27870
rect 50876 27806 50878 27858
rect 50930 27806 50932 27858
rect 50876 27636 50932 27806
rect 50876 27570 50932 27580
rect 50652 27246 50654 27298
rect 50706 27246 50708 27298
rect 50652 27234 50708 27246
rect 49644 27010 49700 27020
rect 49084 26852 49140 26862
rect 48748 26850 49140 26852
rect 48748 26798 49086 26850
rect 49138 26798 49140 26850
rect 48748 26796 49140 26798
rect 47964 26086 48020 26124
rect 47852 25900 48020 25956
rect 47740 25566 47742 25618
rect 47794 25566 47796 25618
rect 47740 25554 47796 25566
rect 47852 25508 47908 25518
rect 47852 24722 47908 25452
rect 47852 24670 47854 24722
rect 47906 24670 47908 24722
rect 47068 23884 47348 23940
rect 47404 24610 47460 24622
rect 47404 24558 47406 24610
rect 47458 24558 47460 24610
rect 46844 23716 46900 23726
rect 46844 23622 46900 23660
rect 46956 23044 47012 23054
rect 46956 22950 47012 22988
rect 46620 22194 46676 22204
rect 46732 22820 46788 22830
rect 46732 22036 46788 22764
rect 47068 22372 47124 23884
rect 47404 23828 47460 24558
rect 47628 24612 47684 24622
rect 47628 24518 47684 24556
rect 47404 23762 47460 23772
rect 47628 24164 47684 24174
rect 47180 23714 47236 23726
rect 47180 23662 47182 23714
rect 47234 23662 47236 23714
rect 47180 23268 47236 23662
rect 47628 23378 47684 24108
rect 47852 24162 47908 24670
rect 47852 24110 47854 24162
rect 47906 24110 47908 24162
rect 47852 24098 47908 24110
rect 47964 23940 48020 25900
rect 48188 25732 48244 25742
rect 48188 25282 48244 25676
rect 48636 25508 48692 25518
rect 48636 25414 48692 25452
rect 48188 25230 48190 25282
rect 48242 25230 48244 25282
rect 48188 24948 48244 25230
rect 48188 24882 48244 24892
rect 48636 24724 48692 24734
rect 48188 24722 48692 24724
rect 48188 24670 48638 24722
rect 48690 24670 48692 24722
rect 48188 24668 48692 24670
rect 48188 24610 48244 24668
rect 48636 24658 48692 24668
rect 48188 24558 48190 24610
rect 48242 24558 48244 24610
rect 48188 24546 48244 24558
rect 48748 24612 48804 26796
rect 49084 26786 49140 26796
rect 49308 26852 49476 26908
rect 49532 26964 49588 26974
rect 49308 26628 49364 26852
rect 49084 26402 49140 26414
rect 49084 26350 49086 26402
rect 49138 26350 49140 26402
rect 48972 26178 49028 26190
rect 48972 26126 48974 26178
rect 49026 26126 49028 26178
rect 48860 24612 48916 24622
rect 48748 24610 48916 24612
rect 48748 24558 48862 24610
rect 48914 24558 48916 24610
rect 48748 24556 48916 24558
rect 48860 24546 48916 24556
rect 48636 24164 48692 24174
rect 48524 24108 48636 24164
rect 48524 24050 48580 24108
rect 48636 24098 48692 24108
rect 48524 23998 48526 24050
rect 48578 23998 48580 24050
rect 48524 23986 48580 23998
rect 47628 23326 47630 23378
rect 47682 23326 47684 23378
rect 47628 23314 47684 23326
rect 47852 23884 48020 23940
rect 48188 23938 48244 23950
rect 48188 23886 48190 23938
rect 48242 23886 48244 23938
rect 47180 23202 47236 23212
rect 47404 23266 47460 23278
rect 47404 23214 47406 23266
rect 47458 23214 47460 23266
rect 46284 21868 46452 21924
rect 46508 21980 46788 22036
rect 46956 22316 47124 22372
rect 47292 23154 47348 23166
rect 47292 23102 47294 23154
rect 47346 23102 47348 23154
rect 46172 21812 46228 21822
rect 46172 21718 46228 21756
rect 46060 21634 46116 21644
rect 45836 21586 45892 21598
rect 45836 21534 45838 21586
rect 45890 21534 45892 21586
rect 45836 20804 45892 21534
rect 45948 21586 46004 21598
rect 45948 21534 45950 21586
rect 46002 21534 46004 21586
rect 45948 21364 46004 21534
rect 46284 21586 46340 21868
rect 46284 21534 46286 21586
rect 46338 21534 46340 21586
rect 45948 21140 46004 21308
rect 45948 21074 46004 21084
rect 46060 21474 46116 21486
rect 46060 21422 46062 21474
rect 46114 21422 46116 21474
rect 46060 21028 46116 21422
rect 46060 20972 46228 21028
rect 46060 20804 46116 20814
rect 45836 20802 46116 20804
rect 45836 20750 46062 20802
rect 46114 20750 46116 20802
rect 45836 20748 46116 20750
rect 46060 20692 46116 20748
rect 45724 20636 45892 20692
rect 45836 19236 45892 20636
rect 46060 20626 46116 20636
rect 46172 20580 46228 20972
rect 46172 20514 46228 20524
rect 46284 20244 46340 21534
rect 46396 21700 46452 21710
rect 46396 20914 46452 21644
rect 46396 20862 46398 20914
rect 46450 20862 46452 20914
rect 46396 20850 46452 20862
rect 45612 19180 45892 19236
rect 45948 20188 46340 20244
rect 45612 18340 45668 19180
rect 45724 19012 45780 19050
rect 45948 19012 46004 20188
rect 46508 20020 46564 21980
rect 46844 21812 46900 21822
rect 46620 21810 46900 21812
rect 46620 21758 46846 21810
rect 46898 21758 46900 21810
rect 46620 21756 46900 21758
rect 46620 20692 46676 21756
rect 46844 21746 46900 21756
rect 46732 21586 46788 21598
rect 46732 21534 46734 21586
rect 46786 21534 46788 21586
rect 46732 21252 46788 21534
rect 46844 21364 46900 21374
rect 46844 21270 46900 21308
rect 46732 21186 46788 21196
rect 46956 21140 47012 22316
rect 47068 22148 47124 22158
rect 47180 22148 47236 22158
rect 47068 22146 47180 22148
rect 47068 22094 47070 22146
rect 47122 22094 47180 22146
rect 47068 22092 47180 22094
rect 47068 21588 47124 22092
rect 47180 22082 47236 22092
rect 47292 21700 47348 23102
rect 47404 23044 47460 23214
rect 47404 22484 47460 22988
rect 47404 22418 47460 22428
rect 47404 22260 47460 22270
rect 47404 22166 47460 22204
rect 47740 22146 47796 22158
rect 47740 22094 47742 22146
rect 47794 22094 47796 22146
rect 47740 21924 47796 22094
rect 47852 22148 47908 23884
rect 47964 23716 48020 23726
rect 47964 23378 48020 23660
rect 47964 23326 47966 23378
rect 48018 23326 48020 23378
rect 47964 23314 48020 23326
rect 48188 23268 48244 23886
rect 48188 23202 48244 23212
rect 48300 23716 48356 23726
rect 48076 23156 48132 23166
rect 48076 23062 48132 23100
rect 48188 23044 48244 23054
rect 48188 22950 48244 22988
rect 48300 22820 48356 23660
rect 48188 22764 48356 22820
rect 48524 23044 48580 23054
rect 48076 22708 48132 22718
rect 47852 22082 47908 22092
rect 47964 22260 48020 22270
rect 47404 21868 47796 21924
rect 47404 21700 47460 21868
rect 47068 21522 47124 21532
rect 47180 21698 47460 21700
rect 47180 21646 47406 21698
rect 47458 21646 47460 21698
rect 47180 21644 47460 21646
rect 47180 21364 47236 21644
rect 47404 21634 47460 21644
rect 47516 21700 47572 21710
rect 47516 21606 47572 21644
rect 47964 21698 48020 22204
rect 48076 22258 48132 22652
rect 48076 22206 48078 22258
rect 48130 22206 48132 22258
rect 48076 22194 48132 22206
rect 47964 21646 47966 21698
rect 48018 21646 48020 21698
rect 47964 21634 48020 21646
rect 48076 21700 48132 21710
rect 48076 21606 48132 21644
rect 47852 21476 47908 21486
rect 48076 21476 48132 21486
rect 46844 21084 47012 21140
rect 47068 21308 47236 21364
rect 47516 21364 47572 21374
rect 47516 21362 47684 21364
rect 47516 21310 47518 21362
rect 47570 21310 47684 21362
rect 47516 21308 47684 21310
rect 46620 20598 46676 20636
rect 46732 20690 46788 20702
rect 46732 20638 46734 20690
rect 46786 20638 46788 20690
rect 46620 20020 46676 20030
rect 46564 20018 46676 20020
rect 46564 19966 46622 20018
rect 46674 19966 46676 20018
rect 46564 19964 46676 19966
rect 46508 19926 46564 19964
rect 46620 19954 46676 19964
rect 45724 18946 45780 18956
rect 45836 19010 46004 19012
rect 45836 18958 45950 19010
rect 46002 18958 46004 19010
rect 45836 18956 46004 18958
rect 45724 18340 45780 18350
rect 45612 18338 45780 18340
rect 45612 18286 45726 18338
rect 45778 18286 45780 18338
rect 45612 18284 45780 18286
rect 45724 18116 45780 18284
rect 45612 17668 45668 17678
rect 45724 17668 45780 18060
rect 45612 17666 45780 17668
rect 45612 17614 45614 17666
rect 45666 17614 45780 17666
rect 45612 17612 45780 17614
rect 45612 17602 45668 17612
rect 45724 17442 45780 17454
rect 45724 17390 45726 17442
rect 45778 17390 45780 17442
rect 45612 16994 45668 17006
rect 45612 16942 45614 16994
rect 45666 16942 45668 16994
rect 45612 16660 45668 16942
rect 45724 16996 45780 17390
rect 45724 16930 45780 16940
rect 45612 16594 45668 16604
rect 45500 15934 45502 15986
rect 45554 15934 45556 15986
rect 45500 15876 45556 15934
rect 45500 15810 45556 15820
rect 45724 16098 45780 16110
rect 45724 16046 45726 16098
rect 45778 16046 45780 16098
rect 45724 15988 45780 16046
rect 45164 15652 45220 15662
rect 44940 15314 45108 15316
rect 44940 15262 44942 15314
rect 44994 15262 45108 15314
rect 44940 15260 45108 15262
rect 44940 15250 44996 15260
rect 44324 13244 44548 13300
rect 44604 15092 44772 15148
rect 44604 13746 44660 15092
rect 44940 14642 44996 14654
rect 44940 14590 44942 14642
rect 44994 14590 44996 14642
rect 44940 13860 44996 14590
rect 44940 13794 44996 13804
rect 44604 13694 44606 13746
rect 44658 13694 44660 13746
rect 44268 12962 44324 13244
rect 44604 13076 44660 13694
rect 44716 13076 44772 13086
rect 44604 13020 44716 13076
rect 44716 13010 44772 13020
rect 44268 12910 44270 12962
rect 44322 12910 44324 12962
rect 44268 12898 44324 12910
rect 43932 12738 43988 12750
rect 43932 12686 43934 12738
rect 43986 12686 43988 12738
rect 43820 12178 43876 12190
rect 43820 12126 43822 12178
rect 43874 12126 43876 12178
rect 43820 12068 43876 12126
rect 43820 12002 43876 12012
rect 43484 11454 43486 11506
rect 43538 11454 43540 11506
rect 43260 11284 43316 11294
rect 42924 10782 42926 10834
rect 42978 10782 42980 10834
rect 42924 10770 42980 10782
rect 43036 11170 43092 11182
rect 43036 11118 43038 11170
rect 43090 11118 43092 11170
rect 42812 10210 42868 10220
rect 42812 10052 42868 10062
rect 42812 9826 42868 9996
rect 43036 10052 43092 11118
rect 43260 10834 43316 11228
rect 43260 10782 43262 10834
rect 43314 10782 43316 10834
rect 43260 10770 43316 10782
rect 43036 9986 43092 9996
rect 43148 10610 43204 10622
rect 43148 10558 43150 10610
rect 43202 10558 43204 10610
rect 42812 9774 42814 9826
rect 42866 9774 42868 9826
rect 42812 9762 42868 9774
rect 42028 9044 42084 9054
rect 42252 9044 42308 9436
rect 42028 9042 42308 9044
rect 42028 8990 42030 9042
rect 42082 8990 42308 9042
rect 42028 8988 42308 8990
rect 42364 9602 42420 9614
rect 42364 9550 42366 9602
rect 42418 9550 42420 9602
rect 42028 8978 42084 8988
rect 42364 8484 42420 9550
rect 42476 9604 42532 9614
rect 42700 9604 42756 9614
rect 42476 8820 42532 9548
rect 42588 9548 42700 9604
rect 42588 9156 42644 9548
rect 42700 9510 42756 9548
rect 43148 9604 43204 10558
rect 43148 9510 43204 9548
rect 43260 10498 43316 10510
rect 43260 10446 43262 10498
rect 43314 10446 43316 10498
rect 42588 9042 42644 9100
rect 42588 8990 42590 9042
rect 42642 8990 42644 9042
rect 42588 8978 42644 8990
rect 43036 9044 43092 9054
rect 43036 8950 43092 8988
rect 43036 8820 43092 8830
rect 42476 8764 42644 8820
rect 42364 8428 42532 8484
rect 42140 8146 42196 8158
rect 42140 8094 42142 8146
rect 42194 8094 42196 8146
rect 42028 6916 42084 6926
rect 41916 6860 42028 6916
rect 42028 6850 42084 6860
rect 42140 6692 42196 8094
rect 42364 8036 42420 8046
rect 42364 7474 42420 7980
rect 42364 7422 42366 7474
rect 42418 7422 42420 7474
rect 42364 7410 42420 7422
rect 42476 6804 42532 8428
rect 42588 8258 42644 8764
rect 42588 8206 42590 8258
rect 42642 8206 42644 8258
rect 42588 7700 42644 8206
rect 42588 7634 42644 7644
rect 42476 6738 42532 6748
rect 42812 7362 42868 7374
rect 42812 7310 42814 7362
rect 42866 7310 42868 7362
rect 42140 6626 42196 6636
rect 42364 6690 42420 6702
rect 42364 6638 42366 6690
rect 42418 6638 42420 6690
rect 41300 5964 41636 6020
rect 41692 6580 41748 6590
rect 41244 5926 41300 5964
rect 41692 5796 41748 6524
rect 42364 6580 42420 6638
rect 42364 6514 42420 6524
rect 42140 6468 42196 6478
rect 41692 5730 41748 5740
rect 41916 6466 42196 6468
rect 41916 6414 42142 6466
rect 42194 6414 42196 6466
rect 41916 6412 42196 6414
rect 41132 5294 41134 5346
rect 41186 5294 41188 5346
rect 41132 5282 41188 5294
rect 41804 5236 41860 5246
rect 39900 5070 39902 5122
rect 39954 5070 39956 5122
rect 39900 5012 39956 5070
rect 39900 4946 39956 4956
rect 40348 5124 40404 5134
rect 40348 5010 40404 5068
rect 40684 5124 40740 5134
rect 40684 5030 40740 5068
rect 41132 5068 41524 5124
rect 40348 4958 40350 5010
rect 40402 4958 40404 5010
rect 40348 4946 40404 4958
rect 41020 5012 41076 5022
rect 41020 4918 41076 4956
rect 41132 5010 41188 5068
rect 41132 4958 41134 5010
rect 41186 4958 41188 5010
rect 41132 4946 41188 4958
rect 41468 5012 41524 5068
rect 41692 5012 41748 5022
rect 41468 5010 41748 5012
rect 41468 4958 41694 5010
rect 41746 4958 41748 5010
rect 41468 4956 41748 4958
rect 41692 4946 41748 4956
rect 39228 4722 39284 4732
rect 40236 4900 40292 4910
rect 40124 4676 40180 4686
rect 40124 4450 40180 4620
rect 40236 4562 40292 4844
rect 40236 4510 40238 4562
rect 40290 4510 40292 4562
rect 40236 4498 40292 4510
rect 41468 4676 41524 4686
rect 40124 4398 40126 4450
rect 40178 4398 40180 4450
rect 40124 4386 40180 4398
rect 39340 4340 39396 4350
rect 39340 4246 39396 4284
rect 40460 4340 40516 4350
rect 40460 4246 40516 4284
rect 41132 4340 41188 4350
rect 41132 4246 41188 4284
rect 39116 4174 39118 4226
rect 39170 4174 39172 4226
rect 39116 4162 39172 4174
rect 40796 4228 40852 4238
rect 41468 4228 41524 4620
rect 40796 3778 40852 4172
rect 41244 4226 41524 4228
rect 41244 4174 41470 4226
rect 41522 4174 41524 4226
rect 41244 4172 41524 4174
rect 41244 4116 41300 4172
rect 41468 4162 41524 4172
rect 40796 3726 40798 3778
rect 40850 3726 40852 3778
rect 40796 3714 40852 3726
rect 41020 4060 41300 4116
rect 38556 3614 38558 3666
rect 38610 3614 38612 3666
rect 38556 3602 38612 3614
rect 41020 3442 41076 4060
rect 41132 3666 41188 3678
rect 41132 3614 41134 3666
rect 41186 3614 41188 3666
rect 41132 3556 41188 3614
rect 41804 3668 41860 5180
rect 41916 5122 41972 6412
rect 42140 6402 42196 6412
rect 42476 5908 42532 5918
rect 42476 5814 42532 5852
rect 41916 5070 41918 5122
rect 41970 5070 41972 5122
rect 41916 5058 41972 5070
rect 42364 5124 42420 5134
rect 42364 5010 42420 5068
rect 42364 4958 42366 5010
rect 42418 4958 42420 5010
rect 42364 4946 42420 4958
rect 42700 4900 42756 4910
rect 42700 4806 42756 4844
rect 42812 4676 42868 7310
rect 43036 6802 43092 8764
rect 43260 8708 43316 10446
rect 43484 10164 43540 11454
rect 43596 11732 43652 11742
rect 43596 10612 43652 11676
rect 43932 11284 43988 12686
rect 44132 12572 44396 12582
rect 44188 12516 44236 12572
rect 44292 12516 44340 12572
rect 44132 12506 44396 12516
rect 44044 12404 44100 12414
rect 44044 12310 44100 12348
rect 45052 12404 45108 15260
rect 45164 15314 45220 15596
rect 45724 15540 45780 15932
rect 45724 15474 45780 15484
rect 45836 15316 45892 18956
rect 45948 18946 46004 18956
rect 46060 19908 46116 19918
rect 46060 19012 46116 19852
rect 45948 17668 46004 17678
rect 45948 17574 46004 17612
rect 45948 17220 46004 17230
rect 45948 17106 46004 17164
rect 45948 17054 45950 17106
rect 46002 17054 46004 17106
rect 45948 17042 46004 17054
rect 46060 16884 46116 18956
rect 46284 19124 46340 19134
rect 46620 19124 46676 19134
rect 46732 19124 46788 20638
rect 46284 19122 46732 19124
rect 46284 19070 46286 19122
rect 46338 19070 46622 19122
rect 46674 19070 46732 19122
rect 46284 19068 46732 19070
rect 46284 18450 46340 19068
rect 46620 19058 46676 19068
rect 46732 19030 46788 19068
rect 46844 18900 46900 21084
rect 46508 18844 46900 18900
rect 46956 19236 47012 19246
rect 46956 19122 47012 19180
rect 46956 19070 46958 19122
rect 47010 19070 47012 19122
rect 46508 18564 46564 18844
rect 46284 18398 46286 18450
rect 46338 18398 46340 18450
rect 46284 18386 46340 18398
rect 46396 18562 46564 18564
rect 46396 18510 46510 18562
rect 46562 18510 46564 18562
rect 46396 18508 46564 18510
rect 45164 15262 45166 15314
rect 45218 15262 45220 15314
rect 45164 15250 45220 15262
rect 45388 15260 45892 15316
rect 45948 16828 46116 16884
rect 46172 16996 46228 17006
rect 46172 16882 46228 16940
rect 46172 16830 46174 16882
rect 46226 16830 46228 16882
rect 45388 14530 45444 15260
rect 45948 15204 46004 16828
rect 46172 16818 46228 16830
rect 46172 16100 46228 16110
rect 46172 16006 46228 16044
rect 46284 15988 46340 15998
rect 46284 15894 46340 15932
rect 46060 15876 46116 15886
rect 46116 15820 46228 15876
rect 46060 15810 46116 15820
rect 46060 15316 46116 15326
rect 46060 15222 46116 15260
rect 45836 15148 46004 15204
rect 45500 15090 45556 15102
rect 45500 15038 45502 15090
rect 45554 15038 45556 15090
rect 45500 14644 45556 15038
rect 45500 14578 45556 14588
rect 45388 14478 45390 14530
rect 45442 14478 45444 14530
rect 45388 14466 45444 14478
rect 45276 13860 45332 13870
rect 45276 13300 45332 13804
rect 45612 13524 45668 13534
rect 45276 13244 45444 13300
rect 45164 13076 45220 13086
rect 45164 12850 45220 13020
rect 45164 12798 45166 12850
rect 45218 12798 45220 12850
rect 45164 12786 45220 12798
rect 45276 12962 45332 12974
rect 45276 12910 45278 12962
rect 45330 12910 45332 12962
rect 44380 12290 44436 12302
rect 44380 12238 44382 12290
rect 44434 12238 44436 12290
rect 44380 12068 44436 12238
rect 44716 12292 44772 12302
rect 44716 12198 44772 12236
rect 45052 12178 45108 12348
rect 45052 12126 45054 12178
rect 45106 12126 45108 12178
rect 45052 12114 45108 12126
rect 45164 12516 45220 12526
rect 44380 12002 44436 12012
rect 45164 11620 45220 12460
rect 43932 11218 43988 11228
rect 45052 11564 45220 11620
rect 45276 12180 45332 12910
rect 45052 11060 45108 11564
rect 45164 11284 45220 11294
rect 45276 11284 45332 12124
rect 45388 12292 45444 13244
rect 45388 12178 45444 12236
rect 45388 12126 45390 12178
rect 45442 12126 45444 12178
rect 45388 12114 45444 12126
rect 45500 13074 45556 13086
rect 45500 13022 45502 13074
rect 45554 13022 45556 13074
rect 45388 11956 45444 11966
rect 45388 11394 45444 11900
rect 45388 11342 45390 11394
rect 45442 11342 45444 11394
rect 45388 11330 45444 11342
rect 45220 11228 45332 11284
rect 45164 11190 45220 11228
rect 44132 11004 44396 11014
rect 45052 11004 45332 11060
rect 44188 10948 44236 11004
rect 44292 10948 44340 11004
rect 44132 10938 44396 10948
rect 45164 10836 45220 10846
rect 43596 10546 43652 10556
rect 44268 10834 45220 10836
rect 44268 10782 45166 10834
rect 45218 10782 45220 10834
rect 44268 10780 45220 10782
rect 44268 10610 44324 10780
rect 45164 10770 45220 10780
rect 44268 10558 44270 10610
rect 44322 10558 44324 10610
rect 43484 10108 43652 10164
rect 43596 10052 43652 10108
rect 44268 10052 44324 10558
rect 43596 9996 44100 10052
rect 43596 9940 43652 9996
rect 43596 9874 43652 9884
rect 43484 9828 43540 9838
rect 43932 9828 43988 9838
rect 43484 9714 43540 9772
rect 43820 9772 43932 9828
rect 43484 9662 43486 9714
rect 43538 9662 43540 9714
rect 43484 9650 43540 9662
rect 43708 9716 43764 9726
rect 43260 8642 43316 8652
rect 43372 8818 43428 8830
rect 43372 8766 43374 8818
rect 43426 8766 43428 8818
rect 43036 6750 43038 6802
rect 43090 6750 43092 6802
rect 43036 6738 43092 6750
rect 43260 7586 43316 7598
rect 43260 7534 43262 7586
rect 43314 7534 43316 7586
rect 43260 6692 43316 7534
rect 43372 7364 43428 8766
rect 43708 8146 43764 9660
rect 43820 9268 43876 9772
rect 43932 9762 43988 9772
rect 44044 9828 44100 9996
rect 44268 9986 44324 9996
rect 44604 10610 44660 10622
rect 44604 10558 44606 10610
rect 44658 10558 44660 10610
rect 44044 9826 44548 9828
rect 44044 9774 44046 9826
rect 44098 9774 44548 9826
rect 44044 9772 44548 9774
rect 44044 9762 44100 9772
rect 43932 9602 43988 9614
rect 43932 9550 43934 9602
rect 43986 9550 43988 9602
rect 43932 9492 43988 9550
rect 43932 9426 43988 9436
rect 44132 9436 44396 9446
rect 44188 9380 44236 9436
rect 44292 9380 44340 9436
rect 44132 9370 44396 9380
rect 43932 9268 43988 9278
rect 43820 9266 43988 9268
rect 43820 9214 43934 9266
rect 43986 9214 43988 9266
rect 43820 9212 43988 9214
rect 43932 9202 43988 9212
rect 44492 9266 44548 9772
rect 44492 9214 44494 9266
rect 44546 9214 44548 9266
rect 44492 9202 44548 9214
rect 43932 9044 43988 9054
rect 43932 8818 43988 8988
rect 43932 8766 43934 8818
rect 43986 8766 43988 8818
rect 43932 8754 43988 8766
rect 44044 9042 44100 9054
rect 44044 8990 44046 9042
rect 44098 8990 44100 9042
rect 44044 8484 44100 8990
rect 44044 8418 44100 8428
rect 44604 8484 44660 10558
rect 44716 10612 44772 10622
rect 45052 10612 45108 10622
rect 45276 10612 45332 11004
rect 44716 10518 44772 10556
rect 44828 10610 45332 10612
rect 44828 10558 45054 10610
rect 45106 10558 45332 10610
rect 44828 10556 45332 10558
rect 44716 10164 44772 10174
rect 44716 9268 44772 10108
rect 44828 9826 44884 10556
rect 45052 10546 45108 10556
rect 45164 10388 45220 10398
rect 45164 10386 45332 10388
rect 45164 10334 45166 10386
rect 45218 10334 45332 10386
rect 45164 10332 45332 10334
rect 45164 10322 45220 10332
rect 44828 9774 44830 9826
rect 44882 9774 44884 9826
rect 44828 9762 44884 9774
rect 45052 10052 45108 10062
rect 45276 10052 45332 10332
rect 45276 9996 45444 10052
rect 45052 9826 45108 9996
rect 45052 9774 45054 9826
rect 45106 9774 45108 9826
rect 45052 9762 45108 9774
rect 45164 9938 45220 9950
rect 45164 9886 45166 9938
rect 45218 9886 45220 9938
rect 44940 9268 44996 9278
rect 44716 9266 44996 9268
rect 44716 9214 44942 9266
rect 44994 9214 44996 9266
rect 44716 9212 44996 9214
rect 45164 9268 45220 9886
rect 45276 9828 45332 9838
rect 45276 9714 45332 9772
rect 45276 9662 45278 9714
rect 45330 9662 45332 9714
rect 45276 9650 45332 9662
rect 45388 9716 45444 9996
rect 45388 9650 45444 9660
rect 45276 9268 45332 9278
rect 45164 9266 45332 9268
rect 45164 9214 45278 9266
rect 45330 9214 45332 9266
rect 45164 9212 45332 9214
rect 45500 9268 45556 13022
rect 45612 12402 45668 13468
rect 45612 12350 45614 12402
rect 45666 12350 45668 12402
rect 45612 12292 45668 12350
rect 45836 12404 45892 15148
rect 46172 14532 46228 15820
rect 46396 15764 46452 18508
rect 46508 18498 46564 18508
rect 46844 18450 46900 18462
rect 46844 18398 46846 18450
rect 46898 18398 46900 18450
rect 46844 18228 46900 18398
rect 46844 18162 46900 18172
rect 46956 17668 47012 19070
rect 46620 17612 47012 17668
rect 46508 17554 46564 17566
rect 46508 17502 46510 17554
rect 46562 17502 46564 17554
rect 46508 17108 46564 17502
rect 46508 17042 46564 17052
rect 46508 16660 46564 16670
rect 46508 16098 46564 16604
rect 46508 16046 46510 16098
rect 46562 16046 46564 16098
rect 46508 16034 46564 16046
rect 46284 15708 46452 15764
rect 46284 15148 46340 15708
rect 46396 15540 46452 15550
rect 46396 15314 46452 15484
rect 46396 15262 46398 15314
rect 46450 15262 46452 15314
rect 46396 15250 46452 15262
rect 46620 15428 46676 17612
rect 46844 17444 46900 17454
rect 47068 17444 47124 21308
rect 47516 21298 47572 21308
rect 47628 21252 47684 21308
rect 47628 21186 47684 21196
rect 47180 21140 47236 21150
rect 47180 20802 47236 21084
rect 47180 20750 47182 20802
rect 47234 20750 47236 20802
rect 47180 20738 47236 20750
rect 47852 21028 47908 21420
rect 47852 20802 47908 20972
rect 47852 20750 47854 20802
rect 47906 20750 47908 20802
rect 47852 20738 47908 20750
rect 47964 21420 48076 21476
rect 47628 20692 47684 20702
rect 47628 20598 47684 20636
rect 47404 20578 47460 20590
rect 47404 20526 47406 20578
rect 47458 20526 47460 20578
rect 47404 19908 47460 20526
rect 47852 20132 47908 20142
rect 47852 20038 47908 20076
rect 47404 19842 47460 19852
rect 47180 19572 47236 19582
rect 47180 18562 47236 19516
rect 47404 19348 47460 19358
rect 47292 19124 47348 19134
rect 47292 19030 47348 19068
rect 47404 19122 47460 19292
rect 47852 19236 47908 19246
rect 47852 19142 47908 19180
rect 47404 19070 47406 19122
rect 47458 19070 47460 19122
rect 47404 19058 47460 19070
rect 47964 19122 48020 21420
rect 48076 21410 48132 21420
rect 48188 20468 48244 22764
rect 48524 22594 48580 22988
rect 48860 23044 48916 23054
rect 48860 22950 48916 22988
rect 48972 22820 49028 26126
rect 49084 25732 49140 26350
rect 49308 26292 49364 26572
rect 49308 26226 49364 26236
rect 49140 25676 49252 25732
rect 49084 25666 49140 25676
rect 49084 25506 49140 25518
rect 49084 25454 49086 25506
rect 49138 25454 49140 25506
rect 49084 24612 49140 25454
rect 49196 25284 49252 25676
rect 49532 25618 49588 26908
rect 50540 26964 50596 26974
rect 50540 26870 50596 26908
rect 50652 26908 50708 26918
rect 50652 26906 50820 26908
rect 49868 26852 49924 26862
rect 50652 26854 50654 26906
rect 50706 26854 50820 26906
rect 50652 26852 50820 26854
rect 49868 26850 50260 26852
rect 49868 26798 49870 26850
rect 49922 26798 50260 26850
rect 50652 26842 50708 26852
rect 49868 26796 50260 26798
rect 49868 26786 49924 26796
rect 49532 25566 49534 25618
rect 49586 25566 49588 25618
rect 49532 25554 49588 25566
rect 50204 25956 50260 26796
rect 50764 26786 50820 26796
rect 50428 26292 50484 26302
rect 50428 26198 50484 26236
rect 50092 25396 50148 25406
rect 49196 25218 49252 25228
rect 49532 25394 50148 25396
rect 49532 25342 50094 25394
rect 50146 25342 50148 25394
rect 49532 25340 50148 25342
rect 49420 24836 49476 24846
rect 49420 24722 49476 24780
rect 49420 24670 49422 24722
rect 49474 24670 49476 24722
rect 49420 24658 49476 24670
rect 49084 23938 49140 24556
rect 49308 24610 49364 24622
rect 49308 24558 49310 24610
rect 49362 24558 49364 24610
rect 49308 24164 49364 24558
rect 49308 24098 49364 24108
rect 49084 23886 49086 23938
rect 49138 23886 49140 23938
rect 49084 23874 49140 23886
rect 49420 23940 49476 23950
rect 49532 23940 49588 25340
rect 50092 25330 50148 25340
rect 50204 25284 50260 25900
rect 50204 25282 50372 25284
rect 50204 25230 50206 25282
rect 50258 25230 50372 25282
rect 50204 25228 50372 25230
rect 50204 25218 50260 25228
rect 50316 24500 50372 25228
rect 50428 25282 50484 25294
rect 50428 25230 50430 25282
rect 50482 25230 50484 25282
rect 50428 24948 50484 25230
rect 51100 25284 51156 32396
rect 51436 32386 51492 32396
rect 51548 32340 51604 33516
rect 51660 32676 51716 34076
rect 52892 34130 52948 34142
rect 52892 34078 52894 34130
rect 52946 34078 52948 34130
rect 52892 33236 52948 34078
rect 53340 34132 53396 34142
rect 53340 34038 53396 34076
rect 53228 33572 53284 33582
rect 53116 33460 53172 33470
rect 53116 33366 53172 33404
rect 53228 33346 53284 33516
rect 53228 33294 53230 33346
rect 53282 33294 53284 33346
rect 53228 33282 53284 33294
rect 53564 33348 53620 33358
rect 53788 33348 53844 33358
rect 53564 33346 53844 33348
rect 53564 33294 53566 33346
rect 53618 33294 53790 33346
rect 53842 33294 53844 33346
rect 53564 33292 53844 33294
rect 53564 33282 53620 33292
rect 53788 33282 53844 33292
rect 51772 33124 51828 33134
rect 51772 33030 51828 33068
rect 51996 32676 52052 32686
rect 51660 32674 52052 32676
rect 51660 32622 51998 32674
rect 52050 32622 52052 32674
rect 51660 32620 52052 32622
rect 51548 32284 51716 32340
rect 51286 32172 51550 32182
rect 51342 32116 51390 32172
rect 51446 32116 51494 32172
rect 51286 32106 51550 32116
rect 51660 31948 51716 32284
rect 51324 31892 51716 31948
rect 51996 31948 52052 32620
rect 52892 32562 52948 33180
rect 53004 33122 53060 33134
rect 53004 33070 53006 33122
rect 53058 33070 53060 33122
rect 53004 32900 53060 33070
rect 53004 32844 53284 32900
rect 53228 32786 53284 32844
rect 53228 32734 53230 32786
rect 53282 32734 53284 32786
rect 53228 32722 53284 32734
rect 52892 32510 52894 32562
rect 52946 32510 52948 32562
rect 52892 32498 52948 32510
rect 53116 32564 53172 32574
rect 51996 31892 52276 31948
rect 51324 31890 51380 31892
rect 51324 31838 51326 31890
rect 51378 31838 51380 31890
rect 51324 31826 51380 31838
rect 51996 31778 52052 31790
rect 51996 31726 51998 31778
rect 52050 31726 52052 31778
rect 51996 31668 52052 31726
rect 51884 31612 52052 31668
rect 51772 31554 51828 31566
rect 51772 31502 51774 31554
rect 51826 31502 51828 31554
rect 51660 30994 51716 31006
rect 51660 30942 51662 30994
rect 51714 30942 51716 30994
rect 51286 30604 51550 30614
rect 51342 30548 51390 30604
rect 51446 30548 51494 30604
rect 51286 30538 51550 30548
rect 51548 29538 51604 29550
rect 51548 29486 51550 29538
rect 51602 29486 51604 29538
rect 51212 29316 51268 29326
rect 51548 29316 51604 29486
rect 51660 29540 51716 30942
rect 51772 30882 51828 31502
rect 51772 30830 51774 30882
rect 51826 30830 51828 30882
rect 51772 30818 51828 30830
rect 51660 29474 51716 29484
rect 51772 29986 51828 29998
rect 51772 29934 51774 29986
rect 51826 29934 51828 29986
rect 51772 29428 51828 29934
rect 51772 29362 51828 29372
rect 51548 29260 51716 29316
rect 51212 29222 51268 29260
rect 51660 29204 51716 29260
rect 51884 29204 51940 31612
rect 52220 31556 52276 31892
rect 51660 29148 51940 29204
rect 51996 31500 52276 31556
rect 51286 29036 51550 29046
rect 51342 28980 51390 29036
rect 51446 28980 51494 29036
rect 51286 28970 51550 28980
rect 51548 28868 51604 28878
rect 51436 28644 51492 28654
rect 51436 28550 51492 28588
rect 51436 27860 51492 27870
rect 51436 27766 51492 27804
rect 51548 27746 51604 28812
rect 51660 28084 51716 29148
rect 51884 28756 51940 28766
rect 51884 28642 51940 28700
rect 51884 28590 51886 28642
rect 51938 28590 51940 28642
rect 51884 28196 51940 28590
rect 51996 28308 52052 31500
rect 53004 30994 53060 31006
rect 53004 30942 53006 30994
rect 53058 30942 53060 30994
rect 52668 30210 52724 30222
rect 52668 30158 52670 30210
rect 52722 30158 52724 30210
rect 52668 28868 52724 30158
rect 52780 29988 52836 29998
rect 52780 29894 52836 29932
rect 53004 29988 53060 30942
rect 53004 29922 53060 29932
rect 53004 29428 53060 29438
rect 53004 29334 53060 29372
rect 52668 28802 52724 28812
rect 52780 28756 52836 28766
rect 52780 28662 52836 28700
rect 52108 28532 52164 28542
rect 52108 28438 52164 28476
rect 51996 28252 52276 28308
rect 51884 28140 52052 28196
rect 51772 28084 51828 28094
rect 51660 28028 51772 28084
rect 51772 28018 51828 28028
rect 51548 27694 51550 27746
rect 51602 27694 51604 27746
rect 51548 27682 51604 27694
rect 51884 27972 51940 27982
rect 51286 27468 51550 27478
rect 51342 27412 51390 27468
rect 51446 27412 51494 27468
rect 51286 27402 51550 27412
rect 51884 27300 51940 27916
rect 51884 27234 51940 27244
rect 51548 27074 51604 27086
rect 51548 27022 51550 27074
rect 51602 27022 51604 27074
rect 51548 26852 51604 27022
rect 51884 27074 51940 27086
rect 51884 27022 51886 27074
rect 51938 27022 51940 27074
rect 51884 26964 51940 27022
rect 51884 26898 51940 26908
rect 51548 26180 51604 26796
rect 51660 26628 51716 26638
rect 51660 26402 51716 26572
rect 51884 26628 51940 26638
rect 51996 26628 52052 28140
rect 52220 28082 52276 28252
rect 52220 28030 52222 28082
rect 52274 28030 52276 28082
rect 52220 28018 52276 28030
rect 52556 28196 52612 28206
rect 52444 27970 52500 27982
rect 52444 27918 52446 27970
rect 52498 27918 52500 27970
rect 52108 27748 52164 27758
rect 52108 27186 52164 27692
rect 52444 27636 52500 27918
rect 52444 27570 52500 27580
rect 52556 27970 52612 28140
rect 52556 27918 52558 27970
rect 52610 27918 52612 27970
rect 52108 27134 52110 27186
rect 52162 27134 52164 27186
rect 52108 27122 52164 27134
rect 51940 26572 52052 26628
rect 52556 27076 52612 27918
rect 53004 27860 53060 27870
rect 53004 27766 53060 27804
rect 52892 27748 52948 27758
rect 52892 27654 52948 27692
rect 52780 27300 52836 27310
rect 52780 27206 52836 27244
rect 51884 26562 51940 26572
rect 51660 26350 51662 26402
rect 51714 26350 51716 26402
rect 51660 26338 51716 26350
rect 52556 26402 52612 27020
rect 52892 26962 52948 26974
rect 52892 26910 52894 26962
rect 52946 26910 52948 26962
rect 52556 26350 52558 26402
rect 52610 26350 52612 26402
rect 52556 26338 52612 26350
rect 52780 26850 52836 26862
rect 52780 26798 52782 26850
rect 52834 26798 52836 26850
rect 52108 26180 52164 26190
rect 52220 26180 52276 26190
rect 51548 26124 51716 26180
rect 51286 25900 51550 25910
rect 51342 25844 51390 25900
rect 51446 25844 51494 25900
rect 51286 25834 51550 25844
rect 51212 25732 51268 25742
rect 51212 25506 51268 25676
rect 51212 25454 51214 25506
rect 51266 25454 51268 25506
rect 51212 25442 51268 25454
rect 51548 25620 51604 25630
rect 51548 25506 51604 25564
rect 51660 25618 51716 26124
rect 52108 26178 52220 26180
rect 52108 26126 52110 26178
rect 52162 26126 52220 26178
rect 52108 26124 52220 26126
rect 52108 26114 52164 26124
rect 51660 25566 51662 25618
rect 51714 25566 51716 25618
rect 51660 25554 51716 25566
rect 51772 25732 51828 25742
rect 51548 25454 51550 25506
rect 51602 25454 51604 25506
rect 51548 25442 51604 25454
rect 51100 25228 51492 25284
rect 50428 24882 50484 24892
rect 50540 24836 50596 24846
rect 50596 24780 50708 24836
rect 50540 24742 50596 24780
rect 50428 24724 50484 24734
rect 50428 24630 50484 24668
rect 50316 24444 50596 24500
rect 49756 24276 49812 24286
rect 49756 23940 49812 24220
rect 49420 23938 49588 23940
rect 49420 23886 49422 23938
rect 49474 23886 49588 23938
rect 49420 23884 49588 23886
rect 49644 23938 49812 23940
rect 49644 23886 49758 23938
rect 49810 23886 49812 23938
rect 49644 23884 49812 23886
rect 49308 23714 49364 23726
rect 49308 23662 49310 23714
rect 49362 23662 49364 23714
rect 49308 23380 49364 23662
rect 49308 23314 49364 23324
rect 49084 23268 49140 23278
rect 49084 23154 49140 23212
rect 49084 23102 49086 23154
rect 49138 23102 49140 23154
rect 49084 23090 49140 23102
rect 48972 22754 49028 22764
rect 48524 22542 48526 22594
rect 48578 22542 48580 22594
rect 48524 22530 48580 22542
rect 48412 22484 48468 22494
rect 48412 22260 48468 22428
rect 48972 22372 49028 22382
rect 48524 22260 48580 22270
rect 48412 22258 48580 22260
rect 48412 22206 48526 22258
rect 48578 22206 48580 22258
rect 48412 22204 48580 22206
rect 48300 21588 48356 21598
rect 48300 21494 48356 21532
rect 48412 21364 48468 21374
rect 48188 20412 48356 20468
rect 47964 19070 47966 19122
rect 48018 19070 48020 19122
rect 47964 19058 48020 19070
rect 48076 20020 48132 20030
rect 47180 18510 47182 18562
rect 47234 18510 47236 18562
rect 47180 18452 47236 18510
rect 47628 19010 47684 19022
rect 47628 18958 47630 19010
rect 47682 18958 47684 19010
rect 47180 18386 47236 18396
rect 47516 18450 47572 18462
rect 47516 18398 47518 18450
rect 47570 18398 47572 18450
rect 47516 18004 47572 18398
rect 47516 17938 47572 17948
rect 46844 17442 47124 17444
rect 46844 17390 46846 17442
rect 46898 17390 47124 17442
rect 46844 17388 47124 17390
rect 47516 17442 47572 17454
rect 47516 17390 47518 17442
rect 47570 17390 47572 17442
rect 46732 16996 46788 17006
rect 46732 16660 46788 16940
rect 46844 16884 46900 17388
rect 47516 17220 47572 17390
rect 47404 17164 47572 17220
rect 46956 17108 47012 17118
rect 46956 16994 47012 17052
rect 46956 16942 46958 16994
rect 47010 16942 47012 16994
rect 46956 16930 47012 16942
rect 47292 16996 47348 17006
rect 47292 16902 47348 16940
rect 46844 16818 46900 16828
rect 46956 16772 47012 16782
rect 46732 16604 46900 16660
rect 46620 15314 46676 15372
rect 46620 15262 46622 15314
rect 46674 15262 46676 15314
rect 46620 15250 46676 15262
rect 46732 15986 46788 15998
rect 46732 15934 46734 15986
rect 46786 15934 46788 15986
rect 46732 15316 46788 15934
rect 46844 15986 46900 16604
rect 46844 15934 46846 15986
rect 46898 15934 46900 15986
rect 46844 15922 46900 15934
rect 46956 16436 47012 16716
rect 46956 15540 47012 16380
rect 47068 16212 47124 16222
rect 47068 16098 47124 16156
rect 47404 16100 47460 17164
rect 47628 17108 47684 18958
rect 47852 18900 47908 18910
rect 47852 18674 47908 18844
rect 47852 18622 47854 18674
rect 47906 18622 47908 18674
rect 47852 18610 47908 18622
rect 47964 18788 48020 18798
rect 47964 18452 48020 18732
rect 48076 18564 48132 19964
rect 48188 19236 48244 19246
rect 48188 19142 48244 19180
rect 48188 18788 48244 18798
rect 48300 18788 48356 20412
rect 48244 18732 48356 18788
rect 48188 18722 48244 18732
rect 48188 18564 48244 18574
rect 48076 18508 48188 18564
rect 48244 18508 48356 18564
rect 48188 18498 48244 18508
rect 47852 17556 47908 17566
rect 47852 17462 47908 17500
rect 47964 17332 48020 18396
rect 48300 17444 48356 18508
rect 48412 17668 48468 21308
rect 48524 20914 48580 22204
rect 48636 22260 48692 22270
rect 48972 22260 49028 22316
rect 48636 22258 49028 22260
rect 48636 22206 48638 22258
rect 48690 22206 48974 22258
rect 49026 22206 49028 22258
rect 48636 22204 49028 22206
rect 48636 22194 48692 22204
rect 48524 20862 48526 20914
rect 48578 20862 48580 20914
rect 48524 20850 48580 20862
rect 48860 21474 48916 21486
rect 48860 21422 48862 21474
rect 48914 21422 48916 21474
rect 48860 20804 48916 21422
rect 48972 20916 49028 22204
rect 49308 22260 49364 22270
rect 49420 22260 49476 23884
rect 49364 22204 49476 22260
rect 49644 23268 49700 23884
rect 49756 23874 49812 23884
rect 50428 24052 50484 24062
rect 50428 23938 50484 23996
rect 50428 23886 50430 23938
rect 50482 23886 50484 23938
rect 49868 23716 49924 23726
rect 49868 23622 49924 23660
rect 50092 23716 50148 23726
rect 50092 23622 50148 23660
rect 49756 23604 49812 23614
rect 49756 23380 49812 23548
rect 50204 23380 50260 23390
rect 49756 23324 49924 23380
rect 49308 22166 49364 22204
rect 49644 21364 49700 23212
rect 49756 23044 49812 23054
rect 49756 22950 49812 22988
rect 49868 22370 49924 23324
rect 50204 23286 50260 23324
rect 50428 22708 50484 23886
rect 50540 23940 50596 24444
rect 50652 24164 50708 24780
rect 51436 24834 51492 25228
rect 51436 24782 51438 24834
rect 51490 24782 51492 24834
rect 51436 24770 51492 24782
rect 51548 24948 51604 24958
rect 50764 24724 50820 24734
rect 51324 24724 51380 24734
rect 50764 24722 51380 24724
rect 50764 24670 50766 24722
rect 50818 24670 51326 24722
rect 51378 24670 51380 24722
rect 50764 24668 51380 24670
rect 50764 24658 50820 24668
rect 51100 24164 51156 24668
rect 51324 24658 51380 24668
rect 51548 24724 51604 24892
rect 51548 24722 51716 24724
rect 51548 24670 51550 24722
rect 51602 24670 51716 24722
rect 51548 24668 51716 24670
rect 51548 24658 51604 24668
rect 51286 24332 51550 24342
rect 51342 24276 51390 24332
rect 51446 24276 51494 24332
rect 51286 24266 51550 24276
rect 50652 24108 51044 24164
rect 51100 24108 51380 24164
rect 50540 23884 50932 23940
rect 50540 23716 50596 23726
rect 50540 23622 50596 23660
rect 50764 23716 50820 23726
rect 50764 23622 50820 23660
rect 50652 23268 50708 23278
rect 50652 23174 50708 23212
rect 50484 22652 50596 22708
rect 50428 22642 50484 22652
rect 50428 22372 50484 22382
rect 49868 22318 49870 22370
rect 49922 22318 49924 22370
rect 49868 22306 49924 22318
rect 50092 22370 50484 22372
rect 50092 22318 50430 22370
rect 50482 22318 50484 22370
rect 50092 22316 50484 22318
rect 49980 22146 50036 22158
rect 49980 22094 49982 22146
rect 50034 22094 50036 22146
rect 49756 21700 49812 21710
rect 49980 21700 50036 22094
rect 49812 21644 50036 21700
rect 49756 21586 49812 21644
rect 49756 21534 49758 21586
rect 49810 21534 49812 21586
rect 49756 21522 49812 21534
rect 49644 21308 49924 21364
rect 48972 20850 49028 20860
rect 49308 20804 49364 20814
rect 48636 20748 48916 20804
rect 49084 20802 49364 20804
rect 49084 20750 49310 20802
rect 49362 20750 49364 20802
rect 49084 20748 49364 20750
rect 48636 19124 48692 20748
rect 49084 20692 49140 20748
rect 49308 20738 49364 20748
rect 49644 20802 49700 20814
rect 49644 20750 49646 20802
rect 49698 20750 49700 20802
rect 48748 20636 49140 20692
rect 48748 20018 48804 20636
rect 49196 20578 49252 20590
rect 49196 20526 49198 20578
rect 49250 20526 49252 20578
rect 49196 20468 49252 20526
rect 49196 20402 49252 20412
rect 49420 20578 49476 20590
rect 49420 20526 49422 20578
rect 49474 20526 49476 20578
rect 48748 19966 48750 20018
rect 48802 19966 48804 20018
rect 48748 19684 48804 19966
rect 48748 19618 48804 19628
rect 48860 20356 48916 20366
rect 48860 19460 48916 20300
rect 49420 20244 49476 20526
rect 49420 20178 49476 20188
rect 49532 20578 49588 20590
rect 49532 20526 49534 20578
rect 49586 20526 49588 20578
rect 48636 19058 48692 19068
rect 48748 19404 48916 19460
rect 48972 20020 49028 20030
rect 48972 19460 49028 19964
rect 48748 18788 48804 19404
rect 48972 19394 49028 19404
rect 49084 20018 49140 20030
rect 49084 19966 49086 20018
rect 49138 19966 49140 20018
rect 48860 19236 48916 19246
rect 49084 19236 49140 19966
rect 49532 20018 49588 20526
rect 49644 20132 49700 20750
rect 49644 20066 49700 20076
rect 49532 19966 49534 20018
rect 49586 19966 49588 20018
rect 49532 19572 49588 19966
rect 49756 20020 49812 20030
rect 49756 19926 49812 19964
rect 49868 19796 49924 21308
rect 50092 21252 50148 22316
rect 50428 22260 50484 22316
rect 50428 22194 50484 22204
rect 50204 22148 50260 22158
rect 50204 22054 50260 22092
rect 50092 21186 50148 21196
rect 50316 22036 50372 22046
rect 50316 20802 50372 21980
rect 50316 20750 50318 20802
rect 50370 20750 50372 20802
rect 49532 19506 49588 19516
rect 49644 19740 49924 19796
rect 50204 20468 50260 20478
rect 50204 20018 50260 20412
rect 50316 20356 50372 20750
rect 50428 21586 50484 21598
rect 50428 21534 50430 21586
rect 50482 21534 50484 21586
rect 50428 20804 50484 21534
rect 50540 21476 50596 22652
rect 50652 22370 50708 22382
rect 50652 22318 50654 22370
rect 50706 22318 50708 22370
rect 50652 21924 50708 22318
rect 50876 22148 50932 23884
rect 50988 23378 51044 24108
rect 51324 24050 51380 24108
rect 51324 23998 51326 24050
rect 51378 23998 51380 24050
rect 51324 23986 51380 23998
rect 51660 23938 51716 24668
rect 51660 23886 51662 23938
rect 51714 23886 51716 23938
rect 51660 23874 51716 23886
rect 50988 23326 50990 23378
rect 51042 23326 51044 23378
rect 50988 23314 51044 23326
rect 51324 23828 51380 23838
rect 51324 23604 51380 23772
rect 51324 23154 51380 23548
rect 51548 23716 51604 23726
rect 51548 23266 51604 23660
rect 51548 23214 51550 23266
rect 51602 23214 51604 23266
rect 51548 23202 51604 23214
rect 51324 23102 51326 23154
rect 51378 23102 51380 23154
rect 51324 23090 51380 23102
rect 51286 22764 51550 22774
rect 51342 22708 51390 22764
rect 51446 22708 51494 22764
rect 51286 22698 51550 22708
rect 50988 22372 51044 22382
rect 51548 22372 51604 22382
rect 50988 22370 51604 22372
rect 50988 22318 50990 22370
rect 51042 22318 51550 22370
rect 51602 22318 51604 22370
rect 50988 22316 51604 22318
rect 50988 22306 51044 22316
rect 51548 22306 51604 22316
rect 51772 22260 51828 25676
rect 52108 25284 52164 25294
rect 52108 25190 52164 25228
rect 52220 25060 52276 26124
rect 52780 25732 52836 26798
rect 52780 25666 52836 25676
rect 52892 25620 52948 26910
rect 53116 25620 53172 32508
rect 53340 32004 53396 32042
rect 53340 31938 53396 31948
rect 53900 31948 53956 34748
rect 54236 34738 54292 34748
rect 54572 34356 54628 34862
rect 54236 34300 54628 34356
rect 54236 34130 54292 34300
rect 54236 34078 54238 34130
rect 54290 34078 54292 34130
rect 54236 34066 54292 34078
rect 54460 33572 54516 34300
rect 54684 34242 54740 35084
rect 55132 34692 55188 36204
rect 55916 35924 55972 36428
rect 56028 36260 56084 36270
rect 56028 36166 56084 36204
rect 56028 35924 56084 35934
rect 55916 35922 56084 35924
rect 55916 35870 56030 35922
rect 56082 35870 56084 35922
rect 55916 35868 56084 35870
rect 56028 35858 56084 35868
rect 55580 35812 55636 35822
rect 55580 35718 55636 35756
rect 55244 35700 55300 35710
rect 55244 35606 55300 35644
rect 55692 35588 55748 35598
rect 55356 35476 55412 35486
rect 55356 34916 55412 35420
rect 55356 34850 55412 34860
rect 55468 34914 55524 34926
rect 55468 34862 55470 34914
rect 55522 34862 55524 34914
rect 55132 34354 55188 34636
rect 55132 34302 55134 34354
rect 55186 34302 55188 34354
rect 55132 34290 55188 34302
rect 54684 34190 54686 34242
rect 54738 34190 54740 34242
rect 54684 34178 54740 34190
rect 54572 34132 54628 34142
rect 54572 34038 54628 34076
rect 55468 34132 55524 34862
rect 55468 34066 55524 34076
rect 55692 34916 55748 35532
rect 54460 33478 54516 33516
rect 55692 33460 55748 34860
rect 56140 35252 56196 35262
rect 56140 34802 56196 35196
rect 56252 35028 56308 37212
rect 56364 37156 56420 37166
rect 56364 35476 56420 37100
rect 56476 36372 56532 36382
rect 56476 36278 56532 36316
rect 56700 36036 56756 39200
rect 56924 36596 56980 36606
rect 56924 36502 56980 36540
rect 56588 35980 56756 36036
rect 58439 36092 58703 36102
rect 58495 36036 58543 36092
rect 58599 36036 58647 36092
rect 58439 36026 58703 36036
rect 56476 35700 56532 35710
rect 56476 35606 56532 35644
rect 56364 35420 56532 35476
rect 56252 34962 56308 34972
rect 56140 34750 56142 34802
rect 56194 34750 56196 34802
rect 56140 34356 56196 34750
rect 56140 34300 56308 34356
rect 55916 34132 55972 34142
rect 55804 33460 55860 33470
rect 55692 33458 55860 33460
rect 55692 33406 55806 33458
rect 55858 33406 55860 33458
rect 55692 33404 55860 33406
rect 55804 33394 55860 33404
rect 54124 33236 54180 33246
rect 54572 33236 54628 33246
rect 54124 33234 54404 33236
rect 54124 33182 54126 33234
rect 54178 33182 54404 33234
rect 54124 33180 54404 33182
rect 54124 33170 54180 33180
rect 54012 33122 54068 33134
rect 54012 33070 54014 33122
rect 54066 33070 54068 33122
rect 54012 33012 54068 33070
rect 54012 32956 54180 33012
rect 54124 32564 54180 32956
rect 54236 32564 54292 32574
rect 54124 32508 54236 32564
rect 54236 32470 54292 32508
rect 54012 32450 54068 32462
rect 54012 32398 54014 32450
rect 54066 32398 54068 32450
rect 54012 32340 54068 32398
rect 54348 32340 54404 33180
rect 54572 33234 54964 33236
rect 54572 33182 54574 33234
rect 54626 33182 54964 33234
rect 54572 33180 54964 33182
rect 54572 33170 54628 33180
rect 54908 32674 54964 33180
rect 55916 32900 55972 34076
rect 54908 32622 54910 32674
rect 54962 32622 54964 32674
rect 54908 32610 54964 32622
rect 55804 32844 55972 32900
rect 56028 33346 56084 33358
rect 56028 33294 56030 33346
rect 56082 33294 56084 33346
rect 55804 32674 55860 32844
rect 56028 32788 56084 33294
rect 56140 32788 56196 32798
rect 56028 32786 56196 32788
rect 56028 32734 56142 32786
rect 56194 32734 56196 32786
rect 56028 32732 56196 32734
rect 56140 32722 56196 32732
rect 55804 32622 55806 32674
rect 55858 32622 55860 32674
rect 54068 32284 54404 32340
rect 55132 32452 55188 32462
rect 54012 32274 54068 32284
rect 53676 31890 53732 31902
rect 53900 31892 54068 31948
rect 53676 31838 53678 31890
rect 53730 31838 53732 31890
rect 53564 31780 53620 31790
rect 53564 31686 53620 31724
rect 53676 30436 53732 31838
rect 53676 30370 53732 30380
rect 53788 30994 53844 31006
rect 53788 30942 53790 30994
rect 53842 30942 53844 30994
rect 53228 30210 53284 30222
rect 53228 30158 53230 30210
rect 53282 30158 53284 30210
rect 53228 29428 53284 30158
rect 53788 30212 53844 30942
rect 53228 29362 53284 29372
rect 53340 30098 53396 30110
rect 53340 30046 53342 30098
rect 53394 30046 53396 30098
rect 53340 29316 53396 30046
rect 53788 29538 53844 30156
rect 53788 29486 53790 29538
rect 53842 29486 53844 29538
rect 53788 29474 53844 29486
rect 53340 29250 53396 29260
rect 54012 29204 54068 31892
rect 54908 31892 54964 31902
rect 54684 31778 54740 31790
rect 54684 31726 54686 31778
rect 54738 31726 54740 31778
rect 54236 30884 54292 30894
rect 54460 30884 54516 30894
rect 54236 30882 54460 30884
rect 54236 30830 54238 30882
rect 54290 30830 54460 30882
rect 54236 30828 54460 30830
rect 54236 30818 54292 30828
rect 54460 30818 54516 30828
rect 54460 30324 54516 30334
rect 54460 30230 54516 30268
rect 54012 29138 54068 29148
rect 54124 30100 54180 30110
rect 53788 29092 53844 29102
rect 53228 28644 53284 28654
rect 53228 28550 53284 28588
rect 53788 28644 53844 29036
rect 54124 28868 54180 30044
rect 54236 29988 54292 29998
rect 54348 29988 54404 29998
rect 54292 29986 54404 29988
rect 54292 29934 54350 29986
rect 54402 29934 54404 29986
rect 54292 29932 54404 29934
rect 54236 29092 54292 29932
rect 54348 29922 54404 29932
rect 54348 29540 54404 29550
rect 54348 29446 54404 29484
rect 54572 29428 54628 29438
rect 54572 29334 54628 29372
rect 54236 29026 54292 29036
rect 54012 28812 54180 28868
rect 54684 28868 54740 31726
rect 54908 31778 54964 31836
rect 54908 31726 54910 31778
rect 54962 31726 54964 31778
rect 54908 31714 54964 31726
rect 55132 31778 55188 32396
rect 55468 32450 55524 32462
rect 55468 32398 55470 32450
rect 55522 32398 55524 32450
rect 55468 31892 55524 32398
rect 55804 32002 55860 32622
rect 55916 32676 55972 32686
rect 55916 32582 55972 32620
rect 55804 31950 55806 32002
rect 55858 31950 55860 32002
rect 55804 31938 55860 31950
rect 56252 31948 56308 34300
rect 56476 32676 56532 35420
rect 56588 35140 56644 35980
rect 56700 35868 56980 35924
rect 56700 35810 56756 35868
rect 56700 35758 56702 35810
rect 56754 35758 56756 35810
rect 56700 35746 56756 35758
rect 56812 35698 56868 35710
rect 56812 35646 56814 35698
rect 56866 35646 56868 35698
rect 56588 35074 56644 35084
rect 56700 35252 56756 35262
rect 56812 35252 56868 35646
rect 56756 35196 56868 35252
rect 56700 35026 56756 35196
rect 56700 34974 56702 35026
rect 56754 34974 56756 35026
rect 56700 34962 56756 34974
rect 56924 35028 56980 35868
rect 58156 35028 58212 35038
rect 56924 34972 57204 35028
rect 57148 34914 57204 34972
rect 57148 34862 57150 34914
rect 57202 34862 57204 34914
rect 56588 34804 56644 34814
rect 56588 34242 56644 34748
rect 57148 34692 57204 34862
rect 56588 34190 56590 34242
rect 56642 34190 56644 34242
rect 56588 34178 56644 34190
rect 57036 34636 57204 34692
rect 57260 35026 58324 35028
rect 57260 34974 58158 35026
rect 58210 34974 58324 35026
rect 57260 34972 58324 34974
rect 56700 34132 56756 34142
rect 56700 34038 56756 34076
rect 56588 32676 56644 32686
rect 56476 32674 56644 32676
rect 56476 32622 56590 32674
rect 56642 32622 56644 32674
rect 56476 32620 56644 32622
rect 56588 32610 56644 32620
rect 55468 31826 55524 31836
rect 56028 31892 56308 31948
rect 57036 31948 57092 34636
rect 57260 34130 57316 34972
rect 58156 34962 58212 34972
rect 57260 34078 57262 34130
rect 57314 34078 57316 34130
rect 57260 34066 57316 34078
rect 57596 34802 57652 34814
rect 57596 34750 57598 34802
rect 57650 34750 57652 34802
rect 57596 33458 57652 34750
rect 58156 34020 58212 34030
rect 57596 33406 57598 33458
rect 57650 33406 57652 33458
rect 57596 33394 57652 33406
rect 58044 34018 58212 34020
rect 58044 33966 58158 34018
rect 58210 33966 58212 34018
rect 58044 33964 58212 33966
rect 57932 33348 57988 33358
rect 58044 33348 58100 33964
rect 58156 33954 58212 33964
rect 57932 33346 58100 33348
rect 57932 33294 57934 33346
rect 57986 33294 58100 33346
rect 57932 33292 58100 33294
rect 57932 33282 57988 33292
rect 57484 32562 57540 32574
rect 57484 32510 57486 32562
rect 57538 32510 57540 32562
rect 57148 32452 57204 32462
rect 57148 32358 57204 32396
rect 57036 31892 57316 31948
rect 55132 31726 55134 31778
rect 55186 31726 55188 31778
rect 55132 31332 55188 31726
rect 56028 31778 56084 31892
rect 56028 31726 56030 31778
rect 56082 31726 56084 31778
rect 56028 31714 56084 31726
rect 56588 31780 56644 31790
rect 55132 31276 55412 31332
rect 55244 31106 55300 31118
rect 55244 31054 55246 31106
rect 55298 31054 55300 31106
rect 55244 30884 55300 31054
rect 55244 30818 55300 30828
rect 55356 30434 55412 31276
rect 56588 31106 56644 31724
rect 56924 31780 56980 31790
rect 56924 31686 56980 31724
rect 57260 31778 57316 31892
rect 57260 31726 57262 31778
rect 57314 31726 57316 31778
rect 56588 31054 56590 31106
rect 56642 31054 56644 31106
rect 56588 31042 56644 31054
rect 55356 30382 55358 30434
rect 55410 30382 55412 30434
rect 55356 30370 55412 30382
rect 55468 30994 55524 31006
rect 55468 30942 55470 30994
rect 55522 30942 55524 30994
rect 55468 30100 55524 30942
rect 57036 30994 57092 31006
rect 57036 30942 57038 30994
rect 57090 30942 57092 30994
rect 56140 30882 56196 30894
rect 56140 30830 56142 30882
rect 56194 30830 56196 30882
rect 55692 30212 55748 30222
rect 55692 30118 55748 30156
rect 55468 30034 55524 30044
rect 55804 30100 55860 30110
rect 55804 29538 55860 30044
rect 56140 29652 56196 30830
rect 56700 30324 56756 30334
rect 57036 30324 57092 30942
rect 56756 30268 57092 30324
rect 57148 30324 57204 30334
rect 56700 30210 56756 30268
rect 56700 30158 56702 30210
rect 56754 30158 56756 30210
rect 56700 30146 56756 30158
rect 56140 29586 56196 29596
rect 56924 29652 56980 29662
rect 55804 29486 55806 29538
rect 55858 29486 55860 29538
rect 54796 29426 54852 29438
rect 54796 29374 54798 29426
rect 54850 29374 54852 29426
rect 54796 29316 54852 29374
rect 54796 29250 54852 29260
rect 54012 28756 54068 28812
rect 54684 28802 54740 28812
rect 55692 28868 55748 28878
rect 55692 28774 55748 28812
rect 54012 28690 54068 28700
rect 54124 28700 54628 28756
rect 53788 27748 53844 28588
rect 54124 27970 54180 28700
rect 54572 28642 54628 28700
rect 54572 28590 54574 28642
rect 54626 28590 54628 28642
rect 54348 28532 54404 28542
rect 54236 28084 54292 28094
rect 54236 27990 54292 28028
rect 54124 27918 54126 27970
rect 54178 27918 54180 27970
rect 54124 27906 54180 27918
rect 54348 27858 54404 28476
rect 54572 28084 54628 28590
rect 55020 28644 55076 28654
rect 55020 28550 55076 28588
rect 55804 28644 55860 29486
rect 55916 29540 55972 29550
rect 55916 29446 55972 29484
rect 56924 29538 56980 29596
rect 56924 29486 56926 29538
rect 56978 29486 56980 29538
rect 56140 29428 56196 29438
rect 56588 29428 56644 29438
rect 56140 29426 56644 29428
rect 56140 29374 56142 29426
rect 56194 29374 56590 29426
rect 56642 29374 56644 29426
rect 56140 29372 56644 29374
rect 56140 29362 56196 29372
rect 56588 29362 56644 29372
rect 55804 28578 55860 28588
rect 55916 29204 55972 29214
rect 54572 28028 55076 28084
rect 55020 27970 55076 28028
rect 55020 27918 55022 27970
rect 55074 27918 55076 27970
rect 55020 27906 55076 27918
rect 54348 27806 54350 27858
rect 54402 27806 54404 27858
rect 54348 27794 54404 27806
rect 54684 27858 54740 27870
rect 54684 27806 54686 27858
rect 54738 27806 54740 27858
rect 53788 27682 53844 27692
rect 53900 27746 53956 27758
rect 53900 27694 53902 27746
rect 53954 27694 53956 27746
rect 53900 27524 53956 27694
rect 54572 27748 54628 27758
rect 53900 27468 54068 27524
rect 53340 26962 53396 26974
rect 53340 26910 53342 26962
rect 53394 26910 53396 26962
rect 53340 26404 53396 26910
rect 53452 26964 53508 26974
rect 53452 26962 53620 26964
rect 53452 26910 53454 26962
rect 53506 26910 53620 26962
rect 53452 26908 53620 26910
rect 53452 26898 53508 26908
rect 53340 26338 53396 26348
rect 53452 26628 53508 26638
rect 53228 26290 53284 26302
rect 53228 26238 53230 26290
rect 53282 26238 53284 26290
rect 53228 26180 53284 26238
rect 53452 26290 53508 26572
rect 53452 26238 53454 26290
rect 53506 26238 53508 26290
rect 53452 26180 53508 26238
rect 53228 26114 53284 26124
rect 53340 26124 53508 26180
rect 53228 25620 53284 25630
rect 53116 25618 53284 25620
rect 53116 25566 53230 25618
rect 53282 25566 53284 25618
rect 53116 25564 53284 25566
rect 52892 25554 52948 25564
rect 53228 25554 53284 25564
rect 53340 25508 53396 26124
rect 53340 25442 53396 25452
rect 53452 25396 53508 25406
rect 53564 25396 53620 26908
rect 53676 26850 53732 26862
rect 53676 26798 53678 26850
rect 53730 26798 53732 26850
rect 53676 25506 53732 26798
rect 53676 25454 53678 25506
rect 53730 25454 53732 25506
rect 53676 25442 53732 25454
rect 53900 26852 53956 26862
rect 53508 25340 53620 25396
rect 52108 25004 52276 25060
rect 53116 25282 53172 25294
rect 53116 25230 53118 25282
rect 53170 25230 53172 25282
rect 51996 24164 52052 24174
rect 51996 24070 52052 24108
rect 51884 22930 51940 22942
rect 51884 22878 51886 22930
rect 51938 22878 51940 22930
rect 51884 22370 51940 22878
rect 51884 22318 51886 22370
rect 51938 22318 51940 22370
rect 51884 22306 51940 22318
rect 51660 22204 51828 22260
rect 51996 22260 52052 22270
rect 51324 22148 51380 22158
rect 50876 22092 51268 22148
rect 50876 21924 50932 21934
rect 50652 21868 50876 21924
rect 50876 21858 50932 21868
rect 50988 21812 51044 21822
rect 50652 21700 50708 21710
rect 50652 21588 50708 21644
rect 50988 21698 51044 21756
rect 50988 21646 50990 21698
rect 51042 21646 51044 21698
rect 50988 21634 51044 21646
rect 51100 21698 51156 21710
rect 51100 21646 51102 21698
rect 51154 21646 51156 21698
rect 51100 21588 51156 21646
rect 50652 21532 50932 21588
rect 50876 21476 50932 21532
rect 51100 21522 51156 21532
rect 50540 21420 50820 21476
rect 50876 21420 51044 21476
rect 50652 21252 50708 21262
rect 50428 20578 50484 20748
rect 50428 20526 50430 20578
rect 50482 20526 50484 20578
rect 50428 20468 50484 20526
rect 50428 20402 50484 20412
rect 50540 21196 50652 21252
rect 50316 20290 50372 20300
rect 50540 20188 50596 21196
rect 50652 21186 50708 21196
rect 50652 20804 50708 20814
rect 50764 20804 50820 21420
rect 50876 20916 50932 20926
rect 50876 20804 50932 20860
rect 50764 20802 50932 20804
rect 50764 20750 50878 20802
rect 50930 20750 50932 20802
rect 50764 20748 50932 20750
rect 50652 20710 50708 20748
rect 50876 20738 50932 20748
rect 50988 20690 51044 21420
rect 51212 21364 51268 22092
rect 51324 22054 51380 22092
rect 51436 22148 51492 22158
rect 51660 22148 51716 22204
rect 51436 22146 51716 22148
rect 51436 22094 51438 22146
rect 51490 22094 51716 22146
rect 51436 22092 51716 22094
rect 51436 22082 51492 22092
rect 51324 21924 51380 21934
rect 51324 21810 51380 21868
rect 51324 21758 51326 21810
rect 51378 21758 51380 21810
rect 51324 21746 51380 21758
rect 51996 21698 52052 22204
rect 51996 21646 51998 21698
rect 52050 21646 52052 21698
rect 51996 21634 52052 21646
rect 50988 20638 50990 20690
rect 51042 20638 51044 20690
rect 50988 20626 51044 20638
rect 51100 21308 51268 21364
rect 50316 20132 50596 20188
rect 50876 20468 50932 20478
rect 50876 20242 50932 20412
rect 50876 20190 50878 20242
rect 50930 20190 50932 20242
rect 50876 20178 50932 20190
rect 50316 20038 50372 20076
rect 50204 19966 50206 20018
rect 50258 19966 50260 20018
rect 48860 19234 49140 19236
rect 48860 19182 48862 19234
rect 48914 19182 49140 19234
rect 48860 19180 49140 19182
rect 49532 19234 49588 19246
rect 49532 19182 49534 19234
rect 49586 19182 49588 19234
rect 48860 19012 48916 19180
rect 49420 19124 49476 19134
rect 48860 18946 48916 18956
rect 49084 19010 49140 19022
rect 49084 18958 49086 19010
rect 49138 18958 49140 19010
rect 49084 18900 49140 18958
rect 48748 18732 49028 18788
rect 48412 17612 48580 17668
rect 48412 17444 48468 17454
rect 48300 17442 48468 17444
rect 48300 17390 48414 17442
rect 48466 17390 48468 17442
rect 48300 17388 48468 17390
rect 48412 17378 48468 17388
rect 47964 17266 48020 17276
rect 47516 17052 47684 17108
rect 47740 17220 47796 17230
rect 47740 17106 47796 17164
rect 47740 17054 47742 17106
rect 47794 17054 47796 17106
rect 47516 16772 47572 17052
rect 47740 17042 47796 17054
rect 47852 16996 47908 17006
rect 47628 16884 47684 16894
rect 47628 16790 47684 16828
rect 47516 16706 47572 16716
rect 47068 16046 47070 16098
rect 47122 16046 47124 16098
rect 47068 16034 47124 16046
rect 47292 16044 47460 16100
rect 47740 16658 47796 16670
rect 47740 16606 47742 16658
rect 47794 16606 47796 16658
rect 46956 15474 47012 15484
rect 47292 15540 47348 16044
rect 47404 15876 47460 15886
rect 47516 15876 47572 15886
rect 47404 15874 47516 15876
rect 47404 15822 47406 15874
rect 47458 15822 47516 15874
rect 47404 15820 47516 15822
rect 47404 15810 47460 15820
rect 47404 15540 47460 15550
rect 47292 15538 47460 15540
rect 47292 15486 47406 15538
rect 47458 15486 47460 15538
rect 47292 15484 47460 15486
rect 46732 15250 46788 15260
rect 47292 15316 47348 15484
rect 47404 15474 47460 15484
rect 47292 15250 47348 15260
rect 46284 15092 46900 15148
rect 46172 14438 46228 14476
rect 46620 14644 46676 14654
rect 46284 14420 46340 14430
rect 46284 14418 46452 14420
rect 46284 14366 46286 14418
rect 46338 14366 46452 14418
rect 46284 14364 46452 14366
rect 46284 14354 46340 14364
rect 46284 13858 46340 13870
rect 46284 13806 46286 13858
rect 46338 13806 46340 13858
rect 46060 13634 46116 13646
rect 46060 13582 46062 13634
rect 46114 13582 46116 13634
rect 46060 12964 46116 13582
rect 46060 12898 46116 12908
rect 46284 13412 46340 13806
rect 46284 12962 46340 13356
rect 46284 12910 46286 12962
rect 46338 12910 46340 12962
rect 46284 12898 46340 12910
rect 46396 12964 46452 14364
rect 46396 12898 46452 12908
rect 46172 12852 46228 12862
rect 46172 12738 46228 12796
rect 46172 12686 46174 12738
rect 46226 12686 46228 12738
rect 46172 12674 46228 12686
rect 45836 12348 46004 12404
rect 45612 11956 45668 12236
rect 45836 12180 45892 12190
rect 45836 12086 45892 12124
rect 45724 12066 45780 12078
rect 45724 12014 45726 12066
rect 45778 12014 45780 12066
rect 45724 11956 45780 12014
rect 45836 11956 45892 11966
rect 45724 11900 45836 11956
rect 45612 11890 45668 11900
rect 45836 11890 45892 11900
rect 45948 11788 46004 12348
rect 46172 12178 46228 12190
rect 46172 12126 46174 12178
rect 46226 12126 46228 12178
rect 46172 12068 46228 12126
rect 46396 12180 46452 12218
rect 46396 12114 46452 12124
rect 46620 12178 46676 14588
rect 46844 14530 46900 15092
rect 46956 15092 47012 15102
rect 46956 14998 47012 15036
rect 46844 14478 46846 14530
rect 46898 14478 46900 14530
rect 46844 14466 46900 14478
rect 46956 14644 47012 14654
rect 46956 14532 47012 14588
rect 47292 14532 47348 14542
rect 46956 14530 47348 14532
rect 46956 14478 47294 14530
rect 47346 14478 47348 14530
rect 46956 14476 47348 14478
rect 47292 14466 47348 14476
rect 47404 14306 47460 14318
rect 47404 14254 47406 14306
rect 47458 14254 47460 14306
rect 47292 13860 47348 13870
rect 47292 13766 47348 13804
rect 46844 12964 46900 12974
rect 46900 12908 47012 12964
rect 46844 12870 46900 12908
rect 46620 12126 46622 12178
rect 46674 12126 46676 12178
rect 46620 12114 46676 12126
rect 46844 12292 46900 12302
rect 46172 12002 46228 12012
rect 46284 12066 46340 12078
rect 46284 12014 46286 12066
rect 46338 12014 46340 12066
rect 45724 11732 45780 11742
rect 45724 11618 45780 11676
rect 45724 11566 45726 11618
rect 45778 11566 45780 11618
rect 45724 11554 45780 11566
rect 45836 11732 46004 11788
rect 46060 11844 46116 11854
rect 45724 11394 45780 11406
rect 45724 11342 45726 11394
rect 45778 11342 45780 11394
rect 45724 11284 45780 11342
rect 45612 9716 45668 9726
rect 45612 9622 45668 9660
rect 45724 9714 45780 11228
rect 45836 10052 45892 11732
rect 45948 11396 46004 11406
rect 45948 11170 46004 11340
rect 45948 11118 45950 11170
rect 46002 11118 46004 11170
rect 45948 10610 46004 11118
rect 45948 10558 45950 10610
rect 46002 10558 46004 10610
rect 45948 10546 46004 10558
rect 45948 10052 46004 10062
rect 45836 9996 45948 10052
rect 45948 9986 46004 9996
rect 45948 9828 46004 9838
rect 45948 9734 46004 9772
rect 45724 9662 45726 9714
rect 45778 9662 45780 9714
rect 45724 9650 45780 9662
rect 46060 9268 46116 11788
rect 46284 11732 46340 12014
rect 46508 11956 46564 11966
rect 46508 11788 46564 11900
rect 46172 11676 46284 11732
rect 46172 10610 46228 11676
rect 46284 11666 46340 11676
rect 46396 11732 46564 11788
rect 46620 11844 46676 11854
rect 46396 11284 46452 11732
rect 46620 11508 46676 11788
rect 46732 11508 46788 11518
rect 46620 11506 46788 11508
rect 46620 11454 46734 11506
rect 46786 11454 46788 11506
rect 46620 11452 46788 11454
rect 46732 11442 46788 11452
rect 46396 10722 46452 11228
rect 46844 10724 46900 12236
rect 46956 11508 47012 12908
rect 47180 12404 47236 12414
rect 47180 12310 47236 12348
rect 47292 12180 47348 12190
rect 47068 12178 47348 12180
rect 47068 12126 47294 12178
rect 47346 12126 47348 12178
rect 47068 12124 47348 12126
rect 47068 12068 47124 12124
rect 47292 12114 47348 12124
rect 47068 12002 47124 12012
rect 47404 12068 47460 14254
rect 47516 13636 47572 15820
rect 47740 14532 47796 16606
rect 47852 16098 47908 16940
rect 48412 16212 48468 16222
rect 48412 16118 48468 16156
rect 47852 16046 47854 16098
rect 47906 16046 47908 16098
rect 47852 16034 47908 16046
rect 48188 16100 48244 16110
rect 48188 16006 48244 16044
rect 47964 15988 48020 15998
rect 48020 15932 48132 15988
rect 47964 15894 48020 15932
rect 48076 15538 48132 15932
rect 48076 15486 48078 15538
rect 48130 15486 48132 15538
rect 48076 15474 48132 15486
rect 48188 15428 48244 15438
rect 48188 15334 48244 15372
rect 48524 15148 48580 17612
rect 48748 17666 48804 18732
rect 48972 18450 49028 18732
rect 48972 18398 48974 18450
rect 49026 18398 49028 18450
rect 48972 18386 49028 18398
rect 49084 18228 49140 18844
rect 48748 17614 48750 17666
rect 48802 17614 48804 17666
rect 48748 17556 48804 17614
rect 48748 17490 48804 17500
rect 48972 18172 49140 18228
rect 49308 18228 49364 18238
rect 48860 17442 48916 17454
rect 48860 17390 48862 17442
rect 48914 17390 48916 17442
rect 48748 16772 48804 16782
rect 48636 16100 48692 16110
rect 48636 16006 48692 16044
rect 48076 15092 48132 15102
rect 48412 15092 48580 15148
rect 48636 15092 48692 15102
rect 48076 15090 48356 15092
rect 48076 15038 48078 15090
rect 48130 15038 48356 15090
rect 48076 15036 48356 15038
rect 48076 15026 48132 15036
rect 48076 14532 48132 14542
rect 47740 14476 48076 14532
rect 48076 14418 48132 14476
rect 48076 14366 48078 14418
rect 48130 14366 48132 14418
rect 47516 13570 47572 13580
rect 47852 13746 47908 13758
rect 47852 13694 47854 13746
rect 47906 13694 47908 13746
rect 47852 13300 47908 13694
rect 47852 13234 47908 13244
rect 47516 12964 47572 12974
rect 48076 12964 48132 14366
rect 48300 14420 48356 15036
rect 48300 14326 48356 14364
rect 48188 14308 48244 14318
rect 48188 14214 48244 14252
rect 48300 13636 48356 13646
rect 47516 12962 48132 12964
rect 47516 12910 47518 12962
rect 47570 12910 48132 12962
rect 47516 12908 48132 12910
rect 48188 13412 48244 13422
rect 47516 12898 47572 12908
rect 47852 12404 47908 12414
rect 48188 12404 48244 13356
rect 47852 12402 48244 12404
rect 47852 12350 47854 12402
rect 47906 12350 48244 12402
rect 47852 12348 48244 12350
rect 48300 13076 48356 13580
rect 48300 12402 48356 13020
rect 48300 12350 48302 12402
rect 48354 12350 48356 12402
rect 47852 12338 47908 12348
rect 48300 12338 48356 12350
rect 47404 12002 47460 12012
rect 47180 11956 47236 11966
rect 47180 11862 47236 11900
rect 46956 11396 47012 11452
rect 47964 11508 48020 11518
rect 47964 11414 48020 11452
rect 47068 11396 47124 11406
rect 46956 11394 47124 11396
rect 46956 11342 47070 11394
rect 47122 11342 47124 11394
rect 46956 11340 47124 11342
rect 47068 11330 47124 11340
rect 48188 11396 48244 11406
rect 48188 11302 48244 11340
rect 47628 11284 47684 11294
rect 46396 10670 46398 10722
rect 46450 10670 46452 10722
rect 46396 10658 46452 10670
rect 46508 10668 46900 10724
rect 47516 11282 47684 11284
rect 47516 11230 47630 11282
rect 47682 11230 47684 11282
rect 47516 11228 47684 11230
rect 46172 10558 46174 10610
rect 46226 10558 46228 10610
rect 46172 10546 46228 10558
rect 45500 9212 45668 9268
rect 44940 9202 44996 9212
rect 45276 9202 45332 9212
rect 45500 9044 45556 9054
rect 45388 8932 45444 8970
rect 45500 8950 45556 8988
rect 45388 8866 45444 8876
rect 44604 8418 44660 8428
rect 45388 8708 45444 8718
rect 45388 8370 45444 8652
rect 45388 8318 45390 8370
rect 45442 8318 45444 8370
rect 45388 8306 45444 8318
rect 45612 8372 45668 9212
rect 46060 9202 46116 9212
rect 46284 10498 46340 10510
rect 46284 10446 46286 10498
rect 46338 10446 46340 10498
rect 46284 9266 46340 10446
rect 46508 10164 46564 10668
rect 47068 10610 47124 10622
rect 47068 10558 47070 10610
rect 47122 10558 47124 10610
rect 46844 10498 46900 10510
rect 46844 10446 46846 10498
rect 46898 10446 46900 10498
rect 46284 9214 46286 9266
rect 46338 9214 46340 9266
rect 46284 9202 46340 9214
rect 46396 10108 46564 10164
rect 46732 10386 46788 10398
rect 46732 10334 46734 10386
rect 46786 10334 46788 10386
rect 45948 9044 46004 9054
rect 45948 9042 46228 9044
rect 45948 8990 45950 9042
rect 46002 8990 46228 9042
rect 45948 8988 46228 8990
rect 45948 8978 46004 8988
rect 46172 8596 46228 8988
rect 46284 8930 46340 8942
rect 46284 8878 46286 8930
rect 46338 8878 46340 8930
rect 46284 8820 46340 8878
rect 46284 8754 46340 8764
rect 46396 8708 46452 10108
rect 46620 10052 46676 10062
rect 46508 9996 46620 10052
rect 46508 9714 46564 9996
rect 46620 9986 46676 9996
rect 46620 9828 46676 9838
rect 46732 9828 46788 10334
rect 46676 9772 46788 9828
rect 46620 9734 46676 9772
rect 46508 9662 46510 9714
rect 46562 9662 46564 9714
rect 46508 9650 46564 9662
rect 46844 9380 46900 10446
rect 47068 10164 47124 10558
rect 46956 10108 47236 10164
rect 46956 10052 47012 10108
rect 46956 9986 47012 9996
rect 47068 9938 47124 9950
rect 47068 9886 47070 9938
rect 47122 9886 47124 9938
rect 46956 9714 47012 9726
rect 46956 9662 46958 9714
rect 47010 9662 47012 9714
rect 46956 9604 47012 9662
rect 46956 9538 47012 9548
rect 46508 9324 46900 9380
rect 46508 9154 46564 9324
rect 46508 9102 46510 9154
rect 46562 9102 46564 9154
rect 46508 9090 46564 9102
rect 47068 8820 47124 9886
rect 47068 8754 47124 8764
rect 46396 8652 46900 8708
rect 46172 8540 46564 8596
rect 45612 8306 45668 8316
rect 46396 8372 46452 8382
rect 45724 8258 45780 8270
rect 45724 8206 45726 8258
rect 45778 8206 45780 8258
rect 43708 8094 43710 8146
rect 43762 8094 43764 8146
rect 43708 8036 43764 8094
rect 43932 8148 43988 8158
rect 43932 8054 43988 8092
rect 44828 8146 44884 8158
rect 44828 8094 44830 8146
rect 44882 8094 44884 8146
rect 43708 7970 43764 7980
rect 44716 8036 44772 8046
rect 44132 7868 44396 7878
rect 44188 7812 44236 7868
rect 44292 7812 44340 7868
rect 44132 7802 44396 7812
rect 43484 7476 43540 7486
rect 43820 7476 43876 7486
rect 43484 7382 43540 7420
rect 43596 7474 43876 7476
rect 43596 7422 43822 7474
rect 43874 7422 43876 7474
rect 43596 7420 43876 7422
rect 43372 7298 43428 7308
rect 43260 6626 43316 6636
rect 43596 6690 43652 7420
rect 43820 7410 43876 7420
rect 44604 7476 44660 7486
rect 44716 7476 44772 7980
rect 44828 7924 44884 8094
rect 44940 8036 44996 8046
rect 44940 7942 44996 7980
rect 44828 7858 44884 7868
rect 44828 7700 44884 7710
rect 44828 7606 44884 7644
rect 44940 7476 44996 7486
rect 44716 7474 44996 7476
rect 44716 7422 44942 7474
rect 44994 7422 44996 7474
rect 44716 7420 44996 7422
rect 44604 7382 44660 7420
rect 44940 7410 44996 7420
rect 45724 7476 45780 8206
rect 46060 8260 46116 8270
rect 46060 8166 46116 8204
rect 46396 8258 46452 8316
rect 46508 8370 46564 8540
rect 46508 8318 46510 8370
rect 46562 8318 46564 8370
rect 46508 8306 46564 8318
rect 46396 8206 46398 8258
rect 46450 8206 46452 8258
rect 46396 8194 46452 8206
rect 45724 7410 45780 7420
rect 46172 8148 46228 8158
rect 44380 7362 44436 7374
rect 44380 7310 44382 7362
rect 44434 7310 44436 7362
rect 44380 7028 44436 7310
rect 46172 7364 46228 8092
rect 46620 8036 46676 8046
rect 46620 7942 46676 7980
rect 46396 7476 46452 7486
rect 46396 7382 46452 7420
rect 46508 7364 46564 7374
rect 46172 7362 46340 7364
rect 46172 7310 46174 7362
rect 46226 7310 46340 7362
rect 46172 7308 46340 7310
rect 46172 7298 46228 7308
rect 44380 6962 44436 6972
rect 45724 7028 45780 7038
rect 44156 6804 44212 6814
rect 43596 6638 43598 6690
rect 43650 6638 43652 6690
rect 43596 6018 43652 6638
rect 44044 6692 44100 6702
rect 44044 6598 44100 6636
rect 44156 6690 44212 6748
rect 44156 6638 44158 6690
rect 44210 6638 44212 6690
rect 44156 6626 44212 6638
rect 43596 5966 43598 6018
rect 43650 5966 43652 6018
rect 43596 5954 43652 5966
rect 43708 6578 43764 6590
rect 43708 6526 43710 6578
rect 43762 6526 43764 6578
rect 43484 5236 43540 5246
rect 43484 5142 43540 5180
rect 43708 5236 43764 6526
rect 45724 6578 45780 6972
rect 45948 6804 46004 6814
rect 45948 6710 46004 6748
rect 45724 6526 45726 6578
rect 45778 6526 45780 6578
rect 45724 6514 45780 6526
rect 45836 6690 45892 6702
rect 45836 6638 45838 6690
rect 45890 6638 45892 6690
rect 44132 6300 44396 6310
rect 44188 6244 44236 6300
rect 44292 6244 44340 6300
rect 44132 6234 44396 6244
rect 44268 5906 44324 5918
rect 44268 5854 44270 5906
rect 44322 5854 44324 5906
rect 44268 5348 44324 5854
rect 44268 5282 44324 5292
rect 44716 5906 44772 5918
rect 44716 5854 44718 5906
rect 44770 5854 44772 5906
rect 43708 5142 43764 5180
rect 43708 4898 43764 4910
rect 43708 4846 43710 4898
rect 43762 4846 43764 4898
rect 43708 4788 43764 4846
rect 44716 4900 44772 5854
rect 45836 5794 45892 6638
rect 46284 6692 46340 7308
rect 46284 5906 46340 6636
rect 46284 5854 46286 5906
rect 46338 5854 46340 5906
rect 46284 5842 46340 5854
rect 46508 5906 46564 7308
rect 46508 5854 46510 5906
rect 46562 5854 46564 5906
rect 46508 5842 46564 5854
rect 46732 7364 46788 7374
rect 45836 5742 45838 5794
rect 45890 5742 45892 5794
rect 45388 5348 45444 5358
rect 44828 5236 44884 5246
rect 44828 5122 44884 5180
rect 44828 5070 44830 5122
rect 44882 5070 44884 5122
rect 44828 5058 44884 5070
rect 45164 4900 45220 4910
rect 44716 4834 44772 4844
rect 45052 4898 45220 4900
rect 45052 4846 45166 4898
rect 45218 4846 45220 4898
rect 45052 4844 45220 4846
rect 43764 4732 43988 4788
rect 43708 4722 43764 4732
rect 42812 4610 42868 4620
rect 43596 4676 43652 4686
rect 43260 4452 43316 4462
rect 43260 4358 43316 4396
rect 42140 4340 42196 4350
rect 41916 3668 41972 3678
rect 41804 3666 41972 3668
rect 41804 3614 41918 3666
rect 41970 3614 41972 3666
rect 41804 3612 41972 3614
rect 41916 3602 41972 3612
rect 41468 3556 41524 3566
rect 41132 3554 41524 3556
rect 41132 3502 41470 3554
rect 41522 3502 41524 3554
rect 41132 3500 41524 3502
rect 41468 3490 41524 3500
rect 41020 3390 41022 3442
rect 41074 3390 41076 3442
rect 41020 3378 41076 3390
rect 42140 3442 42196 4284
rect 42476 4338 42532 4350
rect 42476 4286 42478 4338
rect 42530 4286 42532 4338
rect 42476 4228 42532 4286
rect 42476 4162 42532 4172
rect 42588 3556 42644 3566
rect 43484 3556 43540 3566
rect 42588 3554 43540 3556
rect 42588 3502 42590 3554
rect 42642 3502 43486 3554
rect 43538 3502 43540 3554
rect 42588 3500 43540 3502
rect 42588 3490 42644 3500
rect 43484 3490 43540 3500
rect 42140 3390 42142 3442
rect 42194 3390 42196 3442
rect 42140 3378 42196 3390
rect 43596 3444 43652 4620
rect 43820 4228 43876 4238
rect 43820 3554 43876 4172
rect 43932 4226 43988 4732
rect 44132 4732 44396 4742
rect 44188 4676 44236 4732
rect 44292 4676 44340 4732
rect 44132 4666 44396 4676
rect 43932 4174 43934 4226
rect 43986 4174 43988 4226
rect 43932 4162 43988 4174
rect 44604 4450 44660 4462
rect 44604 4398 44606 4450
rect 44658 4398 44660 4450
rect 44604 3780 44660 4398
rect 44604 3714 44660 3724
rect 43820 3502 43822 3554
rect 43874 3502 43876 3554
rect 43820 3490 43876 3502
rect 45052 3554 45108 4844
rect 45164 4834 45220 4844
rect 45388 4338 45444 5292
rect 45388 4286 45390 4338
rect 45442 4286 45444 4338
rect 45388 4274 45444 4286
rect 45052 3502 45054 3554
rect 45106 3502 45108 3554
rect 45052 3490 45108 3502
rect 45724 4228 45780 4238
rect 43708 3444 43764 3454
rect 43596 3442 43764 3444
rect 43596 3390 43710 3442
rect 43762 3390 43764 3442
rect 43596 3388 43764 3390
rect 43708 3378 43764 3388
rect 45052 3332 45108 3342
rect 45052 3238 45108 3276
rect 44132 3164 44396 3174
rect 44188 3108 44236 3164
rect 44292 3108 44340 3164
rect 44132 3098 44396 3108
rect 45724 2772 45780 4172
rect 45836 3554 45892 5742
rect 46620 5122 46676 5134
rect 46620 5070 46622 5122
rect 46674 5070 46676 5122
rect 46620 4452 46676 5070
rect 46732 4562 46788 7308
rect 46844 7028 46900 8652
rect 47068 8260 47124 8270
rect 47180 8260 47236 10108
rect 47404 9826 47460 9838
rect 47404 9774 47406 9826
rect 47458 9774 47460 9826
rect 47404 9716 47460 9774
rect 47404 9266 47460 9660
rect 47404 9214 47406 9266
rect 47458 9214 47460 9266
rect 47404 9202 47460 9214
rect 47516 9268 47572 11228
rect 47628 11218 47684 11228
rect 48076 9602 48132 9614
rect 48076 9550 48078 9602
rect 48130 9550 48132 9602
rect 47516 9212 47796 9268
rect 47404 9044 47460 9054
rect 47292 8372 47348 8382
rect 47292 8278 47348 8316
rect 47404 8370 47460 8988
rect 47516 8930 47572 9212
rect 47516 8878 47518 8930
rect 47570 8878 47572 8930
rect 47516 8866 47572 8878
rect 47628 9042 47684 9054
rect 47628 8990 47630 9042
rect 47682 8990 47684 9042
rect 47404 8318 47406 8370
rect 47458 8318 47460 8370
rect 47404 8306 47460 8318
rect 47124 8204 47236 8260
rect 47068 8166 47124 8204
rect 47516 8148 47572 8186
rect 47516 8082 47572 8092
rect 47628 7698 47684 8990
rect 47628 7646 47630 7698
rect 47682 7646 47684 7698
rect 46956 7588 47012 7598
rect 46956 7494 47012 7532
rect 47628 7588 47684 7646
rect 47628 7522 47684 7532
rect 47516 7474 47572 7486
rect 47516 7422 47518 7474
rect 47570 7422 47572 7474
rect 47516 7364 47572 7422
rect 47740 7364 47796 9212
rect 48076 8148 48132 9550
rect 48188 9604 48244 9614
rect 48188 8258 48244 9548
rect 48412 9156 48468 15092
rect 48636 13860 48692 15036
rect 48748 14756 48804 16716
rect 48860 16436 48916 17390
rect 48972 17444 49028 18172
rect 49308 17778 49364 18172
rect 49308 17726 49310 17778
rect 49362 17726 49364 17778
rect 49308 17714 49364 17726
rect 49084 17556 49140 17566
rect 49084 17462 49140 17500
rect 48972 17378 49028 17388
rect 48860 16370 48916 16380
rect 48972 16882 49028 16894
rect 48972 16830 48974 16882
rect 49026 16830 49028 16882
rect 48972 16322 49028 16830
rect 49196 16882 49252 16894
rect 49196 16830 49198 16882
rect 49250 16830 49252 16882
rect 48972 16270 48974 16322
rect 49026 16270 49028 16322
rect 48972 16258 49028 16270
rect 49084 16770 49140 16782
rect 49084 16718 49086 16770
rect 49138 16718 49140 16770
rect 48860 16212 48916 16222
rect 48860 15202 48916 16156
rect 49084 15316 49140 16718
rect 49196 15988 49252 16830
rect 49308 16212 49364 16222
rect 49308 16118 49364 16156
rect 49196 15426 49252 15932
rect 49196 15374 49198 15426
rect 49250 15374 49252 15426
rect 49196 15362 49252 15374
rect 49084 15250 49140 15260
rect 48860 15150 48862 15202
rect 48914 15150 48916 15202
rect 48860 15138 48916 15150
rect 48748 14700 49252 14756
rect 48748 14532 48804 14542
rect 48748 14438 48804 14476
rect 48860 14420 48916 14430
rect 48860 14308 48916 14364
rect 48860 14306 49028 14308
rect 48860 14254 48862 14306
rect 48914 14254 49028 14306
rect 48860 14252 49028 14254
rect 48860 14242 48916 14252
rect 48748 13860 48804 13870
rect 48636 13858 48804 13860
rect 48636 13806 48750 13858
rect 48802 13806 48804 13858
rect 48636 13804 48804 13806
rect 48636 12850 48692 13804
rect 48748 13794 48804 13804
rect 48636 12798 48638 12850
rect 48690 12798 48692 12850
rect 48636 12786 48692 12798
rect 48860 13300 48916 13310
rect 48860 12402 48916 13244
rect 48972 13074 49028 14252
rect 49084 14306 49140 14318
rect 49084 14254 49086 14306
rect 49138 14254 49140 14306
rect 49084 13746 49140 14254
rect 49084 13694 49086 13746
rect 49138 13694 49140 13746
rect 49084 13682 49140 13694
rect 48972 13022 48974 13074
rect 49026 13022 49028 13074
rect 48972 13010 49028 13022
rect 48860 12350 48862 12402
rect 48914 12350 48916 12402
rect 48860 12338 48916 12350
rect 48748 11620 48804 11630
rect 48524 11172 48580 11182
rect 48524 11170 48692 11172
rect 48524 11118 48526 11170
rect 48578 11118 48692 11170
rect 48524 11116 48692 11118
rect 48524 11106 48580 11116
rect 48636 10052 48692 11116
rect 48748 10722 48804 11564
rect 48748 10670 48750 10722
rect 48802 10670 48804 10722
rect 48748 10658 48804 10670
rect 48748 10052 48804 10062
rect 48636 10050 48916 10052
rect 48636 9998 48750 10050
rect 48802 9998 48916 10050
rect 48636 9996 48916 9998
rect 48748 9986 48804 9996
rect 48524 9828 48580 9838
rect 48524 9734 48580 9772
rect 48412 9100 48804 9156
rect 48188 8206 48190 8258
rect 48242 8206 48244 8258
rect 48188 8194 48244 8206
rect 48524 8932 48580 8942
rect 48076 8082 48132 8092
rect 48300 8146 48356 8158
rect 48300 8094 48302 8146
rect 48354 8094 48356 8146
rect 48300 7812 48356 8094
rect 47852 7756 48356 7812
rect 47852 7698 47908 7756
rect 47852 7646 47854 7698
rect 47906 7646 47908 7698
rect 47852 7634 47908 7646
rect 48076 7476 48132 7486
rect 47516 7308 47796 7364
rect 47852 7420 48076 7476
rect 46844 6962 46900 6972
rect 46732 4510 46734 4562
rect 46786 4510 46788 4562
rect 46732 4498 46788 4510
rect 46956 6690 47012 6702
rect 46956 6638 46958 6690
rect 47010 6638 47012 6690
rect 46620 4386 46676 4396
rect 45836 3502 45838 3554
rect 45890 3502 45892 3554
rect 45836 3490 45892 3502
rect 45948 3780 46004 3790
rect 45948 3442 46004 3724
rect 46956 3780 47012 6638
rect 47740 6692 47796 6702
rect 47740 6598 47796 6636
rect 47852 6578 47908 7420
rect 48076 7382 48132 7420
rect 48188 7474 48244 7486
rect 48188 7422 48190 7474
rect 48242 7422 48244 7474
rect 48188 7252 48244 7422
rect 48188 7186 48244 7196
rect 47852 6526 47854 6578
rect 47906 6526 47908 6578
rect 47852 6514 47908 6526
rect 48076 6466 48132 6478
rect 48076 6414 48078 6466
rect 48130 6414 48132 6466
rect 47180 5908 47236 5918
rect 47180 5814 47236 5852
rect 47628 5908 47684 5918
rect 47628 5814 47684 5852
rect 47852 5796 47908 5806
rect 47852 5702 47908 5740
rect 47964 5460 48020 5470
rect 47964 5346 48020 5404
rect 47964 5294 47966 5346
rect 48018 5294 48020 5346
rect 47964 5282 48020 5294
rect 47180 5124 47236 5134
rect 48076 5124 48132 6414
rect 48188 5684 48244 5694
rect 48188 5590 48244 5628
rect 47180 5010 47236 5068
rect 47180 4958 47182 5010
rect 47234 4958 47236 5010
rect 47180 4946 47236 4958
rect 47964 5068 48076 5124
rect 47516 4452 47572 4462
rect 47404 4338 47460 4350
rect 47404 4286 47406 4338
rect 47458 4286 47460 4338
rect 46956 3714 47012 3724
rect 47068 4228 47124 4238
rect 47404 4228 47460 4286
rect 47068 4226 47460 4228
rect 47068 4174 47070 4226
rect 47122 4174 47460 4226
rect 47068 4172 47460 4174
rect 45948 3390 45950 3442
rect 46002 3390 46004 3442
rect 45948 3378 46004 3390
rect 45724 2706 45780 2716
rect 38444 2146 38500 2156
rect 47068 800 47124 4172
rect 47404 3780 47460 3790
rect 47404 3666 47460 3724
rect 47404 3614 47406 3666
rect 47458 3614 47460 3666
rect 47404 3602 47460 3614
rect 47516 3554 47572 4396
rect 47852 4228 47908 4238
rect 47852 4134 47908 4172
rect 47516 3502 47518 3554
rect 47570 3502 47572 3554
rect 47516 3490 47572 3502
rect 47964 3554 48020 5068
rect 48076 5058 48132 5068
rect 48524 5122 48580 8876
rect 48748 8708 48804 9100
rect 48860 9042 48916 9996
rect 48972 9826 49028 9838
rect 48972 9774 48974 9826
rect 49026 9774 49028 9826
rect 48972 9716 49028 9774
rect 49028 9660 49140 9716
rect 48972 9650 49028 9660
rect 48860 8990 48862 9042
rect 48914 8990 48916 9042
rect 48860 8978 48916 8990
rect 49084 9042 49140 9660
rect 49084 8990 49086 9042
rect 49138 8990 49140 9042
rect 49084 8978 49140 8990
rect 48748 8652 48916 8708
rect 48748 8148 48804 8158
rect 48748 8054 48804 8092
rect 48748 7924 48804 7934
rect 48748 5908 48804 7868
rect 48860 6690 48916 8652
rect 49196 7476 49252 14700
rect 49420 14642 49476 19068
rect 49532 19012 49588 19182
rect 49532 18564 49588 18956
rect 49532 18498 49588 18508
rect 49532 18340 49588 18350
rect 49644 18340 49700 19740
rect 50204 19684 50260 19966
rect 50540 20018 50596 20030
rect 51100 20020 51156 21308
rect 51286 21196 51550 21206
rect 51342 21140 51390 21196
rect 51446 21140 51494 21196
rect 51286 21130 51550 21140
rect 51548 21028 51604 21038
rect 51212 20916 51268 20926
rect 51268 20860 51380 20916
rect 51212 20850 51268 20860
rect 51212 20578 51268 20590
rect 51212 20526 51214 20578
rect 51266 20526 51268 20578
rect 51212 20132 51268 20526
rect 51324 20242 51380 20860
rect 51548 20914 51604 20972
rect 51548 20862 51550 20914
rect 51602 20862 51604 20914
rect 51548 20850 51604 20862
rect 51996 20578 52052 20590
rect 51996 20526 51998 20578
rect 52050 20526 52052 20578
rect 51996 20468 52052 20526
rect 51996 20402 52052 20412
rect 51324 20190 51326 20242
rect 51378 20190 51380 20242
rect 51324 20178 51380 20190
rect 51212 20066 51268 20076
rect 51996 20132 52052 20142
rect 50540 19966 50542 20018
rect 50594 19966 50596 20018
rect 50428 19684 50484 19694
rect 50204 19628 50372 19684
rect 49980 19572 50036 19582
rect 49756 19124 49812 19134
rect 49756 19030 49812 19068
rect 49980 18788 50036 19516
rect 50204 19460 50260 19470
rect 50204 19346 50260 19404
rect 50204 19294 50206 19346
rect 50258 19294 50260 19346
rect 50204 19282 50260 19294
rect 49532 18338 49700 18340
rect 49532 18286 49534 18338
rect 49586 18286 49700 18338
rect 49532 18284 49700 18286
rect 49868 18732 50036 18788
rect 50316 19124 50372 19628
rect 50428 19124 50484 19628
rect 50540 19348 50596 19966
rect 50876 19964 51156 20020
rect 50540 19282 50596 19292
rect 50764 19794 50820 19806
rect 50764 19742 50766 19794
rect 50818 19742 50820 19794
rect 50764 19236 50820 19742
rect 50652 19234 50820 19236
rect 50652 19182 50766 19234
rect 50818 19182 50820 19234
rect 50652 19180 50820 19182
rect 50428 19068 50596 19124
rect 49868 18450 49924 18732
rect 49980 18564 50036 18574
rect 49980 18562 50148 18564
rect 49980 18510 49982 18562
rect 50034 18510 50148 18562
rect 49980 18508 50148 18510
rect 49980 18498 50036 18508
rect 49868 18398 49870 18450
rect 49922 18398 49924 18450
rect 49868 18340 49924 18398
rect 49868 18284 50036 18340
rect 49532 18274 49588 18284
rect 49532 17666 49588 17678
rect 49532 17614 49534 17666
rect 49586 17614 49588 17666
rect 49532 17444 49588 17614
rect 49532 17378 49588 17388
rect 49868 17442 49924 17454
rect 49868 17390 49870 17442
rect 49922 17390 49924 17442
rect 49868 17108 49924 17390
rect 49868 17042 49924 17052
rect 49980 16996 50036 18284
rect 50092 18228 50148 18508
rect 50204 18452 50260 18462
rect 50204 18358 50260 18396
rect 50092 18162 50148 18172
rect 49980 16930 50036 16940
rect 50092 17444 50148 17454
rect 49644 16884 49700 16894
rect 49644 16882 49924 16884
rect 49644 16830 49646 16882
rect 49698 16830 49924 16882
rect 49644 16828 49924 16830
rect 49644 16818 49700 16828
rect 49868 16322 49924 16828
rect 49980 16772 50036 16782
rect 50092 16772 50148 17388
rect 49980 16770 50148 16772
rect 49980 16718 49982 16770
rect 50034 16718 50148 16770
rect 49980 16716 50148 16718
rect 50204 17442 50260 17454
rect 50204 17390 50206 17442
rect 50258 17390 50260 17442
rect 49980 16706 50036 16716
rect 49868 16270 49870 16322
rect 49922 16270 49924 16322
rect 49868 16258 49924 16270
rect 49532 16100 49588 16110
rect 50092 16100 50148 16110
rect 49532 16006 49588 16044
rect 49980 16098 50148 16100
rect 49980 16046 50094 16098
rect 50146 16046 50148 16098
rect 49980 16044 50148 16046
rect 49980 15988 50036 16044
rect 50092 16034 50148 16044
rect 49980 15922 50036 15932
rect 50204 15148 50260 17390
rect 50316 16884 50372 19068
rect 50540 18674 50596 19068
rect 50540 18622 50542 18674
rect 50594 18622 50596 18674
rect 50428 18564 50484 18574
rect 50428 18470 50484 18508
rect 50540 18340 50596 18622
rect 50428 18284 50596 18340
rect 50428 17220 50484 18284
rect 50540 17892 50596 17902
rect 50652 17892 50708 19180
rect 50764 19170 50820 19180
rect 50876 19236 50932 19964
rect 51772 19906 51828 19918
rect 51772 19854 51774 19906
rect 51826 19854 51828 19906
rect 51772 19796 51828 19854
rect 51772 19794 51940 19796
rect 51772 19742 51774 19794
rect 51826 19742 51940 19794
rect 51772 19740 51940 19742
rect 51772 19730 51828 19740
rect 51286 19628 51550 19638
rect 51342 19572 51390 19628
rect 51446 19572 51494 19628
rect 51286 19562 51550 19572
rect 51548 19348 51604 19358
rect 50876 19180 51268 19236
rect 50876 19122 50932 19180
rect 50876 19070 50878 19122
rect 50930 19070 50932 19122
rect 50876 19058 50932 19070
rect 51100 19012 51156 19022
rect 50988 19010 51156 19012
rect 50988 18958 51102 19010
rect 51154 18958 51156 19010
rect 50988 18956 51156 18958
rect 50764 18452 50820 18462
rect 50764 18358 50820 18396
rect 50540 17890 50708 17892
rect 50540 17838 50542 17890
rect 50594 17838 50708 17890
rect 50540 17836 50708 17838
rect 50540 17826 50596 17836
rect 50428 17106 50484 17164
rect 50428 17054 50430 17106
rect 50482 17054 50484 17106
rect 50428 17042 50484 17054
rect 50316 16828 50484 16884
rect 50316 16436 50372 16446
rect 50316 15986 50372 16380
rect 50316 15934 50318 15986
rect 50370 15934 50372 15986
rect 50316 15922 50372 15934
rect 50428 15986 50484 16828
rect 50652 16772 50708 17836
rect 50652 16706 50708 16716
rect 50764 17666 50820 17678
rect 50764 17614 50766 17666
rect 50818 17614 50820 17666
rect 50764 17332 50820 17614
rect 50988 17444 51044 18956
rect 51100 18946 51156 18956
rect 51100 18676 51156 18686
rect 51212 18676 51268 19180
rect 51100 18674 51268 18676
rect 51100 18622 51102 18674
rect 51154 18622 51268 18674
rect 51100 18620 51268 18622
rect 51100 18610 51156 18620
rect 51548 18338 51604 19292
rect 51772 19236 51828 19246
rect 51772 19142 51828 19180
rect 51548 18286 51550 18338
rect 51602 18286 51604 18338
rect 51548 18274 51604 18286
rect 51286 18060 51550 18070
rect 51342 18004 51390 18060
rect 51446 18004 51494 18060
rect 51286 17994 51550 18004
rect 51772 17780 51828 17790
rect 51884 17780 51940 19740
rect 51996 18562 52052 20076
rect 52108 19796 52164 25004
rect 52220 24836 52276 24846
rect 52220 24722 52276 24780
rect 52220 24670 52222 24722
rect 52274 24670 52276 24722
rect 52220 24658 52276 24670
rect 52556 24724 52612 24734
rect 52556 23938 52612 24668
rect 53116 24724 53172 25230
rect 53340 25284 53396 25294
rect 53340 25190 53396 25228
rect 53116 24164 53172 24668
rect 53116 24098 53172 24108
rect 53452 24834 53508 25340
rect 53452 24782 53454 24834
rect 53506 24782 53508 24834
rect 53340 24052 53396 24062
rect 53340 23958 53396 23996
rect 52556 23886 52558 23938
rect 52610 23886 52612 23938
rect 52556 23874 52612 23886
rect 52892 23828 52948 23838
rect 52892 23734 52948 23772
rect 52780 23716 52836 23726
rect 52780 23622 52836 23660
rect 53452 23492 53508 24782
rect 53340 23436 53508 23492
rect 52444 23042 52500 23054
rect 52444 22990 52446 23042
rect 52498 22990 52500 23042
rect 52220 22930 52276 22942
rect 52220 22878 52222 22930
rect 52274 22878 52276 22930
rect 52220 21924 52276 22878
rect 52444 22260 52500 22990
rect 52892 22372 52948 22382
rect 53228 22372 53284 22382
rect 52948 22370 53284 22372
rect 52948 22318 53230 22370
rect 53282 22318 53284 22370
rect 52948 22316 53284 22318
rect 52892 22278 52948 22316
rect 53228 22306 53284 22316
rect 52444 22194 52500 22204
rect 52220 21586 52276 21868
rect 52220 21534 52222 21586
rect 52274 21534 52276 21586
rect 52220 21522 52276 21534
rect 53116 22148 53172 22158
rect 53116 21586 53172 22092
rect 53116 21534 53118 21586
rect 53170 21534 53172 21586
rect 53116 21522 53172 21534
rect 53116 20802 53172 20814
rect 53116 20750 53118 20802
rect 53170 20750 53172 20802
rect 52892 20692 52948 20702
rect 52892 20580 52948 20636
rect 52668 20524 52948 20580
rect 52108 19730 52164 19740
rect 52444 20018 52500 20030
rect 52444 19966 52446 20018
rect 52498 19966 52500 20018
rect 52108 19460 52164 19470
rect 52444 19460 52500 19966
rect 52556 20020 52612 20030
rect 52668 20020 52724 20524
rect 53116 20244 53172 20750
rect 53116 20178 53172 20188
rect 52780 20132 52836 20142
rect 53004 20132 53060 20142
rect 52836 20076 52948 20132
rect 52780 20066 52836 20076
rect 52612 19964 52724 20020
rect 52892 20018 52948 20076
rect 53004 20038 53060 20076
rect 52892 19966 52894 20018
rect 52946 19966 52948 20018
rect 52556 19954 52612 19964
rect 52892 19954 52948 19966
rect 53116 20018 53172 20030
rect 53116 19966 53118 20018
rect 53170 19966 53172 20018
rect 52108 19458 52500 19460
rect 52108 19406 52110 19458
rect 52162 19406 52500 19458
rect 52108 19404 52500 19406
rect 53116 19460 53172 19966
rect 53228 19460 53284 19470
rect 53116 19458 53284 19460
rect 53116 19406 53230 19458
rect 53282 19406 53284 19458
rect 53116 19404 53284 19406
rect 52108 19394 52164 19404
rect 53228 19394 53284 19404
rect 52668 19348 52724 19358
rect 52668 19254 52724 19292
rect 51996 18510 51998 18562
rect 52050 18510 52052 18562
rect 51996 18498 52052 18510
rect 52892 19236 52948 19246
rect 52892 18452 52948 19180
rect 53004 18452 53060 18462
rect 52892 18450 53060 18452
rect 52892 18398 53006 18450
rect 53058 18398 53060 18450
rect 52892 18396 53060 18398
rect 53004 18386 53060 18396
rect 53340 17890 53396 23436
rect 53676 21810 53732 21822
rect 53676 21758 53678 21810
rect 53730 21758 53732 21810
rect 53676 21700 53732 21758
rect 53676 21634 53732 21644
rect 53900 21140 53956 26796
rect 54012 26628 54068 27468
rect 54012 26562 54068 26572
rect 54124 26964 54180 26974
rect 54012 26404 54068 26414
rect 54012 25730 54068 26348
rect 54124 26180 54180 26908
rect 54124 26114 54180 26124
rect 54012 25678 54014 25730
rect 54066 25678 54068 25730
rect 54012 24722 54068 25678
rect 54236 25396 54292 25406
rect 54236 25302 54292 25340
rect 54124 25284 54180 25294
rect 54124 25190 54180 25228
rect 54572 24948 54628 27692
rect 54684 26180 54740 27806
rect 55132 27860 55188 27870
rect 55468 27860 55524 27870
rect 54796 27636 54852 27646
rect 54796 27188 54852 27580
rect 55132 27300 55188 27804
rect 54796 26962 54852 27132
rect 54796 26910 54798 26962
rect 54850 26910 54852 26962
rect 54796 26898 54852 26910
rect 55020 27244 55188 27300
rect 55244 27858 55524 27860
rect 55244 27806 55470 27858
rect 55522 27806 55524 27858
rect 55244 27804 55524 27806
rect 55020 26908 55076 27244
rect 54908 26852 55076 26908
rect 55132 27074 55188 27086
rect 55132 27022 55134 27074
rect 55186 27022 55188 27074
rect 54796 26404 54852 26414
rect 54908 26404 54964 26852
rect 55132 26628 55188 27022
rect 55132 26562 55188 26572
rect 54796 26402 54964 26404
rect 54796 26350 54798 26402
rect 54850 26350 54964 26402
rect 54796 26348 54964 26350
rect 54796 26338 54852 26348
rect 55132 26292 55188 26302
rect 55244 26292 55300 27804
rect 55468 27794 55524 27804
rect 55916 26908 55972 29148
rect 56364 28644 56420 28654
rect 56364 28550 56420 28588
rect 56924 28532 56980 29486
rect 57148 29314 57204 30268
rect 57148 29262 57150 29314
rect 57202 29262 57204 29314
rect 57148 29250 57204 29262
rect 56924 28466 56980 28476
rect 57260 28082 57316 31726
rect 57372 30882 57428 30894
rect 57372 30830 57374 30882
rect 57426 30830 57428 30882
rect 57372 30212 57428 30830
rect 57372 30146 57428 30156
rect 57484 29764 57540 32510
rect 58044 31108 58100 33292
rect 58156 32788 58212 32798
rect 58268 32788 58324 34972
rect 58439 34524 58703 34534
rect 58495 34468 58543 34524
rect 58599 34468 58647 34524
rect 58439 34458 58703 34468
rect 58439 32956 58703 32966
rect 58495 32900 58543 32956
rect 58599 32900 58647 32956
rect 58439 32890 58703 32900
rect 58156 32786 58324 32788
rect 58156 32734 58158 32786
rect 58210 32734 58324 32786
rect 58156 32732 58324 32734
rect 58156 32722 58212 32732
rect 58268 32676 58324 32732
rect 58044 31014 58100 31052
rect 58156 31892 58212 31902
rect 58156 30884 58212 31836
rect 58044 30828 58212 30884
rect 57932 30210 57988 30222
rect 57932 30158 57934 30210
rect 57986 30158 57988 30210
rect 57596 30100 57652 30110
rect 57596 30006 57652 30044
rect 57708 29986 57764 29998
rect 57708 29934 57710 29986
rect 57762 29934 57764 29986
rect 57484 29708 57652 29764
rect 57260 28030 57262 28082
rect 57314 28030 57316 28082
rect 57260 28018 57316 28030
rect 57372 28532 57428 28542
rect 57036 27858 57092 27870
rect 57036 27806 57038 27858
rect 57090 27806 57092 27858
rect 56028 27076 56084 27086
rect 56028 26982 56084 27020
rect 56700 26964 56756 26974
rect 56700 26962 56868 26964
rect 56700 26910 56702 26962
rect 56754 26910 56868 26962
rect 56700 26908 56868 26910
rect 55916 26852 56084 26908
rect 56700 26898 56756 26908
rect 55132 26290 55300 26292
rect 55132 26238 55134 26290
rect 55186 26238 55300 26290
rect 55132 26236 55300 26238
rect 55132 26226 55188 26236
rect 54908 26180 54964 26190
rect 54684 26178 54964 26180
rect 54684 26126 54910 26178
rect 54962 26126 54964 26178
rect 54684 26124 54964 26126
rect 54908 26114 54964 26124
rect 55132 25508 55188 25546
rect 55132 25442 55188 25452
rect 54572 24892 54852 24948
rect 54012 24670 54014 24722
rect 54066 24670 54068 24722
rect 54012 24658 54068 24670
rect 54684 24724 54740 24734
rect 54684 24630 54740 24668
rect 54684 24500 54740 24510
rect 54348 23156 54404 23166
rect 54348 23062 54404 23100
rect 54460 23044 54516 23054
rect 54236 22932 54292 22942
rect 54236 22370 54292 22876
rect 54460 22482 54516 22988
rect 54460 22430 54462 22482
rect 54514 22430 54516 22482
rect 54460 22418 54516 22430
rect 54236 22318 54238 22370
rect 54290 22318 54292 22370
rect 54236 22306 54292 22318
rect 54348 21812 54404 21822
rect 54348 21718 54404 21756
rect 54460 21698 54516 21710
rect 54460 21646 54462 21698
rect 54514 21646 54516 21698
rect 54236 21362 54292 21374
rect 54236 21310 54238 21362
rect 54290 21310 54292 21362
rect 53900 21084 54068 21140
rect 53452 20916 53508 20926
rect 53900 20916 53956 20926
rect 53452 20914 53956 20916
rect 53452 20862 53454 20914
rect 53506 20862 53902 20914
rect 53954 20862 53956 20914
rect 53452 20860 53956 20862
rect 53452 20850 53508 20860
rect 53564 20580 53620 20590
rect 53564 19458 53620 20524
rect 53900 20130 53956 20860
rect 53900 20078 53902 20130
rect 53954 20078 53956 20130
rect 53900 20066 53956 20078
rect 53564 19406 53566 19458
rect 53618 19406 53620 19458
rect 53564 19394 53620 19406
rect 53788 19908 53844 19918
rect 53788 19122 53844 19852
rect 53900 19460 53956 19470
rect 53900 19366 53956 19404
rect 53788 19070 53790 19122
rect 53842 19070 53844 19122
rect 53340 17838 53342 17890
rect 53394 17838 53396 17890
rect 53340 17826 53396 17838
rect 53676 18338 53732 18350
rect 53676 18286 53678 18338
rect 53730 18286 53732 18338
rect 51100 17778 51940 17780
rect 51100 17726 51774 17778
rect 51826 17726 51940 17778
rect 51100 17724 51940 17726
rect 51100 17666 51156 17724
rect 51100 17614 51102 17666
rect 51154 17614 51156 17666
rect 51100 17602 51156 17614
rect 51212 17444 51268 17454
rect 50988 17378 51044 17388
rect 51100 17442 51268 17444
rect 51100 17390 51214 17442
rect 51266 17390 51268 17442
rect 51100 17388 51268 17390
rect 50764 16212 50820 17276
rect 50876 17220 50932 17230
rect 51100 17220 51156 17388
rect 51212 17378 51268 17388
rect 51436 17442 51492 17454
rect 51436 17390 51438 17442
rect 51490 17390 51492 17442
rect 50932 17164 51156 17220
rect 50876 17154 50932 17164
rect 50988 16322 51044 17164
rect 51212 17108 51268 17118
rect 51212 16884 51268 17052
rect 50988 16270 50990 16322
rect 51042 16270 51044 16322
rect 50988 16258 51044 16270
rect 51100 16882 51268 16884
rect 51100 16830 51214 16882
rect 51266 16830 51268 16882
rect 51100 16828 51268 16830
rect 50876 16212 50932 16222
rect 50764 16210 50932 16212
rect 50764 16158 50878 16210
rect 50930 16158 50932 16210
rect 50764 16156 50932 16158
rect 50876 16146 50932 16156
rect 50428 15934 50430 15986
rect 50482 15934 50484 15986
rect 50428 15428 50484 15934
rect 50428 15362 50484 15372
rect 50652 16100 50708 16110
rect 50652 15426 50708 16044
rect 50652 15374 50654 15426
rect 50706 15374 50708 15426
rect 50652 15362 50708 15374
rect 50988 15202 51044 15214
rect 50988 15150 50990 15202
rect 51042 15150 51044 15202
rect 50988 15148 51044 15150
rect 50092 15092 50260 15148
rect 50540 15092 51044 15148
rect 49420 14590 49422 14642
rect 49474 14590 49476 14642
rect 49420 13412 49476 14590
rect 49868 14980 49924 14990
rect 49868 14642 49924 14924
rect 49868 14590 49870 14642
rect 49922 14590 49924 14642
rect 49868 14578 49924 14590
rect 49644 14308 49700 14318
rect 49644 13746 49700 14252
rect 49644 13694 49646 13746
rect 49698 13694 49700 13746
rect 49644 13682 49700 13694
rect 49756 13970 49812 13982
rect 49756 13918 49758 13970
rect 49810 13918 49812 13970
rect 49420 13346 49476 13356
rect 49532 12964 49588 12974
rect 49308 12908 49532 12964
rect 49308 11396 49364 12908
rect 49532 12870 49588 12908
rect 49756 12850 49812 13918
rect 49868 13076 49924 13086
rect 49868 13074 50036 13076
rect 49868 13022 49870 13074
rect 49922 13022 50036 13074
rect 49868 13020 50036 13022
rect 49868 13010 49924 13020
rect 49756 12798 49758 12850
rect 49810 12798 49812 12850
rect 49420 12178 49476 12190
rect 49420 12126 49422 12178
rect 49474 12126 49476 12178
rect 49420 11732 49476 12126
rect 49756 12068 49812 12798
rect 49420 11666 49476 11676
rect 49532 12066 49812 12068
rect 49532 12014 49758 12066
rect 49810 12014 49812 12066
rect 49532 12012 49812 12014
rect 49420 11396 49476 11406
rect 49308 11394 49476 11396
rect 49308 11342 49422 11394
rect 49474 11342 49476 11394
rect 49308 11340 49476 11342
rect 49420 11330 49476 11340
rect 49532 11282 49588 12012
rect 49756 12002 49812 12012
rect 49756 11396 49812 11406
rect 49756 11302 49812 11340
rect 49980 11394 50036 13020
rect 50092 11732 50148 15092
rect 50204 14644 50260 14654
rect 50204 12962 50260 14588
rect 50428 13860 50484 13870
rect 50316 13636 50372 13646
rect 50316 13542 50372 13580
rect 50204 12910 50206 12962
rect 50258 12910 50260 12962
rect 50204 12898 50260 12910
rect 50428 12962 50484 13804
rect 50428 12910 50430 12962
rect 50482 12910 50484 12962
rect 50428 12898 50484 12910
rect 50540 12964 50596 15092
rect 50540 12898 50596 12908
rect 50652 14980 50708 14990
rect 50652 14644 50708 14924
rect 51100 14756 51156 16828
rect 51212 16818 51268 16828
rect 51436 16770 51492 17390
rect 51436 16718 51438 16770
rect 51490 16718 51492 16770
rect 51436 16706 51492 16718
rect 51286 16492 51550 16502
rect 51342 16436 51390 16492
rect 51446 16436 51494 16492
rect 51286 16426 51550 16436
rect 51324 16322 51380 16334
rect 51324 16270 51326 16322
rect 51378 16270 51380 16322
rect 51324 16210 51380 16270
rect 51548 16324 51604 16334
rect 51604 16268 51716 16324
rect 51548 16258 51604 16268
rect 51324 16158 51326 16210
rect 51378 16158 51380 16210
rect 51324 16146 51380 16158
rect 51548 15316 51604 15326
rect 51548 15222 51604 15260
rect 51660 15204 51716 16268
rect 51772 16210 51828 17724
rect 53116 17668 53172 17678
rect 52780 16882 52836 16894
rect 52780 16830 52782 16882
rect 52834 16830 52836 16882
rect 51884 16772 51940 16782
rect 51884 16678 51940 16716
rect 52780 16660 52836 16830
rect 52780 16594 52836 16604
rect 52892 16772 52948 16782
rect 51772 16158 51774 16210
rect 51826 16158 51828 16210
rect 51772 16146 51828 16158
rect 52668 15988 52724 15998
rect 52444 15986 52724 15988
rect 52444 15934 52670 15986
rect 52722 15934 52724 15986
rect 52444 15932 52724 15934
rect 52444 15428 52500 15932
rect 52668 15922 52724 15932
rect 52892 15988 52948 16716
rect 53116 16770 53172 17612
rect 53116 16718 53118 16770
rect 53170 16718 53172 16770
rect 53116 16706 53172 16718
rect 53340 17666 53396 17678
rect 53340 17614 53342 17666
rect 53394 17614 53396 17666
rect 53340 16660 53396 17614
rect 53564 16884 53620 16894
rect 53564 16770 53620 16828
rect 53564 16718 53566 16770
rect 53618 16718 53620 16770
rect 53564 16706 53620 16718
rect 53340 16594 53396 16604
rect 53676 16436 53732 18286
rect 53564 16380 53732 16436
rect 53004 16212 53060 16222
rect 53004 16210 53172 16212
rect 53004 16158 53006 16210
rect 53058 16158 53172 16210
rect 53004 16156 53172 16158
rect 53004 16146 53060 16156
rect 52892 15986 53060 15988
rect 52892 15934 52894 15986
rect 52946 15934 53060 15986
rect 52892 15932 53060 15934
rect 52892 15922 52948 15932
rect 52444 15334 52500 15372
rect 52892 15316 52948 15326
rect 51660 15138 51716 15148
rect 52556 15204 52612 15214
rect 51286 14924 51550 14934
rect 51342 14868 51390 14924
rect 51446 14868 51494 14924
rect 51286 14858 51550 14868
rect 51156 14700 51380 14756
rect 51100 14662 51156 14700
rect 50988 14644 51044 14654
rect 50652 14642 51044 14644
rect 50652 14590 50654 14642
rect 50706 14590 50990 14642
rect 51042 14590 51044 14642
rect 50652 14588 51044 14590
rect 50652 12850 50708 14588
rect 50988 14578 51044 14588
rect 51324 14530 51380 14700
rect 51324 14478 51326 14530
rect 51378 14478 51380 14530
rect 51324 14466 51380 14478
rect 51772 14530 51828 14542
rect 51772 14478 51774 14530
rect 51826 14478 51828 14530
rect 51100 14420 51156 14430
rect 51100 14418 51268 14420
rect 51100 14366 51102 14418
rect 51154 14366 51268 14418
rect 51100 14364 51268 14366
rect 51100 14354 51156 14364
rect 51100 13860 51156 13870
rect 50764 13858 51156 13860
rect 50764 13806 51102 13858
rect 51154 13806 51156 13858
rect 50764 13804 51156 13806
rect 50764 13186 50820 13804
rect 51100 13794 51156 13804
rect 51212 13524 51268 14364
rect 50764 13134 50766 13186
rect 50818 13134 50820 13186
rect 50764 13122 50820 13134
rect 51100 13468 51268 13524
rect 51660 13746 51716 13758
rect 51660 13694 51662 13746
rect 51714 13694 51716 13746
rect 50652 12798 50654 12850
rect 50706 12798 50708 12850
rect 50652 12786 50708 12798
rect 50764 12964 50820 12974
rect 50764 12178 50820 12908
rect 51100 12852 51156 13468
rect 51286 13356 51550 13366
rect 51342 13300 51390 13356
rect 51446 13300 51494 13356
rect 51286 13290 51550 13300
rect 51100 12786 51156 12796
rect 51212 12962 51268 12974
rect 51212 12910 51214 12962
rect 51266 12910 51268 12962
rect 51212 12292 51268 12910
rect 51212 12226 51268 12236
rect 51436 12964 51492 12974
rect 51660 12964 51716 13694
rect 51772 13636 51828 14478
rect 51996 14532 52052 14542
rect 51996 14438 52052 14476
rect 52556 14530 52612 15148
rect 52780 15204 52836 15214
rect 52780 14642 52836 15148
rect 52780 14590 52782 14642
rect 52834 14590 52836 14642
rect 52780 14578 52836 14590
rect 52556 14478 52558 14530
rect 52610 14478 52612 14530
rect 52556 14466 52612 14478
rect 52892 14530 52948 15260
rect 53004 15314 53060 15932
rect 53004 15262 53006 15314
rect 53058 15262 53060 15314
rect 53004 15250 53060 15262
rect 52892 14478 52894 14530
rect 52946 14478 52948 14530
rect 52892 14466 52948 14478
rect 53116 14530 53172 16156
rect 53228 15428 53284 15438
rect 53228 15202 53284 15372
rect 53228 15150 53230 15202
rect 53282 15150 53284 15202
rect 53228 15138 53284 15150
rect 53564 15148 53620 16380
rect 53788 16324 53844 19070
rect 53116 14478 53118 14530
rect 53170 14478 53172 14530
rect 53116 14466 53172 14478
rect 53452 15092 53620 15148
rect 53676 16268 53844 16324
rect 52444 14196 52500 14206
rect 52332 13748 52388 13758
rect 51772 13188 51828 13580
rect 52220 13746 52388 13748
rect 52220 13694 52334 13746
rect 52386 13694 52388 13746
rect 52220 13692 52388 13694
rect 51772 13132 52052 13188
rect 51996 13076 52052 13132
rect 52108 13076 52164 13086
rect 51996 13074 52164 13076
rect 51996 13022 52110 13074
rect 52162 13022 52164 13074
rect 51996 13020 52164 13022
rect 52108 13010 52164 13020
rect 51436 12962 51716 12964
rect 51436 12910 51438 12962
rect 51490 12910 51716 12962
rect 51436 12908 51716 12910
rect 50764 12126 50766 12178
rect 50818 12126 50820 12178
rect 50764 12114 50820 12126
rect 51100 12068 51156 12078
rect 50764 11956 50820 11966
rect 50092 11666 50148 11676
rect 50652 11732 50708 11742
rect 49980 11342 49982 11394
rect 50034 11342 50036 11394
rect 49980 11330 50036 11342
rect 50540 11396 50596 11406
rect 50540 11302 50596 11340
rect 49532 11230 49534 11282
rect 49586 11230 49588 11282
rect 49532 11218 49588 11230
rect 50652 11282 50708 11676
rect 50652 11230 50654 11282
rect 50706 11230 50708 11282
rect 50652 11218 50708 11230
rect 49308 10610 49364 10622
rect 49308 10558 49310 10610
rect 49362 10558 49364 10610
rect 49308 9826 49364 10558
rect 49308 9774 49310 9826
rect 49362 9774 49364 9826
rect 49308 8370 49364 9774
rect 49308 8318 49310 8370
rect 49362 8318 49364 8370
rect 49308 8306 49364 8318
rect 49532 10498 49588 10510
rect 49532 10446 49534 10498
rect 49586 10446 49588 10498
rect 49532 9826 49588 10446
rect 50652 10052 50708 10062
rect 50652 9958 50708 9996
rect 49532 9774 49534 9826
rect 49586 9774 49588 9826
rect 49532 8258 49588 9774
rect 49756 9828 49812 9838
rect 49756 9156 49812 9772
rect 50540 9826 50596 9838
rect 50764 9828 50820 11900
rect 50988 11506 51044 11518
rect 50988 11454 50990 11506
rect 51042 11454 51044 11506
rect 50988 10052 51044 11454
rect 51100 11284 51156 12012
rect 51436 11956 51492 12908
rect 52108 12292 52164 12302
rect 52220 12292 52276 13692
rect 52332 13682 52388 13692
rect 52164 12236 52276 12292
rect 52332 12290 52388 12302
rect 52332 12238 52334 12290
rect 52386 12238 52388 12290
rect 51548 12068 51604 12078
rect 51772 12068 51828 12078
rect 51548 12066 51716 12068
rect 51548 12014 51550 12066
rect 51602 12014 51716 12066
rect 51548 12012 51716 12014
rect 51548 12002 51604 12012
rect 51436 11890 51492 11900
rect 51286 11788 51550 11798
rect 51342 11732 51390 11788
rect 51446 11732 51494 11788
rect 51286 11722 51550 11732
rect 51548 11620 51604 11630
rect 51660 11620 51716 12012
rect 51548 11618 51716 11620
rect 51548 11566 51550 11618
rect 51602 11566 51716 11618
rect 51548 11564 51716 11566
rect 51100 11228 51380 11284
rect 51324 10610 51380 11228
rect 51324 10558 51326 10610
rect 51378 10558 51380 10610
rect 51324 10546 51380 10558
rect 51548 10498 51604 11564
rect 51772 11282 51828 12012
rect 52108 12066 52164 12236
rect 52108 12014 52110 12066
rect 52162 12014 52164 12066
rect 52108 12002 52164 12014
rect 52332 11956 52388 12238
rect 52332 11890 52388 11900
rect 51772 11230 51774 11282
rect 51826 11230 51828 11282
rect 51772 11218 51828 11230
rect 51548 10446 51550 10498
rect 51602 10446 51604 10498
rect 51548 10434 51604 10446
rect 51660 11170 51716 11182
rect 51660 11118 51662 11170
rect 51714 11118 51716 11170
rect 51286 10220 51550 10230
rect 51342 10164 51390 10220
rect 51446 10164 51494 10220
rect 51286 10154 51550 10164
rect 50988 9996 51156 10052
rect 50540 9774 50542 9826
rect 50594 9774 50596 9826
rect 49756 9042 49812 9100
rect 49756 8990 49758 9042
rect 49810 8990 49812 9042
rect 49756 8978 49812 8990
rect 50204 9380 50260 9390
rect 49532 8206 49534 8258
rect 49586 8206 49588 8258
rect 49532 8194 49588 8206
rect 49980 8820 50036 8830
rect 49980 8258 50036 8764
rect 50204 8370 50260 9324
rect 50540 9268 50596 9774
rect 50316 9212 50596 9268
rect 50652 9772 50820 9828
rect 50988 9826 51044 9838
rect 50988 9774 50990 9826
rect 51042 9774 51044 9826
rect 50316 8820 50372 9212
rect 50316 8754 50372 8764
rect 50204 8318 50206 8370
rect 50258 8318 50260 8370
rect 50204 8306 50260 8318
rect 49980 8206 49982 8258
rect 50034 8206 50036 8258
rect 49980 8194 50036 8206
rect 49196 7362 49252 7420
rect 49532 7588 49588 7598
rect 49532 7474 49588 7532
rect 50316 7588 50372 7598
rect 50316 7494 50372 7532
rect 49532 7422 49534 7474
rect 49586 7422 49588 7474
rect 49532 7410 49588 7422
rect 50540 7476 50596 7486
rect 50540 7382 50596 7420
rect 49196 7310 49198 7362
rect 49250 7310 49252 7362
rect 49196 7298 49252 7310
rect 49532 7250 49588 7262
rect 49532 7198 49534 7250
rect 49586 7198 49588 7250
rect 48860 6638 48862 6690
rect 48914 6638 48916 6690
rect 48860 6580 48916 6638
rect 48860 6514 48916 6524
rect 49308 6914 49364 6926
rect 49308 6862 49310 6914
rect 49362 6862 49364 6914
rect 48860 5908 48916 5918
rect 49308 5908 49364 6862
rect 49532 6804 49588 7198
rect 50092 6804 50148 6814
rect 49532 6802 50148 6804
rect 49532 6750 49534 6802
rect 49586 6750 50094 6802
rect 50146 6750 50148 6802
rect 49532 6748 50148 6750
rect 49532 6738 49588 6748
rect 50092 6738 50148 6748
rect 50428 6802 50484 6814
rect 50428 6750 50430 6802
rect 50482 6750 50484 6802
rect 50428 6692 50484 6750
rect 50428 6626 50484 6636
rect 50316 6580 50372 6590
rect 50316 6486 50372 6524
rect 50428 5908 50484 5918
rect 48748 5906 49252 5908
rect 48748 5854 48862 5906
rect 48914 5854 49252 5906
rect 48748 5852 49252 5854
rect 48860 5842 48916 5852
rect 48972 5684 49028 5694
rect 49196 5684 49252 5852
rect 49308 5906 49700 5908
rect 49308 5854 49310 5906
rect 49362 5854 49700 5906
rect 49308 5852 49700 5854
rect 49308 5842 49364 5852
rect 49196 5628 49476 5684
rect 48972 5348 49028 5628
rect 48972 5254 49028 5292
rect 49420 5346 49476 5628
rect 49420 5294 49422 5346
rect 49474 5294 49476 5346
rect 49420 5282 49476 5294
rect 48524 5070 48526 5122
rect 48578 5070 48580 5122
rect 48524 5058 48580 5070
rect 48748 5124 48804 5134
rect 49644 5124 49700 5852
rect 50428 5814 50484 5852
rect 49756 5796 49812 5806
rect 50092 5796 50148 5806
rect 49812 5794 50148 5796
rect 49812 5742 50094 5794
rect 50146 5742 50148 5794
rect 49812 5740 50148 5742
rect 49756 5702 49812 5740
rect 50092 5730 50148 5740
rect 50204 5794 50260 5806
rect 50204 5742 50206 5794
rect 50258 5742 50260 5794
rect 49756 5460 49812 5470
rect 49756 5346 49812 5404
rect 49756 5294 49758 5346
rect 49810 5294 49812 5346
rect 49756 5282 49812 5294
rect 49756 5124 49812 5134
rect 49644 5122 49812 5124
rect 49644 5070 49758 5122
rect 49810 5070 49812 5122
rect 49644 5068 49812 5070
rect 48748 5030 48804 5068
rect 49756 5058 49812 5068
rect 50204 5124 50260 5742
rect 50204 5058 50260 5068
rect 49084 5012 49140 5022
rect 49308 5012 49364 5022
rect 49084 5010 49308 5012
rect 49084 4958 49086 5010
rect 49138 4958 49308 5010
rect 49084 4956 49308 4958
rect 49084 4946 49140 4956
rect 49308 4946 49364 4956
rect 47964 3502 47966 3554
rect 48018 3502 48020 3554
rect 47964 3490 48020 3502
rect 50652 3332 50708 9772
rect 50988 9380 51044 9774
rect 50988 9314 51044 9324
rect 50988 9156 51044 9166
rect 50988 9062 51044 9100
rect 51100 8484 51156 9996
rect 51660 9828 51716 11118
rect 51660 9762 51716 9772
rect 51996 10498 52052 10510
rect 51996 10446 51998 10498
rect 52050 10446 52052 10498
rect 51884 9716 51940 9726
rect 51996 9716 52052 10446
rect 51940 9660 52052 9716
rect 51660 9042 51716 9054
rect 51660 8990 51662 9042
rect 51714 8990 51716 9042
rect 51286 8652 51550 8662
rect 51342 8596 51390 8652
rect 51446 8596 51494 8652
rect 51286 8586 51550 8596
rect 51660 8484 51716 8990
rect 51884 9042 51940 9660
rect 52332 9380 52388 9390
rect 52332 9154 52388 9324
rect 52332 9102 52334 9154
rect 52386 9102 52388 9154
rect 52332 9090 52388 9102
rect 51884 8990 51886 9042
rect 51938 8990 51940 9042
rect 51884 8978 51940 8990
rect 52108 8596 52164 8606
rect 52108 8484 52164 8540
rect 51100 8428 51492 8484
rect 51660 8428 52164 8484
rect 51436 8260 51492 8428
rect 51436 7362 51492 8204
rect 51772 7588 51828 7598
rect 51436 7310 51438 7362
rect 51490 7310 51492 7362
rect 51436 7298 51492 7310
rect 51548 7474 51604 7486
rect 51548 7422 51550 7474
rect 51602 7422 51604 7474
rect 51548 7364 51604 7422
rect 51548 7298 51604 7308
rect 50876 7250 50932 7262
rect 50876 7198 50878 7250
rect 50930 7198 50932 7250
rect 50876 6914 50932 7198
rect 51772 7140 51828 7532
rect 51286 7084 51550 7094
rect 51342 7028 51390 7084
rect 51446 7028 51494 7084
rect 51286 7018 51550 7028
rect 50876 6862 50878 6914
rect 50930 6862 50932 6914
rect 50876 6850 50932 6862
rect 51772 6690 51828 7084
rect 51772 6638 51774 6690
rect 51826 6638 51828 6690
rect 50876 6580 50932 6590
rect 50876 6486 50932 6524
rect 51324 6580 51380 6590
rect 51324 6486 51380 6524
rect 50988 6018 51044 6030
rect 50988 5966 50990 6018
rect 51042 5966 51044 6018
rect 50876 5794 50932 5806
rect 50876 5742 50878 5794
rect 50930 5742 50932 5794
rect 50764 5682 50820 5694
rect 50764 5630 50766 5682
rect 50818 5630 50820 5682
rect 50764 5236 50820 5630
rect 50764 5170 50820 5180
rect 50876 5012 50932 5742
rect 50988 5460 51044 5966
rect 51660 5796 51716 5806
rect 51772 5796 51828 6638
rect 51884 7028 51940 7038
rect 51884 6914 51940 6972
rect 51884 6862 51886 6914
rect 51938 6862 51940 6914
rect 51884 6018 51940 6862
rect 51884 5966 51886 6018
rect 51938 5966 51940 6018
rect 51884 5954 51940 5966
rect 51660 5794 51828 5796
rect 51660 5742 51662 5794
rect 51714 5742 51828 5794
rect 51660 5740 51828 5742
rect 51660 5730 51716 5740
rect 51286 5516 51550 5526
rect 51342 5460 51390 5516
rect 51446 5460 51494 5516
rect 51286 5450 51550 5460
rect 50988 5394 51044 5404
rect 51100 5348 51156 5358
rect 52108 5348 52164 8428
rect 52444 7700 52500 14140
rect 53004 13860 53060 13870
rect 53004 13766 53060 13804
rect 53340 13636 53396 13646
rect 53340 13542 53396 13580
rect 52556 9826 52612 9838
rect 52556 9774 52558 9826
rect 52610 9774 52612 9826
rect 52556 9716 52612 9774
rect 53116 9828 53172 9838
rect 53116 9734 53172 9772
rect 52556 9650 52612 9660
rect 53004 9714 53060 9726
rect 53004 9662 53006 9714
rect 53058 9662 53060 9714
rect 52892 9602 52948 9614
rect 52892 9550 52894 9602
rect 52946 9550 52948 9602
rect 52892 9156 52948 9550
rect 52892 8930 52948 9100
rect 52892 8878 52894 8930
rect 52946 8878 52948 8930
rect 52892 8866 52948 8878
rect 52892 8596 52948 8606
rect 53004 8596 53060 9662
rect 52948 8540 53060 8596
rect 53116 9044 53172 9054
rect 52892 8530 52948 8540
rect 52444 7634 52500 7644
rect 53004 8372 53060 8382
rect 53004 7474 53060 8316
rect 53004 7422 53006 7474
rect 53058 7422 53060 7474
rect 53004 7410 53060 7422
rect 53116 7250 53172 8988
rect 53116 7198 53118 7250
rect 53170 7198 53172 7250
rect 53116 7186 53172 7198
rect 53228 8372 53284 8382
rect 53452 8372 53508 15092
rect 53564 13748 53620 13758
rect 53676 13748 53732 16268
rect 53564 13746 53732 13748
rect 53564 13694 53566 13746
rect 53618 13694 53732 13746
rect 53564 13692 53732 13694
rect 53788 15090 53844 15102
rect 53788 15038 53790 15090
rect 53842 15038 53844 15090
rect 53564 12178 53620 13692
rect 53564 12126 53566 12178
rect 53618 12126 53620 12178
rect 53564 12114 53620 12126
rect 53788 10388 53844 15038
rect 53900 13972 53956 13982
rect 54012 13972 54068 21084
rect 54124 20804 54180 20814
rect 54124 20242 54180 20748
rect 54124 20190 54126 20242
rect 54178 20190 54180 20242
rect 54124 20178 54180 20190
rect 54236 19906 54292 21310
rect 54460 20692 54516 21646
rect 54460 20626 54516 20636
rect 54236 19854 54238 19906
rect 54290 19854 54292 19906
rect 54236 19842 54292 19854
rect 54684 18116 54740 24444
rect 54796 23042 54852 24892
rect 55244 24162 55300 26236
rect 55916 26402 55972 26414
rect 55916 26350 55918 26402
rect 55970 26350 55972 26402
rect 55916 26292 55972 26350
rect 55916 26226 55972 26236
rect 55692 26180 55748 26190
rect 55356 26124 55692 26180
rect 55356 24834 55412 26124
rect 55692 26086 55748 26124
rect 55804 26178 55860 26190
rect 55804 26126 55806 26178
rect 55858 26126 55860 26178
rect 55804 25508 55860 26126
rect 55804 25442 55860 25452
rect 55916 25620 55972 25630
rect 55916 25506 55972 25564
rect 56028 25618 56084 26852
rect 56028 25566 56030 25618
rect 56082 25566 56084 25618
rect 56028 25554 56084 25566
rect 56476 26516 56532 26526
rect 56476 25618 56532 26460
rect 56700 26180 56756 26190
rect 56700 26086 56756 26124
rect 56476 25566 56478 25618
rect 56530 25566 56532 25618
rect 56476 25554 56532 25566
rect 55916 25454 55918 25506
rect 55970 25454 55972 25506
rect 55916 25442 55972 25454
rect 55356 24782 55358 24834
rect 55410 24782 55412 24834
rect 55356 24770 55412 24782
rect 56140 25394 56196 25406
rect 56140 25342 56142 25394
rect 56194 25342 56196 25394
rect 56140 24836 56196 25342
rect 56588 24836 56644 24846
rect 56140 24834 56644 24836
rect 56140 24782 56590 24834
rect 56642 24782 56644 24834
rect 56140 24780 56644 24782
rect 56588 24770 56644 24780
rect 56028 24722 56084 24734
rect 56028 24670 56030 24722
rect 56082 24670 56084 24722
rect 55804 24610 55860 24622
rect 55804 24558 55806 24610
rect 55858 24558 55860 24610
rect 55692 24500 55748 24510
rect 55244 24110 55246 24162
rect 55298 24110 55300 24162
rect 55244 24098 55300 24110
rect 55468 24498 55748 24500
rect 55468 24446 55694 24498
rect 55746 24446 55748 24498
rect 55468 24444 55748 24446
rect 55356 23714 55412 23726
rect 55356 23662 55358 23714
rect 55410 23662 55412 23714
rect 55020 23266 55076 23278
rect 55020 23214 55022 23266
rect 55074 23214 55076 23266
rect 54796 22990 54798 23042
rect 54850 22990 54852 23042
rect 54796 22978 54852 22990
rect 54908 23154 54964 23166
rect 54908 23102 54910 23154
rect 54962 23102 54964 23154
rect 54908 23044 54964 23102
rect 54908 22978 54964 22988
rect 55020 22932 55076 23214
rect 55020 22866 55076 22876
rect 55020 22596 55076 22606
rect 55020 22502 55076 22540
rect 55356 22484 55412 23662
rect 55468 22708 55524 24444
rect 55692 24434 55748 24444
rect 55580 24164 55636 24174
rect 55804 24164 55860 24558
rect 55580 24162 55860 24164
rect 55580 24110 55582 24162
rect 55634 24110 55860 24162
rect 55580 24108 55860 24110
rect 55580 24098 55636 24108
rect 55468 22642 55524 22652
rect 56028 23156 56084 24670
rect 56812 24722 56868 26908
rect 56812 24670 56814 24722
rect 56866 24670 56868 24722
rect 56812 23938 56868 24670
rect 56812 23886 56814 23938
rect 56866 23886 56868 23938
rect 56812 23874 56868 23886
rect 57036 24722 57092 27806
rect 57148 27746 57204 27758
rect 57148 27694 57150 27746
rect 57202 27694 57204 27746
rect 57148 27298 57204 27694
rect 57148 27246 57150 27298
rect 57202 27246 57204 27298
rect 57148 27234 57204 27246
rect 57260 27076 57316 27086
rect 57260 26982 57316 27020
rect 57372 26852 57428 28476
rect 57596 27748 57652 29708
rect 57708 29426 57764 29934
rect 57708 29374 57710 29426
rect 57762 29374 57764 29426
rect 57708 29362 57764 29374
rect 57932 29540 57988 30158
rect 57820 28868 57876 28878
rect 57820 27970 57876 28812
rect 57820 27918 57822 27970
rect 57874 27918 57876 27970
rect 57708 27748 57764 27758
rect 57596 27746 57764 27748
rect 57596 27694 57710 27746
rect 57762 27694 57764 27746
rect 57596 27692 57764 27694
rect 57708 27682 57764 27692
rect 57484 27300 57540 27310
rect 57484 27074 57540 27244
rect 57484 27022 57486 27074
rect 57538 27022 57540 27074
rect 57484 27010 57540 27022
rect 57372 26786 57428 26796
rect 57036 24670 57038 24722
rect 57090 24670 57092 24722
rect 56028 22596 56084 23100
rect 56252 23828 56308 23838
rect 56140 22596 56196 22606
rect 56028 22594 56196 22596
rect 56028 22542 56142 22594
rect 56194 22542 56196 22594
rect 56028 22540 56196 22542
rect 56140 22530 56196 22540
rect 55356 22428 55636 22484
rect 55244 21588 55300 21598
rect 54796 20690 54852 20702
rect 54796 20638 54798 20690
rect 54850 20638 54852 20690
rect 54796 20468 54852 20638
rect 54796 20402 54852 20412
rect 55244 20020 55300 21532
rect 55580 21474 55636 22428
rect 55916 22482 55972 22494
rect 55916 22430 55918 22482
rect 55970 22430 55972 22482
rect 55804 22372 55860 22382
rect 55692 22370 55860 22372
rect 55692 22318 55806 22370
rect 55858 22318 55860 22370
rect 55692 22316 55860 22318
rect 55692 21812 55748 22316
rect 55804 22306 55860 22316
rect 55692 21718 55748 21756
rect 55916 21700 55972 22430
rect 55916 21606 55972 21644
rect 55580 21422 55582 21474
rect 55634 21422 55636 21474
rect 55580 21410 55636 21422
rect 55804 20804 55860 20814
rect 55468 20802 55860 20804
rect 55468 20750 55806 20802
rect 55858 20750 55860 20802
rect 55468 20748 55860 20750
rect 55356 20690 55412 20702
rect 55356 20638 55358 20690
rect 55410 20638 55412 20690
rect 55356 20188 55412 20638
rect 55468 20690 55524 20748
rect 55804 20738 55860 20748
rect 55468 20638 55470 20690
rect 55522 20638 55524 20690
rect 55468 20626 55524 20638
rect 56140 20690 56196 20702
rect 56140 20638 56142 20690
rect 56194 20638 56196 20690
rect 55692 20580 55748 20590
rect 56028 20580 56084 20590
rect 55692 20486 55748 20524
rect 55804 20578 56084 20580
rect 55804 20526 56030 20578
rect 56082 20526 56084 20578
rect 55804 20524 56084 20526
rect 55356 20132 55748 20188
rect 55692 20130 55748 20132
rect 55692 20078 55694 20130
rect 55746 20078 55748 20130
rect 55692 20066 55748 20078
rect 55804 20132 55860 20524
rect 56028 20514 56084 20524
rect 56140 20468 56196 20638
rect 56140 20402 56196 20412
rect 55804 20066 55860 20076
rect 55916 20130 55972 20142
rect 55916 20078 55918 20130
rect 55970 20078 55972 20130
rect 55244 19964 55412 20020
rect 55020 19346 55076 19358
rect 55020 19294 55022 19346
rect 55074 19294 55076 19346
rect 55020 19236 55076 19294
rect 55020 19170 55076 19180
rect 55132 19234 55188 19246
rect 55132 19182 55134 19234
rect 55186 19182 55188 19234
rect 54796 19122 54852 19134
rect 54796 19070 54798 19122
rect 54850 19070 54852 19122
rect 54796 18340 54852 19070
rect 55132 18452 55188 19182
rect 55132 18358 55188 18396
rect 54796 18274 54852 18284
rect 54684 18060 54852 18116
rect 54460 17780 54516 17790
rect 54460 17666 54516 17724
rect 54460 17614 54462 17666
rect 54514 17614 54516 17666
rect 54460 17602 54516 17614
rect 54684 17556 54740 17566
rect 54348 16884 54404 16894
rect 54348 16770 54404 16828
rect 54684 16882 54740 17500
rect 54684 16830 54686 16882
rect 54738 16830 54740 16882
rect 54684 16818 54740 16830
rect 54348 16718 54350 16770
rect 54402 16718 54404 16770
rect 54348 16706 54404 16718
rect 54796 16660 54852 18060
rect 55244 17780 55300 17790
rect 55244 17686 55300 17724
rect 54908 17666 54964 17678
rect 54908 17614 54910 17666
rect 54962 17614 54964 17666
rect 54908 16884 54964 17614
rect 54908 16818 54964 16828
rect 55132 16884 55188 16894
rect 55132 16790 55188 16828
rect 54796 16604 54964 16660
rect 54796 15314 54852 15326
rect 54796 15262 54798 15314
rect 54850 15262 54852 15314
rect 54796 15204 54852 15262
rect 54796 15138 54852 15148
rect 53900 13970 54068 13972
rect 53900 13918 53902 13970
rect 53954 13918 54068 13970
rect 53900 13916 54068 13918
rect 54684 15090 54740 15102
rect 54684 15038 54686 15090
rect 54738 15038 54740 15090
rect 54684 14418 54740 15038
rect 54908 14644 54964 16604
rect 55244 15986 55300 15998
rect 55244 15934 55246 15986
rect 55298 15934 55300 15986
rect 55132 15428 55188 15438
rect 55132 15202 55188 15372
rect 55132 15150 55134 15202
rect 55186 15150 55188 15202
rect 55132 15138 55188 15150
rect 55020 14756 55076 14766
rect 55244 14756 55300 15934
rect 55020 14754 55300 14756
rect 55020 14702 55022 14754
rect 55074 14702 55300 14754
rect 55020 14700 55300 14702
rect 55020 14690 55076 14700
rect 54908 14578 54964 14588
rect 54684 14366 54686 14418
rect 54738 14366 54740 14418
rect 53900 13906 53956 13916
rect 54684 13634 54740 14366
rect 54908 14306 54964 14318
rect 54908 14254 54910 14306
rect 54962 14254 54964 14306
rect 54908 13860 54964 14254
rect 55356 13972 55412 19964
rect 55916 19460 55972 20078
rect 56028 20018 56084 20030
rect 56028 19966 56030 20018
rect 56082 19966 56084 20018
rect 56028 19908 56084 19966
rect 56028 19842 56084 19852
rect 55916 19394 55972 19404
rect 56252 19346 56308 23772
rect 57036 23828 57092 24670
rect 57036 23762 57092 23772
rect 57148 26292 57204 26302
rect 56252 19294 56254 19346
rect 56306 19294 56308 19346
rect 56252 19282 56308 19294
rect 56476 23716 56532 23726
rect 55468 19234 55524 19246
rect 55468 19182 55470 19234
rect 55522 19182 55524 19234
rect 55468 17892 55524 19182
rect 55692 19236 55748 19246
rect 55692 19142 55748 19180
rect 56028 18450 56084 18462
rect 56028 18398 56030 18450
rect 56082 18398 56084 18450
rect 55580 18340 55636 18350
rect 55580 18246 55636 18284
rect 56028 18340 56084 18398
rect 55580 17892 55636 17902
rect 55468 17890 55636 17892
rect 55468 17838 55582 17890
rect 55634 17838 55636 17890
rect 55468 17836 55636 17838
rect 55580 17826 55636 17836
rect 55692 17892 55748 17902
rect 55916 17892 55972 17902
rect 56028 17892 56084 18284
rect 55748 17836 55860 17892
rect 55692 17826 55748 17836
rect 55580 17668 55636 17678
rect 55580 17444 55636 17612
rect 55580 17378 55636 17388
rect 55804 17108 55860 17836
rect 55916 17890 56084 17892
rect 55916 17838 55918 17890
rect 55970 17838 56084 17890
rect 55916 17836 56084 17838
rect 55916 17826 55972 17836
rect 56252 17556 56308 17566
rect 56140 17554 56308 17556
rect 56140 17502 56254 17554
rect 56306 17502 56308 17554
rect 56140 17500 56308 17502
rect 56028 17444 56084 17454
rect 55916 17108 55972 17118
rect 55804 17052 55916 17108
rect 55916 17014 55972 17052
rect 55692 16884 55748 16894
rect 55692 16770 55748 16828
rect 55692 16718 55694 16770
rect 55746 16718 55748 16770
rect 55692 16706 55748 16718
rect 56028 16770 56084 17388
rect 56028 16718 56030 16770
rect 56082 16718 56084 16770
rect 56028 16706 56084 16718
rect 55580 16324 55636 16334
rect 55580 16322 56084 16324
rect 55580 16270 55582 16322
rect 55634 16270 56084 16322
rect 55580 16268 56084 16270
rect 55580 16258 55636 16268
rect 55580 16100 55636 16110
rect 55580 16098 55748 16100
rect 55580 16046 55582 16098
rect 55634 16046 55748 16098
rect 55580 16044 55748 16046
rect 55580 16034 55636 16044
rect 55692 15202 55748 16044
rect 55916 15540 55972 16268
rect 56028 16210 56084 16268
rect 56028 16158 56030 16210
rect 56082 16158 56084 16210
rect 56028 16146 56084 16158
rect 55692 15150 55694 15202
rect 55746 15150 55748 15202
rect 55692 15138 55748 15150
rect 55804 15426 55860 15438
rect 55804 15374 55806 15426
rect 55858 15374 55860 15426
rect 55804 15204 55860 15374
rect 55804 15138 55860 15148
rect 55916 14756 55972 15484
rect 56028 15428 56084 15438
rect 56140 15428 56196 17500
rect 56252 17490 56308 17500
rect 56084 15372 56196 15428
rect 56252 15986 56308 15998
rect 56252 15934 56254 15986
rect 56306 15934 56308 15986
rect 56028 15334 56084 15372
rect 56140 15204 56196 15214
rect 55692 14700 55972 14756
rect 56028 15092 56196 15148
rect 55692 14196 55748 14700
rect 55804 14532 55860 14542
rect 55804 14438 55860 14476
rect 55692 14140 55972 14196
rect 54908 13746 54964 13804
rect 54908 13694 54910 13746
rect 54962 13694 54964 13746
rect 54908 13682 54964 13694
rect 55244 13916 55412 13972
rect 55916 13970 55972 14140
rect 55916 13918 55918 13970
rect 55970 13918 55972 13970
rect 54684 13582 54686 13634
rect 54738 13582 54740 13634
rect 54684 13570 54740 13582
rect 55244 12292 55300 13916
rect 55916 13906 55972 13918
rect 56028 13858 56084 15092
rect 56140 14644 56196 14682
rect 56140 14578 56196 14588
rect 56252 14532 56308 15934
rect 56252 14466 56308 14476
rect 56028 13806 56030 13858
rect 56082 13806 56084 13858
rect 56028 13794 56084 13806
rect 56140 14418 56196 14430
rect 56140 14366 56142 14418
rect 56194 14366 56196 14418
rect 55244 12226 55300 12236
rect 55356 13746 55412 13758
rect 55356 13694 55358 13746
rect 55410 13694 55412 13746
rect 55356 12404 55412 13694
rect 55916 13524 55972 13534
rect 56140 13524 56196 14366
rect 55916 13522 56196 13524
rect 55916 13470 55918 13522
rect 55970 13470 56196 13522
rect 55916 13468 56196 13470
rect 55916 13458 55972 13468
rect 55468 13076 55524 13086
rect 55468 12982 55524 13020
rect 55468 12404 55524 12414
rect 55356 12402 55524 12404
rect 55356 12350 55470 12402
rect 55522 12350 55524 12402
rect 55356 12348 55524 12350
rect 54908 11956 54964 11966
rect 55244 11956 55300 11966
rect 54908 11862 54964 11900
rect 55132 11954 55300 11956
rect 55132 11902 55246 11954
rect 55298 11902 55300 11954
rect 55132 11900 55300 11902
rect 54796 11396 54852 11406
rect 55132 11396 55188 11900
rect 55244 11890 55300 11900
rect 54796 11394 55188 11396
rect 54796 11342 54798 11394
rect 54850 11342 55188 11394
rect 54796 11340 55188 11342
rect 55244 11396 55300 11406
rect 55356 11396 55412 12348
rect 55468 12338 55524 12348
rect 56140 12292 56196 12302
rect 55580 12068 55636 12078
rect 55580 11974 55636 12012
rect 55244 11394 55412 11396
rect 55244 11342 55246 11394
rect 55298 11342 55412 11394
rect 55244 11340 55412 11342
rect 56140 11844 56196 12236
rect 54572 11282 54628 11294
rect 54572 11230 54574 11282
rect 54626 11230 54628 11282
rect 53900 10836 53956 10846
rect 53900 10742 53956 10780
rect 54460 10612 54516 10622
rect 54572 10612 54628 11230
rect 54460 10610 54628 10612
rect 54460 10558 54462 10610
rect 54514 10558 54628 10610
rect 54460 10556 54628 10558
rect 53788 10332 54404 10388
rect 53900 10164 53956 10174
rect 53900 9266 53956 10108
rect 53900 9214 53902 9266
rect 53954 9214 53956 9266
rect 53900 9202 53956 9214
rect 53788 9156 53844 9166
rect 53788 9062 53844 9100
rect 54012 9154 54068 9166
rect 54012 9102 54014 9154
rect 54066 9102 54068 9154
rect 54012 9044 54068 9102
rect 54012 8978 54068 8988
rect 54348 9156 54404 10332
rect 54460 9828 54516 10556
rect 54460 9762 54516 9772
rect 54796 9716 54852 11340
rect 55244 11330 55300 11340
rect 56140 11282 56196 11788
rect 56140 11230 56142 11282
rect 56194 11230 56196 11282
rect 56140 11218 56196 11230
rect 56252 11170 56308 11182
rect 56252 11118 56254 11170
rect 56306 11118 56308 11170
rect 55356 10724 55412 10734
rect 54908 10722 55412 10724
rect 54908 10670 55358 10722
rect 55410 10670 55412 10722
rect 54908 10668 55412 10670
rect 54908 10164 54964 10668
rect 54908 9938 54964 10108
rect 54908 9886 54910 9938
rect 54962 9886 54964 9938
rect 54908 9874 54964 9886
rect 55132 9828 55188 9838
rect 54796 9660 55076 9716
rect 54796 9156 54852 9166
rect 54348 9154 54852 9156
rect 54348 9102 54798 9154
rect 54850 9102 54852 9154
rect 54348 9100 54852 9102
rect 53228 8370 53508 8372
rect 53228 8318 53230 8370
rect 53282 8318 53508 8370
rect 53228 8316 53508 8318
rect 54348 8482 54404 9100
rect 54796 9090 54852 9100
rect 54908 9154 54964 9166
rect 54908 9102 54910 9154
rect 54962 9102 54964 9154
rect 54908 9044 54964 9102
rect 54908 8978 54964 8988
rect 54348 8430 54350 8482
rect 54402 8430 54404 8482
rect 54348 8372 54404 8430
rect 53228 6804 53284 8316
rect 54348 8306 54404 8316
rect 54572 8932 54628 8942
rect 54572 8260 54628 8876
rect 54908 8818 54964 8830
rect 54908 8766 54910 8818
rect 54962 8766 54964 8818
rect 54684 8372 54740 8382
rect 54684 8278 54740 8316
rect 54572 8146 54628 8204
rect 54908 8258 54964 8766
rect 55020 8372 55076 9660
rect 55132 8820 55188 9772
rect 55356 9042 55412 10668
rect 55916 10498 55972 10510
rect 55916 10446 55918 10498
rect 55970 10446 55972 10498
rect 55916 10052 55972 10446
rect 55916 9986 55972 9996
rect 55804 9826 55860 9838
rect 55804 9774 55806 9826
rect 55858 9774 55860 9826
rect 55356 8990 55358 9042
rect 55410 8990 55412 9042
rect 55356 8978 55412 8990
rect 55468 9602 55524 9614
rect 55468 9550 55470 9602
rect 55522 9550 55524 9602
rect 55468 9044 55524 9550
rect 55692 9044 55748 9054
rect 55468 8988 55692 9044
rect 55692 8978 55748 8988
rect 55580 8820 55636 8830
rect 55132 8818 55636 8820
rect 55132 8766 55582 8818
rect 55634 8766 55636 8818
rect 55132 8764 55636 8766
rect 55580 8754 55636 8764
rect 55356 8484 55412 8494
rect 55804 8484 55860 9774
rect 55916 8820 55972 8830
rect 55916 8726 55972 8764
rect 55916 8484 55972 8494
rect 55804 8482 55972 8484
rect 55804 8430 55918 8482
rect 55970 8430 55972 8482
rect 55804 8428 55972 8430
rect 55132 8372 55188 8382
rect 55020 8370 55188 8372
rect 55020 8318 55134 8370
rect 55186 8318 55188 8370
rect 55020 8316 55188 8318
rect 55132 8306 55188 8316
rect 54908 8206 54910 8258
rect 54962 8206 54964 8258
rect 54908 8194 54964 8206
rect 55244 8258 55300 8270
rect 55244 8206 55246 8258
rect 55298 8206 55300 8258
rect 54572 8094 54574 8146
rect 54626 8094 54628 8146
rect 54572 8082 54628 8094
rect 53340 8036 53396 8046
rect 53340 7942 53396 7980
rect 53452 8034 53508 8046
rect 53452 7982 53454 8034
rect 53506 7982 53508 8034
rect 53452 7028 53508 7982
rect 54124 8034 54180 8046
rect 54124 7982 54126 8034
rect 54178 7982 54180 8034
rect 54124 7588 54180 7982
rect 54124 7494 54180 7532
rect 54908 8036 54964 8046
rect 54348 7474 54404 7486
rect 54348 7422 54350 7474
rect 54402 7422 54404 7474
rect 53508 6972 53732 7028
rect 53452 6962 53508 6972
rect 53676 6804 53732 6972
rect 54012 6804 54068 6814
rect 53676 6748 53844 6804
rect 53004 6692 53060 6702
rect 53004 6598 53060 6636
rect 53228 5906 53284 6748
rect 53564 6690 53620 6702
rect 53564 6638 53566 6690
rect 53618 6638 53620 6690
rect 53228 5854 53230 5906
rect 53282 5854 53284 5906
rect 53228 5842 53284 5854
rect 53452 6580 53508 6590
rect 51100 5346 51828 5348
rect 51100 5294 51102 5346
rect 51154 5294 51828 5346
rect 51100 5292 51828 5294
rect 51100 5282 51156 5292
rect 51436 5124 51492 5134
rect 51436 5030 51492 5068
rect 51660 5124 51716 5134
rect 51660 5030 51716 5068
rect 51772 5122 51828 5292
rect 52108 5282 52164 5292
rect 53116 5348 53172 5358
rect 51772 5070 51774 5122
rect 51826 5070 51828 5122
rect 51772 5058 51828 5070
rect 51996 5122 52052 5134
rect 51996 5070 51998 5122
rect 52050 5070 52052 5122
rect 51100 5012 51156 5022
rect 50876 5010 51156 5012
rect 50876 4958 51102 5010
rect 51154 4958 51156 5010
rect 50876 4956 51156 4958
rect 51100 4452 51156 4956
rect 51212 5012 51268 5022
rect 51212 4918 51268 4956
rect 51996 4676 52052 5070
rect 53116 5122 53172 5292
rect 53452 5234 53508 6524
rect 53564 6132 53620 6638
rect 53676 6580 53732 6590
rect 53676 6486 53732 6524
rect 53788 6356 53844 6748
rect 54012 6690 54068 6748
rect 54012 6638 54014 6690
rect 54066 6638 54068 6690
rect 54012 6626 54068 6638
rect 54124 6692 54180 6702
rect 54180 6636 54292 6692
rect 54124 6626 54180 6636
rect 54124 6466 54180 6478
rect 54124 6414 54126 6466
rect 54178 6414 54180 6466
rect 54124 6356 54180 6414
rect 53788 6300 54180 6356
rect 54124 6132 54180 6142
rect 54236 6132 54292 6636
rect 54348 6690 54404 7422
rect 54908 7474 54964 7980
rect 55020 7700 55076 7710
rect 55020 7606 55076 7644
rect 54908 7422 54910 7474
rect 54962 7422 54964 7474
rect 54908 7410 54964 7422
rect 55244 7364 55300 8206
rect 55244 7298 55300 7308
rect 54348 6638 54350 6690
rect 54402 6638 54404 6690
rect 54348 6626 54404 6638
rect 53564 6130 54068 6132
rect 53564 6078 53566 6130
rect 53618 6078 54068 6130
rect 53564 6076 54068 6078
rect 53564 6066 53620 6076
rect 54012 6018 54068 6076
rect 54124 6130 54292 6132
rect 54124 6078 54126 6130
rect 54178 6078 54292 6130
rect 54124 6076 54292 6078
rect 54796 6580 54852 6590
rect 54124 6066 54180 6076
rect 54012 5966 54014 6018
rect 54066 5966 54068 6018
rect 54012 5954 54068 5966
rect 54684 6018 54740 6030
rect 54684 5966 54686 6018
rect 54738 5966 54740 6018
rect 54460 5906 54516 5918
rect 54460 5854 54462 5906
rect 54514 5854 54516 5906
rect 54124 5684 54180 5694
rect 54124 5682 54292 5684
rect 54124 5630 54126 5682
rect 54178 5630 54292 5682
rect 54124 5628 54292 5630
rect 54124 5618 54180 5628
rect 53452 5182 53454 5234
rect 53506 5182 53508 5234
rect 53452 5170 53508 5182
rect 53116 5070 53118 5122
rect 53170 5070 53172 5122
rect 53116 5058 53172 5070
rect 54012 5124 54068 5134
rect 54012 5030 54068 5068
rect 51100 4386 51156 4396
rect 51884 4620 52052 4676
rect 52220 5012 52276 5022
rect 52668 5012 52724 5022
rect 52276 5010 52724 5012
rect 52276 4958 52670 5010
rect 52722 4958 52724 5010
rect 52276 4956 52724 4958
rect 51884 4226 51940 4620
rect 51996 4452 52052 4462
rect 51996 4358 52052 4396
rect 52220 4450 52276 4956
rect 52668 4946 52724 4956
rect 54236 5010 54292 5628
rect 54348 5124 54404 5134
rect 54460 5124 54516 5854
rect 54684 5348 54740 5966
rect 54796 6018 54852 6524
rect 54796 5966 54798 6018
rect 54850 5966 54852 6018
rect 54796 5954 54852 5966
rect 54684 5282 54740 5292
rect 55244 5348 55300 5358
rect 55356 5348 55412 8428
rect 55916 8418 55972 8428
rect 55468 8372 55524 8382
rect 55468 8258 55524 8316
rect 56252 8372 56308 11118
rect 56476 9940 56532 23660
rect 57148 23380 57204 26236
rect 57596 26178 57652 26190
rect 57596 26126 57598 26178
rect 57650 26126 57652 26178
rect 57596 25620 57652 26126
rect 57260 25506 57316 25518
rect 57260 25454 57262 25506
rect 57314 25454 57316 25506
rect 57260 24612 57316 25454
rect 57260 23716 57316 24556
rect 57596 23938 57652 25564
rect 57708 25508 57764 25518
rect 57820 25508 57876 27918
rect 57708 25506 57876 25508
rect 57708 25454 57710 25506
rect 57762 25454 57876 25506
rect 57708 25452 57876 25454
rect 57932 28754 57988 29484
rect 57932 28702 57934 28754
rect 57986 28702 57988 28754
rect 57708 25442 57764 25452
rect 57932 24276 57988 28702
rect 58044 27634 58100 30828
rect 58156 29314 58212 29326
rect 58156 29262 58158 29314
rect 58210 29262 58212 29314
rect 58156 28532 58212 29262
rect 58156 28466 58212 28476
rect 58044 27582 58046 27634
rect 58098 27582 58100 27634
rect 58044 26178 58100 27582
rect 58044 26126 58046 26178
rect 58098 26126 58100 26178
rect 58044 24612 58100 26126
rect 58156 24612 58212 24622
rect 58044 24556 58156 24612
rect 58156 24518 58212 24556
rect 57932 24220 58100 24276
rect 57596 23886 57598 23938
rect 57650 23886 57652 23938
rect 57596 23874 57652 23886
rect 57260 23650 57316 23660
rect 57148 23324 57428 23380
rect 56924 23156 56980 23166
rect 56924 23062 56980 23100
rect 56700 23042 56756 23054
rect 56700 22990 56702 23042
rect 56754 22990 56756 23042
rect 56700 22596 56756 22990
rect 56700 22530 56756 22540
rect 57036 22372 57092 22382
rect 56812 22370 57092 22372
rect 56812 22318 57038 22370
rect 57090 22318 57092 22370
rect 56812 22316 57092 22318
rect 56812 20804 56868 22316
rect 57036 22306 57092 22316
rect 57260 22372 57316 22382
rect 57260 22036 57316 22316
rect 57036 21980 57316 22036
rect 57036 20914 57092 21980
rect 57372 21924 57428 23324
rect 57596 23042 57652 23054
rect 57596 22990 57598 23042
rect 57650 22990 57652 23042
rect 57596 22372 57652 22990
rect 57596 22306 57652 22316
rect 57596 22148 57652 22158
rect 57596 22146 57876 22148
rect 57596 22094 57598 22146
rect 57650 22094 57876 22146
rect 57596 22092 57876 22094
rect 57596 22082 57652 22092
rect 57372 21868 57764 21924
rect 57036 20862 57038 20914
rect 57090 20862 57092 20914
rect 57036 20850 57092 20862
rect 57260 21698 57316 21710
rect 57260 21646 57262 21698
rect 57314 21646 57316 21698
rect 56924 20804 56980 20814
rect 56812 20802 56980 20804
rect 56812 20750 56926 20802
rect 56978 20750 56980 20802
rect 56812 20748 56980 20750
rect 56812 20580 56868 20748
rect 56924 20738 56980 20748
rect 56812 20514 56868 20524
rect 56700 20468 56756 20478
rect 56700 20018 56756 20412
rect 56700 19966 56702 20018
rect 56754 19966 56756 20018
rect 56700 19954 56756 19966
rect 57036 20132 57092 20142
rect 57036 20018 57092 20076
rect 57036 19966 57038 20018
rect 57090 19966 57092 20018
rect 57036 19954 57092 19966
rect 56588 19908 56644 19918
rect 56588 19684 56644 19852
rect 56588 19628 56980 19684
rect 56812 19460 56868 19470
rect 56812 19234 56868 19404
rect 56924 19346 56980 19628
rect 56924 19294 56926 19346
rect 56978 19294 56980 19346
rect 56924 19282 56980 19294
rect 56812 19182 56814 19234
rect 56866 19182 56868 19234
rect 56812 19170 56868 19182
rect 57148 18450 57204 18462
rect 57148 18398 57150 18450
rect 57202 18398 57204 18450
rect 56812 18340 56868 18350
rect 56812 18246 56868 18284
rect 56700 18226 56756 18238
rect 56700 18174 56702 18226
rect 56754 18174 56756 18226
rect 56700 17778 56756 18174
rect 56700 17726 56702 17778
rect 56754 17726 56756 17778
rect 56700 15426 56756 17726
rect 56924 17666 56980 17678
rect 56924 17614 56926 17666
rect 56978 17614 56980 17666
rect 56812 16884 56868 16894
rect 56812 16790 56868 16828
rect 56924 16658 56980 17614
rect 57148 17668 57204 18398
rect 57148 17602 57204 17612
rect 56924 16606 56926 16658
rect 56978 16606 56980 16658
rect 56924 15538 56980 16606
rect 56924 15486 56926 15538
rect 56978 15486 56980 15538
rect 56924 15474 56980 15486
rect 57036 17556 57092 17566
rect 56700 15374 56702 15426
rect 56754 15374 56756 15426
rect 56700 15362 56756 15374
rect 57036 15202 57092 17500
rect 57148 17108 57204 17118
rect 57148 16882 57204 17052
rect 57148 16830 57150 16882
rect 57202 16830 57204 16882
rect 57148 16818 57204 16830
rect 57036 15150 57038 15202
rect 57090 15150 57092 15202
rect 57036 15138 57092 15150
rect 57260 14420 57316 21646
rect 57372 21588 57428 21598
rect 57372 21494 57428 21532
rect 57484 19460 57540 19470
rect 57372 19458 57540 19460
rect 57372 19406 57486 19458
rect 57538 19406 57540 19458
rect 57372 19404 57540 19406
rect 57372 15148 57428 19404
rect 57484 19394 57540 19404
rect 57708 17780 57764 21868
rect 57820 21586 57876 22092
rect 57932 21812 57988 21822
rect 58044 21812 58100 24220
rect 57932 21810 58100 21812
rect 57932 21758 57934 21810
rect 57986 21758 58100 21810
rect 57932 21756 58100 21758
rect 58156 23826 58212 23838
rect 58156 23774 58158 23826
rect 58210 23774 58212 23826
rect 57932 21746 57988 21756
rect 57820 21534 57822 21586
rect 57874 21534 57876 21586
rect 57820 21522 57876 21534
rect 58044 21588 58100 21598
rect 58044 20914 58100 21532
rect 58044 20862 58046 20914
rect 58098 20862 58100 20914
rect 58044 20850 58100 20862
rect 57820 17780 57876 17790
rect 57708 17778 57876 17780
rect 57708 17726 57822 17778
rect 57874 17726 57876 17778
rect 57708 17724 57876 17726
rect 57820 17714 57876 17724
rect 57708 17556 57764 17566
rect 57708 17462 57764 17500
rect 57932 17444 57988 17454
rect 57932 17350 57988 17388
rect 58156 17220 58212 23774
rect 57932 17164 58212 17220
rect 57932 16100 57988 17164
rect 57708 16044 57988 16100
rect 57484 15540 57540 15550
rect 57484 15446 57540 15484
rect 57708 15426 57764 16044
rect 57932 15986 57988 16044
rect 57932 15934 57934 15986
rect 57986 15934 57988 15986
rect 57932 15922 57988 15934
rect 57708 15374 57710 15426
rect 57762 15374 57764 15426
rect 57596 15202 57652 15214
rect 57596 15150 57598 15202
rect 57650 15150 57652 15202
rect 57372 15092 57540 15148
rect 57260 14364 57428 14420
rect 57260 14196 57316 14206
rect 57148 14140 57260 14196
rect 56700 13746 56756 13758
rect 56700 13694 56702 13746
rect 56754 13694 56756 13746
rect 56588 12962 56644 12974
rect 56588 12910 56590 12962
rect 56642 12910 56644 12962
rect 56588 12292 56644 12910
rect 56700 12402 56756 13694
rect 56700 12350 56702 12402
rect 56754 12350 56756 12402
rect 56700 12338 56756 12350
rect 56588 12198 56644 12236
rect 56812 12290 56868 12302
rect 56812 12238 56814 12290
rect 56866 12238 56868 12290
rect 56812 12068 56868 12238
rect 57148 12292 57204 14140
rect 57260 14130 57316 14140
rect 57372 13860 57428 14364
rect 57484 13972 57540 15092
rect 57596 14530 57652 15150
rect 57708 15204 57764 15374
rect 57708 15138 57764 15148
rect 57820 15874 57876 15886
rect 57820 15822 57822 15874
rect 57874 15822 57876 15874
rect 57596 14478 57598 14530
rect 57650 14478 57652 14530
rect 57596 14466 57652 14478
rect 57820 14196 57876 15822
rect 57820 14130 57876 14140
rect 57484 13916 57764 13972
rect 57372 13804 57540 13860
rect 57260 13746 57316 13758
rect 57260 13694 57262 13746
rect 57314 13694 57316 13746
rect 57260 13300 57316 13694
rect 57372 13300 57428 13310
rect 57260 13244 57372 13300
rect 57372 13234 57428 13244
rect 57484 13188 57540 13804
rect 57484 13122 57540 13132
rect 57596 13746 57652 13758
rect 57596 13694 57598 13746
rect 57650 13694 57652 13746
rect 57372 12850 57428 12862
rect 57372 12798 57374 12850
rect 57426 12798 57428 12850
rect 57260 12292 57316 12302
rect 57204 12290 57316 12292
rect 57204 12238 57262 12290
rect 57314 12238 57316 12290
rect 57204 12236 57316 12238
rect 57148 12198 57204 12236
rect 57260 12226 57316 12236
rect 57372 12290 57428 12798
rect 57596 12402 57652 13694
rect 57596 12350 57598 12402
rect 57650 12350 57652 12402
rect 57596 12338 57652 12350
rect 57372 12238 57374 12290
rect 57426 12238 57428 12290
rect 56812 12002 56868 12012
rect 57372 12068 57428 12238
rect 57372 12002 57428 12012
rect 56812 11844 56868 11854
rect 56812 10498 56868 11788
rect 57148 11844 57204 11854
rect 57148 10610 57204 11788
rect 57148 10558 57150 10610
rect 57202 10558 57204 10610
rect 57148 10546 57204 10558
rect 57484 11282 57540 11294
rect 57484 11230 57486 11282
rect 57538 11230 57540 11282
rect 56812 10446 56814 10498
rect 56866 10446 56868 10498
rect 56812 10434 56868 10446
rect 57484 10388 57540 11230
rect 57708 10612 57764 13916
rect 57820 13636 57876 13646
rect 58268 13636 58324 32620
rect 58439 31388 58703 31398
rect 58495 31332 58543 31388
rect 58599 31332 58647 31388
rect 58439 31322 58703 31332
rect 58439 29820 58703 29830
rect 58495 29764 58543 29820
rect 58599 29764 58647 29820
rect 58439 29754 58703 29764
rect 58439 28252 58703 28262
rect 58495 28196 58543 28252
rect 58599 28196 58647 28252
rect 58439 28186 58703 28196
rect 58439 26684 58703 26694
rect 58495 26628 58543 26684
rect 58599 26628 58647 26684
rect 58439 26618 58703 26628
rect 58439 25116 58703 25126
rect 58495 25060 58543 25116
rect 58599 25060 58647 25116
rect 58439 25050 58703 25060
rect 58439 23548 58703 23558
rect 58495 23492 58543 23548
rect 58599 23492 58647 23548
rect 58439 23482 58703 23492
rect 58439 21980 58703 21990
rect 58495 21924 58543 21980
rect 58599 21924 58647 21980
rect 58439 21914 58703 21924
rect 58439 20412 58703 20422
rect 58495 20356 58543 20412
rect 58599 20356 58647 20412
rect 58439 20346 58703 20356
rect 58439 18844 58703 18854
rect 58495 18788 58543 18844
rect 58599 18788 58647 18844
rect 58439 18778 58703 18788
rect 58439 17276 58703 17286
rect 58495 17220 58543 17276
rect 58599 17220 58647 17276
rect 58439 17210 58703 17220
rect 58439 15708 58703 15718
rect 58495 15652 58543 15708
rect 58599 15652 58647 15708
rect 58439 15642 58703 15652
rect 58439 14140 58703 14150
rect 58495 14084 58543 14140
rect 58599 14084 58647 14140
rect 58439 14074 58703 14084
rect 57820 13634 58324 13636
rect 57820 13582 57822 13634
rect 57874 13582 58324 13634
rect 57820 13580 58324 13582
rect 57820 13570 57876 13580
rect 58044 13300 58100 13310
rect 57820 13188 57876 13198
rect 57820 11844 57876 13132
rect 57820 11508 57876 11788
rect 58044 13074 58100 13244
rect 58044 13022 58046 13074
rect 58098 13022 58100 13074
rect 57932 11508 57988 11518
rect 57820 11506 57988 11508
rect 57820 11454 57934 11506
rect 57986 11454 57988 11506
rect 57820 11452 57988 11454
rect 57932 11442 57988 11452
rect 57708 10556 57876 10612
rect 57596 10500 57652 10510
rect 57596 10498 57764 10500
rect 57596 10446 57598 10498
rect 57650 10446 57764 10498
rect 57596 10444 57764 10446
rect 57596 10434 57652 10444
rect 57148 10332 57540 10388
rect 56700 10052 56756 10062
rect 56588 9940 56644 9950
rect 56476 9938 56644 9940
rect 56476 9886 56590 9938
rect 56642 9886 56644 9938
rect 56476 9884 56644 9886
rect 56588 9874 56644 9884
rect 56700 9154 56756 9996
rect 56700 9102 56702 9154
rect 56754 9102 56756 9154
rect 56700 9090 56756 9102
rect 57148 9826 57204 10332
rect 57148 9774 57150 9826
rect 57202 9774 57204 9826
rect 56588 9044 56644 9054
rect 56588 8950 56644 8988
rect 57148 8482 57204 9774
rect 57708 9714 57764 10444
rect 57708 9662 57710 9714
rect 57762 9662 57764 9714
rect 57708 9650 57764 9662
rect 57820 9492 57876 10556
rect 57148 8430 57150 8482
rect 57202 8430 57204 8482
rect 57148 8418 57204 8430
rect 57372 9436 57876 9492
rect 56252 8278 56308 8316
rect 56924 8372 56980 8382
rect 55468 8206 55470 8258
rect 55522 8206 55524 8258
rect 55468 8194 55524 8206
rect 55804 8260 55860 8270
rect 55804 6802 55860 8204
rect 56476 8260 56532 8270
rect 56476 8166 56532 8204
rect 56924 7474 56980 8316
rect 57372 8370 57428 9436
rect 57484 9268 57540 9278
rect 58044 9268 58100 13022
rect 58439 12572 58703 12582
rect 58495 12516 58543 12572
rect 58599 12516 58647 12572
rect 58439 12506 58703 12516
rect 58439 11004 58703 11014
rect 58495 10948 58543 11004
rect 58599 10948 58647 11004
rect 58439 10938 58703 10948
rect 58439 9436 58703 9446
rect 58495 9380 58543 9436
rect 58599 9380 58647 9436
rect 58439 9370 58703 9380
rect 57484 9266 58100 9268
rect 57484 9214 57486 9266
rect 57538 9214 58100 9266
rect 57484 9212 58100 9214
rect 57484 9202 57540 9212
rect 57484 9042 57540 9054
rect 57484 8990 57486 9042
rect 57538 8990 57540 9042
rect 57484 8820 57540 8990
rect 57484 8754 57540 8764
rect 57372 8318 57374 8370
rect 57426 8318 57428 8370
rect 56924 7422 56926 7474
rect 56978 7422 56980 7474
rect 56924 7410 56980 7422
rect 57148 8258 57204 8270
rect 57148 8206 57150 8258
rect 57202 8206 57204 8258
rect 57148 7700 57204 8206
rect 56812 7362 56868 7374
rect 56812 7310 56814 7362
rect 56866 7310 56868 7362
rect 56812 6916 56868 7310
rect 56812 6850 56868 6860
rect 57036 7364 57092 7374
rect 55804 6750 55806 6802
rect 55858 6750 55860 6802
rect 55804 6738 55860 6750
rect 55692 6466 55748 6478
rect 55692 6414 55694 6466
rect 55746 6414 55748 6466
rect 55692 5794 55748 6414
rect 55916 6466 55972 6478
rect 55916 6414 55918 6466
rect 55970 6414 55972 6466
rect 55916 6244 55972 6414
rect 56140 6468 56196 6478
rect 56140 6374 56196 6412
rect 57036 6356 57092 7308
rect 57148 6690 57204 7644
rect 57260 8260 57316 8270
rect 57260 7474 57316 8204
rect 57260 7422 57262 7474
rect 57314 7422 57316 7474
rect 57260 7410 57316 7422
rect 57260 6804 57316 6814
rect 57372 6804 57428 8318
rect 58044 8258 58100 8270
rect 58044 8206 58046 8258
rect 58098 8206 58100 8258
rect 58044 6914 58100 8206
rect 58439 7868 58703 7878
rect 58495 7812 58543 7868
rect 58599 7812 58647 7868
rect 58439 7802 58703 7812
rect 58044 6862 58046 6914
rect 58098 6862 58100 6914
rect 58044 6850 58100 6862
rect 57260 6802 57428 6804
rect 57260 6750 57262 6802
rect 57314 6750 57428 6802
rect 57260 6748 57428 6750
rect 57260 6738 57316 6748
rect 58156 6692 58212 6702
rect 57148 6638 57150 6690
rect 57202 6638 57204 6690
rect 57148 6626 57204 6638
rect 57596 6690 58212 6692
rect 57596 6638 58158 6690
rect 58210 6638 58212 6690
rect 57596 6636 58212 6638
rect 55916 6188 56308 6244
rect 55692 5742 55694 5794
rect 55746 5742 55748 5794
rect 55692 5730 55748 5742
rect 55804 6018 55860 6030
rect 55804 5966 55806 6018
rect 55858 5966 55860 6018
rect 55244 5346 55412 5348
rect 55244 5294 55246 5346
rect 55298 5294 55412 5346
rect 55244 5292 55412 5294
rect 55244 5282 55300 5292
rect 54348 5122 54516 5124
rect 54348 5070 54350 5122
rect 54402 5070 54516 5122
rect 54348 5068 54516 5070
rect 55692 5124 55748 5134
rect 55804 5124 55860 5966
rect 56028 5908 56084 5918
rect 55748 5068 55860 5124
rect 55916 5852 56028 5908
rect 55916 5122 55972 5852
rect 56028 5814 56084 5852
rect 56252 5236 56308 6188
rect 56588 5908 56644 5918
rect 56588 5814 56644 5852
rect 57036 5906 57092 6300
rect 57596 6578 57652 6636
rect 58156 6626 58212 6636
rect 57596 6526 57598 6578
rect 57650 6526 57652 6578
rect 57036 5854 57038 5906
rect 57090 5854 57092 5906
rect 57036 5842 57092 5854
rect 57484 5908 57540 5918
rect 57596 5908 57652 6526
rect 57820 6468 57876 6478
rect 57820 6130 57876 6412
rect 58044 6466 58100 6478
rect 58044 6414 58046 6466
rect 58098 6414 58100 6466
rect 58044 6356 58100 6414
rect 58044 6290 58100 6300
rect 58439 6300 58703 6310
rect 58495 6244 58543 6300
rect 58599 6244 58647 6300
rect 58439 6234 58703 6244
rect 57820 6078 57822 6130
rect 57874 6078 57876 6130
rect 57820 6066 57876 6078
rect 57484 5906 57652 5908
rect 57484 5854 57486 5906
rect 57538 5854 57652 5906
rect 57484 5852 57652 5854
rect 58044 6018 58100 6030
rect 58044 5966 58046 6018
rect 58098 5966 58100 6018
rect 57484 5842 57540 5852
rect 56252 5170 56308 5180
rect 56924 5236 56980 5246
rect 55916 5070 55918 5122
rect 55970 5070 55972 5122
rect 54348 5058 54404 5068
rect 55692 5058 55748 5068
rect 55916 5058 55972 5070
rect 56588 5124 56644 5134
rect 56588 5030 56644 5068
rect 56924 5122 56980 5180
rect 56924 5070 56926 5122
rect 56978 5070 56980 5122
rect 56924 5058 56980 5070
rect 58044 5124 58100 5966
rect 58156 5908 58212 5918
rect 58156 5814 58212 5852
rect 58044 5058 58100 5068
rect 54236 4958 54238 5010
rect 54290 4958 54292 5010
rect 54236 4946 54292 4958
rect 58439 4732 58703 4742
rect 58495 4676 58543 4732
rect 58599 4676 58647 4732
rect 58439 4666 58703 4676
rect 52220 4398 52222 4450
rect 52274 4398 52276 4450
rect 52220 4386 52276 4398
rect 56588 4564 56644 4574
rect 51884 4174 51886 4226
rect 51938 4174 51940 4226
rect 51884 4162 51940 4174
rect 51286 3948 51550 3958
rect 51342 3892 51390 3948
rect 51446 3892 51494 3948
rect 51286 3882 51550 3892
rect 56588 3668 56644 4508
rect 56588 3666 56980 3668
rect 56588 3614 56590 3666
rect 56642 3614 56980 3666
rect 56588 3612 56980 3614
rect 56588 3602 56644 3612
rect 52780 3554 52836 3566
rect 52780 3502 52782 3554
rect 52834 3502 52836 3554
rect 50652 3266 50708 3276
rect 51996 3444 52052 3482
rect 52220 3444 52276 3454
rect 51996 3442 52276 3444
rect 51996 3390 51998 3442
rect 52050 3390 52222 3442
rect 52274 3390 52276 3442
rect 51996 3388 52276 3390
rect 51996 800 52052 3388
rect 52220 3378 52276 3388
rect 52780 2660 52836 3502
rect 56924 3554 56980 3612
rect 56924 3502 56926 3554
rect 56978 3502 56980 3554
rect 56924 3490 56980 3502
rect 57372 3666 57428 3678
rect 57372 3614 57374 3666
rect 57426 3614 57428 3666
rect 57372 3388 57428 3614
rect 52780 2594 52836 2604
rect 57036 3332 57428 3388
rect 57036 1652 57092 3332
rect 58439 3164 58703 3174
rect 58495 3108 58543 3164
rect 58599 3108 58647 3164
rect 58439 3098 58703 3108
rect 56924 1596 57092 1652
rect 56924 800 56980 1596
rect 2688 0 2800 800
rect 7616 0 7728 800
rect 12544 0 12656 800
rect 17472 0 17584 800
rect 22400 0 22512 800
rect 27328 0 27440 800
rect 32256 0 32368 800
rect 37184 0 37296 800
rect 42112 0 42224 800
rect 47040 0 47152 800
rect 51968 0 52080 800
rect 56896 0 57008 800
<< via2 >>
rect 1820 36482 1876 36484
rect 1820 36430 1822 36482
rect 1822 36430 1874 36482
rect 1874 36430 1876 36482
rect 1820 36428 1876 36430
rect 1708 35532 1764 35588
rect 1484 35308 1540 35364
rect 1372 34860 1428 34916
rect 1148 33740 1204 33796
rect 1036 29260 1092 29316
rect 1148 14364 1204 14420
rect 1260 28812 1316 28868
rect 2156 35308 2212 35364
rect 1708 34972 1764 35028
rect 2268 34914 2324 34916
rect 2268 34862 2270 34914
rect 2270 34862 2322 34914
rect 2322 34862 2324 34914
rect 2268 34860 2324 34862
rect 1820 34300 1876 34356
rect 2604 36092 2660 36148
rect 3500 37212 3556 37268
rect 2604 34636 2660 34692
rect 3052 34242 3108 34244
rect 3052 34190 3054 34242
rect 3054 34190 3106 34242
rect 3106 34190 3108 34242
rect 3052 34188 3108 34190
rect 2380 34076 2436 34132
rect 1708 33852 1764 33908
rect 1708 33404 1764 33460
rect 1820 33346 1876 33348
rect 1820 33294 1822 33346
rect 1822 33294 1874 33346
rect 1874 33294 1876 33346
rect 1820 33292 1876 33294
rect 1596 32732 1652 32788
rect 1820 32674 1876 32676
rect 1820 32622 1822 32674
rect 1822 32622 1874 32674
rect 1874 32622 1876 32674
rect 1820 32620 1876 32622
rect 1484 26012 1540 26068
rect 1596 32060 1652 32116
rect 1820 31778 1876 31780
rect 1820 31726 1822 31778
rect 1822 31726 1874 31778
rect 1874 31726 1876 31778
rect 1820 31724 1876 31726
rect 1708 30994 1764 30996
rect 1708 30942 1710 30994
rect 1710 30942 1762 30994
rect 1762 30942 1764 30994
rect 1708 30940 1764 30942
rect 1708 30492 1764 30548
rect 1708 30098 1764 30100
rect 1708 30046 1710 30098
rect 1710 30046 1762 30098
rect 1762 30046 1764 30098
rect 1708 30044 1764 30046
rect 1708 28252 1764 28308
rect 2716 33852 2772 33908
rect 3052 33068 3108 33124
rect 2268 32284 2324 32340
rect 2940 31948 2996 32004
rect 2828 31836 2884 31892
rect 2268 31164 2324 31220
rect 2044 30492 2100 30548
rect 1932 29260 1988 29316
rect 2268 30380 2324 30436
rect 2492 30268 2548 30324
rect 2156 29036 2212 29092
rect 2492 30044 2548 30100
rect 2380 29986 2436 29988
rect 2380 29934 2382 29986
rect 2382 29934 2434 29986
rect 2434 29934 2436 29986
rect 2380 29932 2436 29934
rect 2380 29372 2436 29428
rect 2604 29148 2660 29204
rect 1820 28364 1876 28420
rect 1820 27132 1876 27188
rect 1596 21868 1652 21924
rect 1708 24220 1764 24276
rect 1372 16716 1428 16772
rect 1484 21196 1540 21252
rect 4620 36594 4676 36596
rect 4620 36542 4622 36594
rect 4622 36542 4674 36594
rect 4674 36542 4676 36594
rect 4620 36540 4676 36542
rect 5404 36540 5460 36596
rect 4172 36428 4228 36484
rect 4956 35868 5012 35924
rect 4172 35698 4228 35700
rect 4172 35646 4174 35698
rect 4174 35646 4226 35698
rect 4226 35646 4228 35698
rect 4172 35644 4228 35646
rect 5068 35644 5124 35700
rect 3836 35308 3892 35364
rect 3500 34914 3556 34916
rect 3500 34862 3502 34914
rect 3502 34862 3554 34914
rect 3554 34862 3556 34914
rect 3500 34860 3556 34862
rect 4060 34914 4116 34916
rect 4060 34862 4062 34914
rect 4062 34862 4114 34914
rect 4114 34862 4116 34914
rect 4060 34860 4116 34862
rect 5180 34860 5236 34916
rect 3164 32060 3220 32116
rect 3276 33292 3332 33348
rect 3500 33740 3556 33796
rect 4060 33906 4116 33908
rect 4060 33854 4062 33906
rect 4062 33854 4114 33906
rect 4114 33854 4116 33906
rect 4060 33852 4116 33854
rect 3724 32956 3780 33012
rect 4396 34130 4452 34132
rect 4396 34078 4398 34130
rect 4398 34078 4450 34130
rect 4450 34078 4452 34130
rect 4396 34076 4452 34078
rect 4620 33740 4676 33796
rect 4620 33292 4676 33348
rect 4172 32844 4228 32900
rect 3388 32620 3444 32676
rect 3276 31836 3332 31892
rect 3276 31666 3332 31668
rect 3276 31614 3278 31666
rect 3278 31614 3330 31666
rect 3330 31614 3332 31666
rect 3276 31612 3332 31614
rect 3164 30716 3220 30772
rect 3052 29932 3108 29988
rect 2940 29484 2996 29540
rect 3052 29148 3108 29204
rect 3948 32508 4004 32564
rect 3836 31948 3892 32004
rect 4172 32284 4228 32340
rect 4620 31836 4676 31892
rect 3276 28642 3332 28644
rect 3276 28590 3278 28642
rect 3278 28590 3330 28642
rect 3330 28590 3332 28642
rect 3276 28588 3332 28590
rect 3948 29986 4004 29988
rect 3948 29934 3950 29986
rect 3950 29934 4002 29986
rect 4002 29934 4004 29986
rect 3948 29932 4004 29934
rect 4732 31612 4788 31668
rect 4508 30156 4564 30212
rect 5180 31948 5236 32004
rect 4620 30716 4676 30772
rect 5628 35308 5684 35364
rect 6636 36370 6692 36372
rect 6636 36318 6638 36370
rect 6638 36318 6690 36370
rect 6690 36318 6692 36370
rect 6636 36316 6692 36318
rect 7868 36316 7924 36372
rect 5852 35644 5908 35700
rect 6972 35756 7028 35812
rect 6636 34354 6692 34356
rect 6636 34302 6638 34354
rect 6638 34302 6690 34354
rect 6690 34302 6692 34354
rect 6636 34300 6692 34302
rect 6188 33458 6244 33460
rect 6188 33406 6190 33458
rect 6190 33406 6242 33458
rect 6242 33406 6244 33458
rect 6188 33404 6244 33406
rect 6748 32844 6804 32900
rect 5964 32396 6020 32452
rect 5180 31500 5236 31556
rect 4956 31052 5012 31108
rect 3724 29820 3780 29876
rect 3724 28812 3780 28868
rect 3948 28812 4004 28868
rect 3724 28642 3780 28644
rect 3724 28590 3726 28642
rect 3726 28590 3778 28642
rect 3778 28590 3780 28642
rect 3724 28588 3780 28590
rect 3388 28476 3444 28532
rect 2044 25676 2100 25732
rect 2156 24946 2212 24948
rect 2156 24894 2158 24946
rect 2158 24894 2210 24946
rect 2210 24894 2212 24946
rect 2156 24892 2212 24894
rect 2492 26684 2548 26740
rect 2268 24108 2324 24164
rect 1932 23436 1988 23492
rect 1820 21756 1876 21812
rect 2156 23714 2212 23716
rect 2156 23662 2158 23714
rect 2158 23662 2210 23714
rect 2210 23662 2212 23714
rect 2156 23660 2212 23662
rect 4060 28140 4116 28196
rect 4396 28530 4452 28532
rect 4396 28478 4398 28530
rect 4398 28478 4450 28530
rect 4450 28478 4452 28530
rect 4396 28476 4452 28478
rect 4956 30268 5012 30324
rect 5068 30940 5124 30996
rect 4732 30098 4788 30100
rect 4732 30046 4734 30098
rect 4734 30046 4786 30098
rect 4786 30046 4788 30098
rect 4732 30044 4788 30046
rect 4956 29036 5012 29092
rect 4732 28812 4788 28868
rect 5180 30492 5236 30548
rect 4732 28642 4788 28644
rect 4732 28590 4734 28642
rect 4734 28590 4786 28642
rect 4786 28590 4788 28642
rect 4732 28588 4788 28590
rect 3276 26290 3332 26292
rect 3276 26238 3278 26290
rect 3278 26238 3330 26290
rect 3330 26238 3332 26290
rect 3276 26236 3332 26238
rect 2492 24444 2548 24500
rect 3388 25116 3444 25172
rect 2268 23548 2324 23604
rect 3164 24668 3220 24724
rect 3276 24220 3332 24276
rect 3164 24108 3220 24164
rect 2828 23660 2884 23716
rect 2604 23548 2660 23604
rect 2492 23042 2548 23044
rect 2492 22990 2494 23042
rect 2494 22990 2546 23042
rect 2546 22990 2548 23042
rect 2492 22988 2548 22990
rect 2604 22258 2660 22260
rect 2604 22206 2606 22258
rect 2606 22206 2658 22258
rect 2658 22206 2660 22258
rect 2604 22204 2660 22206
rect 1708 20412 1764 20468
rect 2268 21308 2324 21364
rect 2044 20412 2100 20468
rect 1708 19964 1764 20020
rect 1708 19234 1764 19236
rect 1708 19182 1710 19234
rect 1710 19182 1762 19234
rect 1762 19182 1764 19234
rect 1708 19180 1764 19182
rect 2044 19852 2100 19908
rect 1932 19180 1988 19236
rect 1708 18172 1764 18228
rect 1708 17666 1764 17668
rect 1708 17614 1710 17666
rect 1710 17614 1762 17666
rect 1762 17614 1764 17666
rect 1708 17612 1764 17614
rect 1820 16828 1876 16884
rect 1708 15932 1764 15988
rect 2492 21698 2548 21700
rect 2492 21646 2494 21698
rect 2494 21646 2546 21698
rect 2546 21646 2548 21698
rect 2492 21644 2548 21646
rect 3052 22988 3108 23044
rect 2828 21980 2884 22036
rect 4060 25564 4116 25620
rect 4732 28140 4788 28196
rect 5292 28364 5348 28420
rect 5628 31666 5684 31668
rect 5628 31614 5630 31666
rect 5630 31614 5682 31666
rect 5682 31614 5684 31666
rect 5628 31612 5684 31614
rect 6412 32562 6468 32564
rect 6412 32510 6414 32562
rect 6414 32510 6466 32562
rect 6466 32510 6468 32562
rect 6412 32508 6468 32510
rect 8365 36874 8421 36876
rect 8365 36822 8367 36874
rect 8367 36822 8419 36874
rect 8419 36822 8421 36874
rect 8365 36820 8421 36822
rect 8469 36874 8525 36876
rect 8469 36822 8471 36874
rect 8471 36822 8523 36874
rect 8523 36822 8525 36874
rect 8469 36820 8525 36822
rect 8573 36874 8629 36876
rect 8573 36822 8575 36874
rect 8575 36822 8627 36874
rect 8627 36822 8629 36874
rect 9660 36876 9716 36932
rect 10668 36876 10724 36932
rect 8573 36820 8629 36822
rect 8876 35420 8932 35476
rect 8988 35532 9044 35588
rect 8365 35306 8421 35308
rect 8365 35254 8367 35306
rect 8367 35254 8419 35306
rect 8419 35254 8421 35306
rect 8365 35252 8421 35254
rect 8469 35306 8525 35308
rect 8469 35254 8471 35306
rect 8471 35254 8523 35306
rect 8523 35254 8525 35306
rect 8469 35252 8525 35254
rect 8573 35306 8629 35308
rect 8573 35254 8575 35306
rect 8575 35254 8627 35306
rect 8627 35254 8629 35306
rect 8573 35252 8629 35254
rect 9772 35532 9828 35588
rect 11228 36764 11284 36820
rect 11116 35586 11172 35588
rect 11116 35534 11118 35586
rect 11118 35534 11170 35586
rect 11170 35534 11172 35586
rect 11116 35532 11172 35534
rect 10444 35308 10500 35364
rect 9996 34636 10052 34692
rect 7084 33122 7140 33124
rect 7084 33070 7086 33122
rect 7086 33070 7138 33122
rect 7138 33070 7140 33122
rect 7084 33068 7140 33070
rect 8204 34130 8260 34132
rect 8204 34078 8206 34130
rect 8206 34078 8258 34130
rect 8258 34078 8260 34130
rect 8204 34076 8260 34078
rect 8365 33738 8421 33740
rect 8365 33686 8367 33738
rect 8367 33686 8419 33738
rect 8419 33686 8421 33738
rect 8365 33684 8421 33686
rect 8469 33738 8525 33740
rect 8469 33686 8471 33738
rect 8471 33686 8523 33738
rect 8523 33686 8525 33738
rect 8469 33684 8525 33686
rect 8573 33738 8629 33740
rect 8573 33686 8575 33738
rect 8575 33686 8627 33738
rect 8627 33686 8629 33738
rect 8573 33684 8629 33686
rect 8876 33516 8932 33572
rect 8204 33458 8260 33460
rect 8204 33406 8206 33458
rect 8206 33406 8258 33458
rect 8258 33406 8260 33458
rect 8204 33404 8260 33406
rect 8540 33292 8596 33348
rect 7196 32844 7252 32900
rect 6524 31836 6580 31892
rect 6972 32620 7028 32676
rect 6076 31724 6132 31780
rect 6188 30994 6244 30996
rect 6188 30942 6190 30994
rect 6190 30942 6242 30994
rect 6242 30942 6244 30994
rect 6188 30940 6244 30942
rect 5964 30210 6020 30212
rect 5964 30158 5966 30210
rect 5966 30158 6018 30210
rect 6018 30158 6020 30210
rect 5964 30156 6020 30158
rect 6412 30098 6468 30100
rect 6412 30046 6414 30098
rect 6414 30046 6466 30098
rect 6466 30046 6468 30098
rect 6412 30044 6468 30046
rect 7196 32284 7252 32340
rect 7644 31948 7700 32004
rect 7756 32956 7812 33012
rect 7196 31890 7252 31892
rect 7196 31838 7198 31890
rect 7198 31838 7250 31890
rect 7250 31838 7252 31890
rect 7196 31836 7252 31838
rect 7532 31890 7588 31892
rect 7532 31838 7534 31890
rect 7534 31838 7586 31890
rect 7586 31838 7588 31890
rect 7532 31836 7588 31838
rect 6748 30268 6804 30324
rect 5516 29820 5572 29876
rect 5740 29820 5796 29876
rect 5516 29260 5572 29316
rect 6076 29036 6132 29092
rect 5516 28642 5572 28644
rect 5516 28590 5518 28642
rect 5518 28590 5570 28642
rect 5570 28590 5572 28642
rect 5516 28588 5572 28590
rect 5964 28642 6020 28644
rect 5964 28590 5966 28642
rect 5966 28590 6018 28642
rect 6018 28590 6020 28642
rect 5964 28588 6020 28590
rect 4620 26402 4676 26404
rect 4620 26350 4622 26402
rect 4622 26350 4674 26402
rect 4674 26350 4676 26402
rect 4620 26348 4676 26350
rect 3948 25116 4004 25172
rect 4060 24834 4116 24836
rect 4060 24782 4062 24834
rect 4062 24782 4114 24834
rect 4114 24782 4116 24834
rect 4060 24780 4116 24782
rect 3388 23826 3444 23828
rect 3388 23774 3390 23826
rect 3390 23774 3442 23826
rect 3442 23774 3444 23826
rect 3388 23772 3444 23774
rect 3388 22988 3444 23044
rect 3948 24722 4004 24724
rect 3948 24670 3950 24722
rect 3950 24670 4002 24722
rect 4002 24670 4004 24722
rect 3948 24668 4004 24670
rect 4060 24498 4116 24500
rect 4060 24446 4062 24498
rect 4062 24446 4114 24498
rect 4114 24446 4116 24498
rect 4060 24444 4116 24446
rect 4284 26012 4340 26068
rect 3724 22988 3780 23044
rect 3948 22988 4004 23044
rect 3164 21420 3220 21476
rect 3836 21362 3892 21364
rect 3836 21310 3838 21362
rect 3838 21310 3890 21362
rect 3890 21310 3892 21362
rect 3836 21308 3892 21310
rect 2492 20690 2548 20692
rect 2492 20638 2494 20690
rect 2494 20638 2546 20690
rect 2546 20638 2548 20690
rect 2492 20636 2548 20638
rect 2828 21084 2884 21140
rect 3164 21084 3220 21140
rect 3276 20636 3332 20692
rect 3724 20188 3780 20244
rect 3388 20076 3444 20132
rect 2604 19906 2660 19908
rect 2604 19854 2606 19906
rect 2606 19854 2658 19906
rect 2658 19854 2660 19906
rect 2604 19852 2660 19854
rect 2716 19292 2772 19348
rect 2492 18620 2548 18676
rect 3724 19794 3780 19796
rect 3724 19742 3726 19794
rect 3726 19742 3778 19794
rect 3778 19742 3780 19794
rect 3724 19740 3780 19742
rect 4172 20860 4228 20916
rect 4060 19740 4116 19796
rect 3612 19292 3668 19348
rect 3612 19068 3668 19124
rect 3500 18674 3556 18676
rect 3500 18622 3502 18674
rect 3502 18622 3554 18674
rect 3554 18622 3556 18674
rect 3500 18620 3556 18622
rect 4620 26066 4676 26068
rect 4620 26014 4622 26066
rect 4622 26014 4674 26066
rect 4674 26014 4676 26066
rect 4620 26012 4676 26014
rect 4396 24668 4452 24724
rect 4620 23996 4676 24052
rect 5292 27020 5348 27076
rect 4956 26236 5012 26292
rect 4844 25618 4900 25620
rect 4844 25566 4846 25618
rect 4846 25566 4898 25618
rect 4898 25566 4900 25618
rect 4844 25564 4900 25566
rect 4508 23714 4564 23716
rect 4508 23662 4510 23714
rect 4510 23662 4562 23714
rect 4562 23662 4564 23714
rect 4508 23660 4564 23662
rect 4620 23042 4676 23044
rect 4620 22990 4622 23042
rect 4622 22990 4674 23042
rect 4674 22990 4676 23042
rect 4620 22988 4676 22990
rect 4620 22540 4676 22596
rect 4508 22370 4564 22372
rect 4508 22318 4510 22370
rect 4510 22318 4562 22370
rect 4562 22318 4564 22370
rect 4508 22316 4564 22318
rect 4732 22204 4788 22260
rect 4620 21586 4676 21588
rect 4620 21534 4622 21586
rect 4622 21534 4674 21586
rect 4674 21534 4676 21586
rect 4620 21532 4676 21534
rect 4844 21810 4900 21812
rect 4844 21758 4846 21810
rect 4846 21758 4898 21810
rect 4898 21758 4900 21810
rect 4844 21756 4900 21758
rect 4732 21196 4788 21252
rect 4620 20914 4676 20916
rect 4620 20862 4622 20914
rect 4622 20862 4674 20914
rect 4674 20862 4676 20914
rect 4620 20860 4676 20862
rect 5292 20860 5348 20916
rect 4396 20076 4452 20132
rect 4508 20412 4564 20468
rect 4284 18844 4340 18900
rect 2828 17948 2884 18004
rect 3500 17948 3556 18004
rect 3500 17500 3556 17556
rect 2044 17276 2100 17332
rect 3724 17442 3780 17444
rect 3724 17390 3726 17442
rect 3726 17390 3778 17442
rect 3778 17390 3780 17442
rect 3724 17388 3780 17390
rect 4956 20130 5012 20132
rect 4956 20078 4958 20130
rect 4958 20078 5010 20130
rect 5010 20078 5012 20130
rect 4956 20076 5012 20078
rect 5068 19964 5124 20020
rect 5180 20188 5236 20244
rect 3948 17554 4004 17556
rect 3948 17502 3950 17554
rect 3950 17502 4002 17554
rect 4002 17502 4004 17554
rect 3948 17500 4004 17502
rect 4844 18450 4900 18452
rect 4844 18398 4846 18450
rect 4846 18398 4898 18450
rect 4898 18398 4900 18450
rect 4844 18396 4900 18398
rect 5180 18060 5236 18116
rect 4172 17388 4228 17444
rect 2604 17052 2660 17108
rect 1484 14252 1540 14308
rect 2156 16716 2212 16772
rect 1820 15036 1876 15092
rect 2044 14306 2100 14308
rect 2044 14254 2046 14306
rect 2046 14254 2098 14306
rect 2098 14254 2100 14306
rect 2044 14252 2100 14254
rect 2044 13916 2100 13972
rect 2716 16994 2772 16996
rect 2716 16942 2718 16994
rect 2718 16942 2770 16994
rect 2770 16942 2772 16994
rect 2716 16940 2772 16942
rect 3052 16882 3108 16884
rect 3052 16830 3054 16882
rect 3054 16830 3106 16882
rect 3106 16830 3108 16882
rect 3052 16828 3108 16830
rect 2380 14924 2436 14980
rect 3500 14642 3556 14644
rect 3500 14590 3502 14642
rect 3502 14590 3554 14642
rect 3554 14590 3556 14642
rect 3500 14588 3556 14590
rect 3388 14530 3444 14532
rect 3388 14478 3390 14530
rect 3390 14478 3442 14530
rect 3442 14478 3444 14530
rect 3388 14476 3444 14478
rect 4956 16268 5012 16324
rect 4620 16044 4676 16100
rect 5068 15986 5124 15988
rect 5068 15934 5070 15986
rect 5070 15934 5122 15986
rect 5122 15934 5124 15986
rect 5068 15932 5124 15934
rect 4956 15372 5012 15428
rect 3948 14700 4004 14756
rect 4508 14754 4564 14756
rect 4508 14702 4510 14754
rect 4510 14702 4562 14754
rect 4562 14702 4564 14754
rect 4508 14700 4564 14702
rect 4060 14588 4116 14644
rect 2156 13804 2212 13860
rect 2716 14418 2772 14420
rect 2716 14366 2718 14418
rect 2718 14366 2770 14418
rect 2770 14366 2772 14418
rect 2716 14364 2772 14366
rect 2716 13858 2772 13860
rect 2716 13806 2718 13858
rect 2718 13806 2770 13858
rect 2770 13806 2772 13858
rect 2716 13804 2772 13806
rect 2268 13692 2324 13748
rect 1260 12796 1316 12852
rect 1036 10780 1092 10836
rect 1708 12572 1764 12628
rect 1708 10722 1764 10724
rect 1708 10670 1710 10722
rect 1710 10670 1762 10722
rect 1762 10670 1764 10722
rect 1708 10668 1764 10670
rect 1932 11676 1988 11732
rect 3836 14252 3892 14308
rect 3500 13970 3556 13972
rect 3500 13918 3502 13970
rect 3502 13918 3554 13970
rect 3554 13918 3556 13970
rect 3500 13916 3556 13918
rect 2940 13692 2996 13748
rect 2380 12850 2436 12852
rect 2380 12798 2382 12850
rect 2382 12798 2434 12850
rect 2434 12798 2436 12850
rect 2380 12796 2436 12798
rect 1932 11452 1988 11508
rect 2156 11340 2212 11396
rect 2044 10834 2100 10836
rect 2044 10782 2046 10834
rect 2046 10782 2098 10834
rect 2098 10782 2100 10834
rect 2044 10780 2100 10782
rect 2492 11394 2548 11396
rect 2492 11342 2494 11394
rect 2494 11342 2546 11394
rect 2546 11342 2548 11394
rect 2492 11340 2548 11342
rect 2156 10220 2212 10276
rect 1820 9996 1876 10052
rect 2156 9266 2212 9268
rect 2156 9214 2158 9266
rect 2158 9214 2210 9266
rect 2210 9214 2212 9266
rect 2156 9212 2212 9214
rect 1820 9100 1876 9156
rect 2492 10108 2548 10164
rect 2268 7868 2324 7924
rect 2380 9660 2436 9716
rect 2268 7698 2324 7700
rect 2268 7646 2270 7698
rect 2270 7646 2322 7698
rect 2322 7646 2324 7698
rect 2268 7644 2324 7646
rect 1932 6130 1988 6132
rect 1932 6078 1934 6130
rect 1934 6078 1986 6130
rect 1986 6078 1988 6130
rect 1932 6076 1988 6078
rect 2716 9324 2772 9380
rect 2716 9154 2772 9156
rect 2716 9102 2718 9154
rect 2718 9102 2770 9154
rect 2770 9102 2772 9154
rect 2716 9100 2772 9102
rect 3052 12908 3108 12964
rect 3052 12738 3108 12740
rect 3052 12686 3054 12738
rect 3054 12686 3106 12738
rect 3106 12686 3108 12738
rect 3052 12684 3108 12686
rect 3724 13858 3780 13860
rect 3724 13806 3726 13858
rect 3726 13806 3778 13858
rect 3778 13806 3780 13858
rect 3724 13804 3780 13806
rect 3500 12796 3556 12852
rect 3724 12850 3780 12852
rect 3724 12798 3726 12850
rect 3726 12798 3778 12850
rect 3778 12798 3780 12850
rect 3724 12796 3780 12798
rect 3724 12236 3780 12292
rect 4396 14476 4452 14532
rect 3052 11452 3108 11508
rect 3388 11394 3444 11396
rect 3388 11342 3390 11394
rect 3390 11342 3442 11394
rect 3442 11342 3444 11394
rect 3388 11340 3444 11342
rect 3276 11116 3332 11172
rect 3388 10668 3444 10724
rect 2940 9660 2996 9716
rect 3052 9996 3108 10052
rect 3052 9100 3108 9156
rect 2828 7980 2884 8036
rect 3276 7868 3332 7924
rect 2044 5180 2100 5236
rect 4172 12796 4228 12852
rect 3612 11564 3668 11620
rect 3612 11228 3668 11284
rect 4060 11452 4116 11508
rect 3948 11170 4004 11172
rect 3948 11118 3950 11170
rect 3950 11118 4002 11170
rect 4002 11118 4004 11170
rect 3948 11116 4004 11118
rect 5180 15202 5236 15204
rect 5180 15150 5182 15202
rect 5182 15150 5234 15202
rect 5234 15150 5236 15202
rect 5180 15148 5236 15150
rect 4844 14530 4900 14532
rect 4844 14478 4846 14530
rect 4846 14478 4898 14530
rect 4898 14478 4900 14530
rect 4844 14476 4900 14478
rect 4508 14252 4564 14308
rect 4956 14364 5012 14420
rect 4508 14028 4564 14084
rect 4508 11282 4564 11284
rect 4508 11230 4510 11282
rect 4510 11230 4562 11282
rect 4562 11230 4564 11282
rect 4508 11228 4564 11230
rect 4844 13356 4900 13412
rect 5292 13580 5348 13636
rect 4732 12348 4788 12404
rect 4844 12684 4900 12740
rect 5180 12290 5236 12292
rect 5180 12238 5182 12290
rect 5182 12238 5234 12290
rect 5234 12238 5236 12290
rect 5180 12236 5236 12238
rect 5180 12012 5236 12068
rect 4732 11564 4788 11620
rect 5068 11788 5124 11844
rect 4284 9884 4340 9940
rect 3500 7644 3556 7700
rect 3836 7868 3892 7924
rect 4620 9660 4676 9716
rect 4844 9324 4900 9380
rect 4620 8988 4676 9044
rect 5852 28364 5908 28420
rect 6748 28642 6804 28644
rect 6748 28590 6750 28642
rect 6750 28590 6802 28642
rect 6802 28590 6804 28642
rect 6748 28588 6804 28590
rect 5628 27074 5684 27076
rect 5628 27022 5630 27074
rect 5630 27022 5682 27074
rect 5682 27022 5684 27074
rect 5628 27020 5684 27022
rect 5740 24722 5796 24724
rect 5740 24670 5742 24722
rect 5742 24670 5794 24722
rect 5794 24670 5796 24722
rect 5740 24668 5796 24670
rect 5628 21756 5684 21812
rect 5516 20188 5572 20244
rect 8316 32674 8372 32676
rect 8316 32622 8318 32674
rect 8318 32622 8370 32674
rect 8370 32622 8372 32674
rect 8316 32620 8372 32622
rect 9324 33404 9380 33460
rect 9212 32844 9268 32900
rect 9212 32284 9268 32340
rect 8365 32170 8421 32172
rect 8365 32118 8367 32170
rect 8367 32118 8419 32170
rect 8419 32118 8421 32170
rect 8365 32116 8421 32118
rect 8469 32170 8525 32172
rect 8469 32118 8471 32170
rect 8471 32118 8523 32170
rect 8523 32118 8525 32170
rect 8469 32116 8525 32118
rect 8573 32170 8629 32172
rect 8573 32118 8575 32170
rect 8575 32118 8627 32170
rect 8627 32118 8629 32170
rect 8573 32116 8629 32118
rect 8316 31666 8372 31668
rect 8316 31614 8318 31666
rect 8318 31614 8370 31666
rect 8370 31614 8372 31666
rect 8316 31612 8372 31614
rect 8428 31778 8484 31780
rect 8428 31726 8430 31778
rect 8430 31726 8482 31778
rect 8482 31726 8484 31778
rect 8428 31724 8484 31726
rect 7980 31164 8036 31220
rect 7196 29820 7252 29876
rect 7756 29260 7812 29316
rect 8988 31612 9044 31668
rect 8876 31554 8932 31556
rect 8876 31502 8878 31554
rect 8878 31502 8930 31554
rect 8930 31502 8932 31554
rect 8876 31500 8932 31502
rect 8365 30602 8421 30604
rect 8365 30550 8367 30602
rect 8367 30550 8419 30602
rect 8419 30550 8421 30602
rect 8365 30548 8421 30550
rect 8469 30602 8525 30604
rect 8469 30550 8471 30602
rect 8471 30550 8523 30602
rect 8523 30550 8525 30602
rect 8469 30548 8525 30550
rect 8573 30602 8629 30604
rect 8573 30550 8575 30602
rect 8575 30550 8627 30602
rect 8627 30550 8629 30602
rect 8573 30548 8629 30550
rect 8092 30268 8148 30324
rect 8540 29596 8596 29652
rect 8204 29314 8260 29316
rect 8204 29262 8206 29314
rect 8206 29262 8258 29314
rect 8258 29262 8260 29314
rect 8204 29260 8260 29262
rect 8316 29148 8372 29204
rect 8365 29034 8421 29036
rect 8365 28982 8367 29034
rect 8367 28982 8419 29034
rect 8419 28982 8421 29034
rect 8365 28980 8421 28982
rect 8469 29034 8525 29036
rect 8469 28982 8471 29034
rect 8471 28982 8523 29034
rect 8523 28982 8525 29034
rect 8469 28980 8525 28982
rect 8573 29034 8629 29036
rect 8573 28982 8575 29034
rect 8575 28982 8627 29034
rect 8627 28982 8629 29034
rect 8573 28980 8629 28982
rect 8316 28866 8372 28868
rect 8316 28814 8318 28866
rect 8318 28814 8370 28866
rect 8370 28814 8372 28866
rect 8316 28812 8372 28814
rect 8652 28866 8708 28868
rect 8652 28814 8654 28866
rect 8654 28814 8706 28866
rect 8706 28814 8708 28866
rect 8652 28812 8708 28814
rect 7308 27916 7364 27972
rect 6076 26290 6132 26292
rect 6076 26238 6078 26290
rect 6078 26238 6130 26290
rect 6130 26238 6132 26290
rect 6076 26236 6132 26238
rect 6524 26290 6580 26292
rect 6524 26238 6526 26290
rect 6526 26238 6578 26290
rect 6578 26238 6580 26290
rect 6524 26236 6580 26238
rect 6188 25676 6244 25732
rect 5964 22258 6020 22260
rect 5964 22206 5966 22258
rect 5966 22206 6018 22258
rect 6018 22206 6020 22258
rect 5964 22204 6020 22206
rect 6412 24444 6468 24500
rect 6300 24108 6356 24164
rect 7196 26572 7252 26628
rect 6972 23772 7028 23828
rect 6748 22876 6804 22932
rect 8092 27804 8148 27860
rect 7420 26460 7476 26516
rect 7532 26348 7588 26404
rect 7644 24556 7700 24612
rect 8428 27858 8484 27860
rect 8428 27806 8430 27858
rect 8430 27806 8482 27858
rect 8482 27806 8484 27858
rect 8428 27804 8484 27806
rect 8365 27466 8421 27468
rect 8365 27414 8367 27466
rect 8367 27414 8419 27466
rect 8419 27414 8421 27466
rect 8365 27412 8421 27414
rect 8469 27466 8525 27468
rect 8469 27414 8471 27466
rect 8471 27414 8523 27466
rect 8523 27414 8525 27466
rect 8469 27412 8525 27414
rect 8573 27466 8629 27468
rect 8573 27414 8575 27466
rect 8575 27414 8627 27466
rect 8627 27414 8629 27466
rect 8573 27412 8629 27414
rect 10220 34130 10276 34132
rect 10220 34078 10222 34130
rect 10222 34078 10274 34130
rect 10274 34078 10276 34130
rect 10220 34076 10276 34078
rect 9996 33404 10052 33460
rect 9660 32786 9716 32788
rect 9660 32734 9662 32786
rect 9662 32734 9714 32786
rect 9714 32734 9716 32786
rect 9660 32732 9716 32734
rect 11116 34018 11172 34020
rect 11116 33966 11118 34018
rect 11118 33966 11170 34018
rect 11170 33966 11172 34018
rect 11116 33964 11172 33966
rect 10668 32844 10724 32900
rect 10332 32732 10388 32788
rect 9436 32562 9492 32564
rect 9436 32510 9438 32562
rect 9438 32510 9490 32562
rect 9490 32510 9492 32562
rect 9436 32508 9492 32510
rect 9324 32396 9380 32452
rect 10668 32562 10724 32564
rect 10668 32510 10670 32562
rect 10670 32510 10722 32562
rect 10722 32510 10724 32562
rect 10668 32508 10724 32510
rect 10668 31778 10724 31780
rect 10668 31726 10670 31778
rect 10670 31726 10722 31778
rect 10722 31726 10724 31778
rect 10668 31724 10724 31726
rect 10332 31554 10388 31556
rect 10332 31502 10334 31554
rect 10334 31502 10386 31554
rect 10386 31502 10388 31554
rect 10332 31500 10388 31502
rect 10780 31554 10836 31556
rect 10780 31502 10782 31554
rect 10782 31502 10834 31554
rect 10834 31502 10836 31554
rect 10780 31500 10836 31502
rect 10108 30994 10164 30996
rect 10108 30942 10110 30994
rect 10110 30942 10162 30994
rect 10162 30942 10164 30994
rect 10108 30940 10164 30942
rect 10332 30380 10388 30436
rect 9660 29820 9716 29876
rect 9996 30210 10052 30212
rect 9996 30158 9998 30210
rect 9998 30158 10050 30210
rect 10050 30158 10052 30210
rect 9996 30156 10052 30158
rect 9436 29484 9492 29540
rect 9436 28642 9492 28644
rect 9436 28590 9438 28642
rect 9438 28590 9490 28642
rect 9490 28590 9492 28642
rect 9436 28588 9492 28590
rect 9548 29036 9604 29092
rect 9324 28140 9380 28196
rect 8988 26460 9044 26516
rect 8652 26290 8708 26292
rect 8652 26238 8654 26290
rect 8654 26238 8706 26290
rect 8706 26238 8708 26290
rect 8652 26236 8708 26238
rect 8204 26124 8260 26180
rect 8365 25898 8421 25900
rect 8365 25846 8367 25898
rect 8367 25846 8419 25898
rect 8419 25846 8421 25898
rect 8365 25844 8421 25846
rect 8469 25898 8525 25900
rect 8469 25846 8471 25898
rect 8471 25846 8523 25898
rect 8523 25846 8525 25898
rect 8469 25844 8525 25846
rect 8573 25898 8629 25900
rect 8573 25846 8575 25898
rect 8575 25846 8627 25898
rect 8627 25846 8629 25898
rect 8573 25844 8629 25846
rect 8540 25730 8596 25732
rect 8540 25678 8542 25730
rect 8542 25678 8594 25730
rect 8594 25678 8596 25730
rect 8540 25676 8596 25678
rect 8204 25618 8260 25620
rect 8204 25566 8206 25618
rect 8206 25566 8258 25618
rect 8258 25566 8260 25618
rect 8204 25564 8260 25566
rect 7532 24162 7588 24164
rect 7532 24110 7534 24162
rect 7534 24110 7586 24162
rect 7586 24110 7588 24162
rect 7532 24108 7588 24110
rect 7644 23938 7700 23940
rect 7644 23886 7646 23938
rect 7646 23886 7698 23938
rect 7698 23886 7700 23938
rect 7644 23884 7700 23886
rect 7196 22428 7252 22484
rect 7308 22764 7364 22820
rect 7868 23826 7924 23828
rect 7868 23774 7870 23826
rect 7870 23774 7922 23826
rect 7922 23774 7924 23826
rect 7868 23772 7924 23774
rect 7532 22764 7588 22820
rect 7756 22594 7812 22596
rect 7756 22542 7758 22594
rect 7758 22542 7810 22594
rect 7810 22542 7812 22594
rect 7756 22540 7812 22542
rect 5740 19234 5796 19236
rect 5740 19182 5742 19234
rect 5742 19182 5794 19234
rect 5794 19182 5796 19234
rect 5740 19180 5796 19182
rect 5516 18450 5572 18452
rect 5516 18398 5518 18450
rect 5518 18398 5570 18450
rect 5570 18398 5572 18450
rect 5516 18396 5572 18398
rect 5628 17442 5684 17444
rect 5628 17390 5630 17442
rect 5630 17390 5682 17442
rect 5682 17390 5684 17442
rect 5628 17388 5684 17390
rect 6076 18956 6132 19012
rect 6300 19122 6356 19124
rect 6300 19070 6302 19122
rect 6302 19070 6354 19122
rect 6354 19070 6356 19122
rect 6300 19068 6356 19070
rect 7420 20076 7476 20132
rect 6748 19740 6804 19796
rect 6524 19234 6580 19236
rect 6524 19182 6526 19234
rect 6526 19182 6578 19234
rect 6578 19182 6580 19234
rect 6524 19180 6580 19182
rect 7420 19516 7476 19572
rect 5516 15426 5572 15428
rect 5516 15374 5518 15426
rect 5518 15374 5570 15426
rect 5570 15374 5572 15426
rect 5516 15372 5572 15374
rect 5628 15036 5684 15092
rect 6524 18450 6580 18452
rect 6524 18398 6526 18450
rect 6526 18398 6578 18450
rect 6578 18398 6580 18450
rect 6524 18396 6580 18398
rect 6188 18172 6244 18228
rect 6412 18284 6468 18340
rect 6412 17666 6468 17668
rect 6412 17614 6414 17666
rect 6414 17614 6466 17666
rect 6466 17614 6468 17666
rect 6412 17612 6468 17614
rect 6300 16828 6356 16884
rect 6300 16268 6356 16324
rect 6076 15874 6132 15876
rect 6076 15822 6078 15874
rect 6078 15822 6130 15874
rect 6130 15822 6132 15874
rect 6076 15820 6132 15822
rect 5964 15314 6020 15316
rect 5964 15262 5966 15314
rect 5966 15262 6018 15314
rect 6018 15262 6020 15314
rect 5964 15260 6020 15262
rect 5740 14476 5796 14532
rect 6524 15426 6580 15428
rect 6524 15374 6526 15426
rect 6526 15374 6578 15426
rect 6578 15374 6580 15426
rect 6524 15372 6580 15374
rect 6076 14306 6132 14308
rect 6076 14254 6078 14306
rect 6078 14254 6130 14306
rect 6130 14254 6132 14306
rect 6076 14252 6132 14254
rect 5852 13692 5908 13748
rect 5852 13468 5908 13524
rect 5740 12850 5796 12852
rect 5740 12798 5742 12850
rect 5742 12798 5794 12850
rect 5794 12798 5796 12850
rect 5740 12796 5796 12798
rect 5516 12572 5572 12628
rect 5516 11788 5572 11844
rect 5740 12012 5796 12068
rect 5628 11340 5684 11396
rect 5404 11004 5460 11060
rect 5740 11228 5796 11284
rect 5964 11340 6020 11396
rect 5852 11116 5908 11172
rect 5292 9660 5348 9716
rect 5068 9212 5124 9268
rect 5180 9548 5236 9604
rect 4956 8764 5012 8820
rect 3612 6860 3668 6916
rect 3948 6076 4004 6132
rect 4732 7308 4788 7364
rect 5404 9042 5460 9044
rect 5404 8990 5406 9042
rect 5406 8990 5458 9042
rect 5458 8990 5460 9042
rect 5404 8988 5460 8990
rect 5852 10220 5908 10276
rect 7196 19180 7252 19236
rect 8316 24780 8372 24836
rect 8092 24556 8148 24612
rect 8652 24610 8708 24612
rect 8652 24558 8654 24610
rect 8654 24558 8706 24610
rect 8706 24558 8708 24610
rect 8652 24556 8708 24558
rect 8365 24330 8421 24332
rect 8365 24278 8367 24330
rect 8367 24278 8419 24330
rect 8419 24278 8421 24330
rect 8365 24276 8421 24278
rect 8469 24330 8525 24332
rect 8469 24278 8471 24330
rect 8471 24278 8523 24330
rect 8523 24278 8525 24330
rect 8469 24276 8525 24278
rect 8573 24330 8629 24332
rect 8573 24278 8575 24330
rect 8575 24278 8627 24330
rect 8627 24278 8629 24330
rect 8573 24276 8629 24278
rect 8204 23938 8260 23940
rect 8204 23886 8206 23938
rect 8206 23886 8258 23938
rect 8258 23886 8260 23938
rect 8204 23884 8260 23886
rect 8092 22764 8148 22820
rect 8365 22762 8421 22764
rect 8365 22710 8367 22762
rect 8367 22710 8419 22762
rect 8419 22710 8421 22762
rect 8365 22708 8421 22710
rect 8469 22762 8525 22764
rect 8469 22710 8471 22762
rect 8471 22710 8523 22762
rect 8523 22710 8525 22762
rect 8469 22708 8525 22710
rect 8573 22762 8629 22764
rect 8573 22710 8575 22762
rect 8575 22710 8627 22762
rect 8627 22710 8629 22762
rect 8573 22708 8629 22710
rect 8764 22316 8820 22372
rect 8988 21868 9044 21924
rect 9212 26908 9268 26964
rect 10220 29820 10276 29876
rect 10108 29036 10164 29092
rect 9772 28588 9828 28644
rect 10780 30098 10836 30100
rect 10780 30046 10782 30098
rect 10782 30046 10834 30098
rect 10834 30046 10836 30098
rect 10780 30044 10836 30046
rect 11116 29820 11172 29876
rect 10668 28700 10724 28756
rect 10780 28082 10836 28084
rect 10780 28030 10782 28082
rect 10782 28030 10834 28082
rect 10834 28030 10836 28082
rect 10780 28028 10836 28030
rect 13804 37324 13860 37380
rect 12236 36988 12292 37044
rect 12124 35308 12180 35364
rect 11564 34412 11620 34468
rect 11676 34300 11732 34356
rect 11900 34354 11956 34356
rect 11900 34302 11902 34354
rect 11902 34302 11954 34354
rect 11954 34302 11956 34354
rect 11900 34300 11956 34302
rect 11788 33628 11844 33684
rect 12012 33458 12068 33460
rect 12012 33406 12014 33458
rect 12014 33406 12066 33458
rect 12066 33406 12068 33458
rect 12012 33404 12068 33406
rect 11788 32786 11844 32788
rect 11788 32734 11790 32786
rect 11790 32734 11842 32786
rect 11842 32734 11844 32786
rect 11788 32732 11844 32734
rect 11452 32450 11508 32452
rect 11452 32398 11454 32450
rect 11454 32398 11506 32450
rect 11506 32398 11508 32450
rect 11452 32396 11508 32398
rect 11340 30210 11396 30212
rect 11340 30158 11342 30210
rect 11342 30158 11394 30210
rect 11394 30158 11396 30210
rect 11340 30156 11396 30158
rect 12572 36594 12628 36596
rect 12572 36542 12574 36594
rect 12574 36542 12626 36594
rect 12626 36542 12628 36594
rect 12572 36540 12628 36542
rect 13244 36258 13300 36260
rect 13244 36206 13246 36258
rect 13246 36206 13298 36258
rect 13298 36206 13300 36258
rect 13244 36204 13300 36206
rect 13692 36258 13748 36260
rect 13692 36206 13694 36258
rect 13694 36206 13746 36258
rect 13746 36206 13748 36258
rect 13692 36204 13748 36206
rect 14364 36540 14420 36596
rect 16380 36876 16436 36932
rect 17388 36876 17444 36932
rect 18060 36540 18116 36596
rect 14028 36316 14084 36372
rect 12796 35532 12852 35588
rect 13132 35420 13188 35476
rect 13020 34802 13076 34804
rect 13020 34750 13022 34802
rect 13022 34750 13074 34802
rect 13074 34750 13076 34802
rect 13020 34748 13076 34750
rect 12796 34300 12852 34356
rect 12908 33964 12964 34020
rect 12572 33628 12628 33684
rect 13020 33180 13076 33236
rect 12908 31500 12964 31556
rect 13916 33234 13972 33236
rect 13916 33182 13918 33234
rect 13918 33182 13970 33234
rect 13970 33182 13972 33234
rect 13916 33180 13972 33182
rect 15820 36370 15876 36372
rect 15820 36318 15822 36370
rect 15822 36318 15874 36370
rect 15874 36318 15876 36370
rect 15820 36316 15876 36318
rect 16492 36316 16548 36372
rect 15148 36204 15204 36260
rect 16156 36258 16212 36260
rect 16156 36206 16158 36258
rect 16158 36206 16210 36258
rect 16210 36206 16212 36258
rect 16156 36204 16212 36206
rect 15518 36090 15574 36092
rect 15518 36038 15520 36090
rect 15520 36038 15572 36090
rect 15572 36038 15574 36090
rect 15518 36036 15574 36038
rect 15622 36090 15678 36092
rect 15622 36038 15624 36090
rect 15624 36038 15676 36090
rect 15676 36038 15678 36090
rect 15622 36036 15678 36038
rect 15726 36090 15782 36092
rect 15726 36038 15728 36090
rect 15728 36038 15780 36090
rect 15780 36038 15782 36090
rect 15726 36036 15782 36038
rect 15932 35586 15988 35588
rect 15932 35534 15934 35586
rect 15934 35534 15986 35586
rect 15986 35534 15988 35586
rect 15932 35532 15988 35534
rect 14140 34802 14196 34804
rect 14140 34750 14142 34802
rect 14142 34750 14194 34802
rect 14194 34750 14196 34802
rect 14140 34748 14196 34750
rect 15932 35084 15988 35140
rect 15518 34522 15574 34524
rect 15518 34470 15520 34522
rect 15520 34470 15572 34522
rect 15572 34470 15574 34522
rect 15518 34468 15574 34470
rect 15622 34522 15678 34524
rect 15622 34470 15624 34522
rect 15624 34470 15676 34522
rect 15676 34470 15678 34522
rect 15622 34468 15678 34470
rect 15726 34522 15782 34524
rect 15726 34470 15728 34522
rect 15728 34470 15780 34522
rect 15780 34470 15782 34522
rect 15726 34468 15782 34470
rect 16940 35532 16996 35588
rect 17724 34748 17780 34804
rect 14588 32562 14644 32564
rect 14588 32510 14590 32562
rect 14590 32510 14642 32562
rect 14642 32510 14644 32562
rect 14588 32508 14644 32510
rect 14700 32284 14756 32340
rect 13244 31724 13300 31780
rect 12796 29036 12852 29092
rect 12908 29596 12964 29652
rect 11452 28642 11508 28644
rect 11452 28590 11454 28642
rect 11454 28590 11506 28642
rect 11506 28590 11508 28642
rect 11452 28588 11508 28590
rect 11228 28364 11284 28420
rect 11452 28418 11508 28420
rect 11452 28366 11454 28418
rect 11454 28366 11506 28418
rect 11506 28366 11508 28418
rect 11452 28364 11508 28366
rect 11452 27858 11508 27860
rect 11452 27806 11454 27858
rect 11454 27806 11506 27858
rect 11506 27806 11508 27858
rect 11452 27804 11508 27806
rect 9996 26962 10052 26964
rect 9996 26910 9998 26962
rect 9998 26910 10050 26962
rect 10050 26910 10052 26962
rect 9996 26908 10052 26910
rect 9772 26178 9828 26180
rect 9772 26126 9774 26178
rect 9774 26126 9826 26178
rect 9826 26126 9828 26178
rect 9772 26124 9828 26126
rect 10332 26962 10388 26964
rect 10332 26910 10334 26962
rect 10334 26910 10386 26962
rect 10386 26910 10388 26962
rect 10332 26908 10388 26910
rect 11228 27074 11284 27076
rect 11228 27022 11230 27074
rect 11230 27022 11282 27074
rect 11282 27022 11284 27074
rect 11228 27020 11284 27022
rect 11788 27074 11844 27076
rect 11788 27022 11790 27074
rect 11790 27022 11842 27074
rect 11842 27022 11844 27074
rect 11788 27020 11844 27022
rect 10220 26124 10276 26180
rect 9996 25282 10052 25284
rect 9996 25230 9998 25282
rect 9998 25230 10050 25282
rect 10050 25230 10052 25282
rect 9996 25228 10052 25230
rect 10444 25282 10500 25284
rect 10444 25230 10446 25282
rect 10446 25230 10498 25282
rect 10498 25230 10500 25282
rect 10444 25228 10500 25230
rect 9212 23212 9268 23268
rect 9100 21756 9156 21812
rect 9212 22876 9268 22932
rect 8540 21362 8596 21364
rect 8540 21310 8542 21362
rect 8542 21310 8594 21362
rect 8594 21310 8596 21362
rect 8540 21308 8596 21310
rect 8365 21194 8421 21196
rect 8365 21142 8367 21194
rect 8367 21142 8419 21194
rect 8419 21142 8421 21194
rect 8365 21140 8421 21142
rect 8469 21194 8525 21196
rect 8469 21142 8471 21194
rect 8471 21142 8523 21194
rect 8523 21142 8525 21194
rect 8469 21140 8525 21142
rect 8573 21194 8629 21196
rect 8573 21142 8575 21194
rect 8575 21142 8627 21194
rect 8627 21142 8629 21194
rect 8573 21140 8629 21142
rect 7756 19516 7812 19572
rect 8092 19404 8148 19460
rect 7308 18338 7364 18340
rect 7308 18286 7310 18338
rect 7310 18286 7362 18338
rect 7362 18286 7364 18338
rect 7308 18284 7364 18286
rect 7196 17724 7252 17780
rect 6972 16940 7028 16996
rect 7196 16604 7252 16660
rect 6748 16044 6804 16100
rect 6636 14924 6692 14980
rect 6412 14028 6468 14084
rect 6300 13580 6356 13636
rect 7532 18956 7588 19012
rect 7532 18620 7588 18676
rect 7644 18172 7700 18228
rect 6972 14588 7028 14644
rect 7084 13580 7140 13636
rect 6636 12850 6692 12852
rect 6636 12798 6638 12850
rect 6638 12798 6690 12850
rect 6690 12798 6692 12850
rect 6636 12796 6692 12798
rect 6748 12684 6804 12740
rect 7308 15036 7364 15092
rect 7308 14364 7364 14420
rect 7308 13858 7364 13860
rect 7308 13806 7310 13858
rect 7310 13806 7362 13858
rect 7362 13806 7364 13858
rect 7308 13804 7364 13806
rect 6300 11676 6356 11732
rect 6636 11340 6692 11396
rect 6412 11116 6468 11172
rect 6748 11228 6804 11284
rect 6188 9548 6244 9604
rect 6748 9324 6804 9380
rect 6300 9212 6356 9268
rect 5852 8988 5908 9044
rect 7084 11676 7140 11732
rect 7756 17164 7812 17220
rect 7644 16770 7700 16772
rect 7644 16718 7646 16770
rect 7646 16718 7698 16770
rect 7698 16718 7700 16770
rect 7644 16716 7700 16718
rect 7756 15932 7812 15988
rect 8652 19740 8708 19796
rect 8365 19626 8421 19628
rect 8365 19574 8367 19626
rect 8367 19574 8419 19626
rect 8419 19574 8421 19626
rect 8365 19572 8421 19574
rect 8469 19626 8525 19628
rect 8469 19574 8471 19626
rect 8471 19574 8523 19626
rect 8523 19574 8525 19626
rect 8469 19572 8525 19574
rect 8573 19626 8629 19628
rect 8573 19574 8575 19626
rect 8575 19574 8627 19626
rect 8627 19574 8629 19626
rect 8573 19572 8629 19574
rect 9100 19964 9156 20020
rect 9324 22652 9380 22708
rect 9772 23436 9828 23492
rect 9324 21868 9380 21924
rect 10220 24108 10276 24164
rect 10108 22204 10164 22260
rect 9772 21980 9828 22036
rect 9996 21362 10052 21364
rect 9996 21310 9998 21362
rect 9998 21310 10050 21362
rect 10050 21310 10052 21362
rect 9996 21308 10052 21310
rect 9772 20524 9828 20580
rect 8204 19292 8260 19348
rect 8316 19122 8372 19124
rect 8316 19070 8318 19122
rect 8318 19070 8370 19122
rect 8370 19070 8372 19122
rect 8316 19068 8372 19070
rect 8988 19068 9044 19124
rect 8652 18674 8708 18676
rect 8652 18622 8654 18674
rect 8654 18622 8706 18674
rect 8706 18622 8708 18674
rect 8652 18620 8708 18622
rect 8365 18058 8421 18060
rect 8365 18006 8367 18058
rect 8367 18006 8419 18058
rect 8419 18006 8421 18058
rect 8365 18004 8421 18006
rect 8469 18058 8525 18060
rect 8469 18006 8471 18058
rect 8471 18006 8523 18058
rect 8523 18006 8525 18058
rect 8469 18004 8525 18006
rect 8573 18058 8629 18060
rect 8573 18006 8575 18058
rect 8575 18006 8627 18058
rect 8627 18006 8629 18058
rect 8573 18004 8629 18006
rect 7644 14530 7700 14532
rect 7644 14478 7646 14530
rect 7646 14478 7698 14530
rect 7698 14478 7700 14530
rect 7644 14476 7700 14478
rect 7980 17724 8036 17780
rect 8540 17666 8596 17668
rect 8540 17614 8542 17666
rect 8542 17614 8594 17666
rect 8594 17614 8596 17666
rect 8540 17612 8596 17614
rect 9212 18396 9268 18452
rect 9436 18396 9492 18452
rect 12796 28700 12852 28756
rect 12012 28642 12068 28644
rect 12012 28590 12014 28642
rect 12014 28590 12066 28642
rect 12066 28590 12068 28642
rect 12012 28588 12068 28590
rect 12236 28588 12292 28644
rect 12124 28364 12180 28420
rect 12012 26962 12068 26964
rect 12012 26910 12014 26962
rect 12014 26910 12066 26962
rect 12066 26910 12068 26962
rect 12012 26908 12068 26910
rect 13020 29148 13076 29204
rect 13356 29372 13412 29428
rect 13132 27916 13188 27972
rect 13244 29036 13300 29092
rect 12684 26962 12740 26964
rect 12684 26910 12686 26962
rect 12686 26910 12738 26962
rect 12738 26910 12740 26962
rect 12684 26908 12740 26910
rect 12012 26460 12068 26516
rect 11900 25564 11956 25620
rect 11228 25394 11284 25396
rect 11228 25342 11230 25394
rect 11230 25342 11282 25394
rect 11282 25342 11284 25394
rect 11228 25340 11284 25342
rect 11676 25394 11732 25396
rect 11676 25342 11678 25394
rect 11678 25342 11730 25394
rect 11730 25342 11732 25394
rect 11676 25340 11732 25342
rect 12460 25618 12516 25620
rect 12460 25566 12462 25618
rect 12462 25566 12514 25618
rect 12514 25566 12516 25618
rect 12460 25564 12516 25566
rect 12012 25506 12068 25508
rect 12012 25454 12014 25506
rect 12014 25454 12066 25506
rect 12066 25454 12068 25506
rect 12012 25452 12068 25454
rect 12796 25228 12852 25284
rect 11004 24220 11060 24276
rect 11116 24108 11172 24164
rect 10892 22652 10948 22708
rect 10444 21586 10500 21588
rect 10444 21534 10446 21586
rect 10446 21534 10498 21586
rect 10498 21534 10500 21586
rect 10444 21532 10500 21534
rect 10668 21756 10724 21812
rect 12012 23826 12068 23828
rect 12012 23774 12014 23826
rect 12014 23774 12066 23826
rect 12066 23774 12068 23826
rect 12012 23772 12068 23774
rect 12572 23826 12628 23828
rect 12572 23774 12574 23826
rect 12574 23774 12626 23826
rect 12626 23774 12628 23826
rect 12572 23772 12628 23774
rect 12124 23660 12180 23716
rect 11340 22204 11396 22260
rect 10668 20914 10724 20916
rect 10668 20862 10670 20914
rect 10670 20862 10722 20914
rect 10722 20862 10724 20914
rect 10668 20860 10724 20862
rect 10892 21308 10948 21364
rect 10332 20412 10388 20468
rect 10780 20018 10836 20020
rect 10780 19966 10782 20018
rect 10782 19966 10834 20018
rect 10834 19966 10836 20018
rect 10780 19964 10836 19966
rect 10332 19516 10388 19572
rect 9548 17724 9604 17780
rect 8988 17164 9044 17220
rect 9100 17052 9156 17108
rect 9436 17164 9492 17220
rect 8876 16940 8932 16996
rect 8204 16658 8260 16660
rect 8204 16606 8206 16658
rect 8206 16606 8258 16658
rect 8258 16606 8260 16658
rect 8204 16604 8260 16606
rect 8365 16490 8421 16492
rect 8365 16438 8367 16490
rect 8367 16438 8419 16490
rect 8419 16438 8421 16490
rect 8365 16436 8421 16438
rect 8469 16490 8525 16492
rect 8469 16438 8471 16490
rect 8471 16438 8523 16490
rect 8523 16438 8525 16490
rect 8469 16436 8525 16438
rect 8573 16490 8629 16492
rect 8573 16438 8575 16490
rect 8575 16438 8627 16490
rect 8627 16438 8629 16490
rect 8573 16436 8629 16438
rect 7980 15036 8036 15092
rect 8876 16156 8932 16212
rect 8988 16716 9044 16772
rect 8540 16098 8596 16100
rect 8540 16046 8542 16098
rect 8542 16046 8594 16098
rect 8594 16046 8596 16098
rect 8540 16044 8596 16046
rect 9324 16156 9380 16212
rect 9212 16044 9268 16100
rect 8204 15932 8260 15988
rect 8764 15986 8820 15988
rect 8764 15934 8766 15986
rect 8766 15934 8818 15986
rect 8818 15934 8820 15986
rect 8764 15932 8820 15934
rect 8316 15874 8372 15876
rect 8316 15822 8318 15874
rect 8318 15822 8370 15874
rect 8370 15822 8372 15874
rect 8316 15820 8372 15822
rect 8092 14588 8148 14644
rect 8204 15260 8260 15316
rect 7868 14476 7924 14532
rect 7644 14028 7700 14084
rect 7980 14252 8036 14308
rect 8652 15148 8708 15204
rect 8365 14922 8421 14924
rect 8365 14870 8367 14922
rect 8367 14870 8419 14922
rect 8419 14870 8421 14922
rect 8365 14868 8421 14870
rect 8469 14922 8525 14924
rect 8469 14870 8471 14922
rect 8471 14870 8523 14922
rect 8523 14870 8525 14922
rect 8469 14868 8525 14870
rect 8573 14922 8629 14924
rect 8573 14870 8575 14922
rect 8575 14870 8627 14922
rect 8627 14870 8629 14922
rect 8573 14868 8629 14870
rect 7980 13356 8036 13412
rect 8092 13580 8148 13636
rect 7868 12796 7924 12852
rect 8092 12402 8148 12404
rect 8092 12350 8094 12402
rect 8094 12350 8146 12402
rect 8146 12350 8148 12402
rect 8092 12348 8148 12350
rect 8764 14364 8820 14420
rect 8988 14924 9044 14980
rect 8988 14700 9044 14756
rect 8428 13468 8484 13524
rect 8365 13354 8421 13356
rect 8365 13302 8367 13354
rect 8367 13302 8419 13354
rect 8419 13302 8421 13354
rect 8365 13300 8421 13302
rect 8469 13354 8525 13356
rect 8469 13302 8471 13354
rect 8471 13302 8523 13354
rect 8523 13302 8525 13354
rect 8469 13300 8525 13302
rect 8573 13354 8629 13356
rect 8573 13302 8575 13354
rect 8575 13302 8627 13354
rect 8627 13302 8629 13354
rect 8573 13300 8629 13302
rect 8316 13132 8372 13188
rect 9324 15260 9380 15316
rect 9100 13468 9156 13524
rect 8988 12684 9044 12740
rect 7644 11676 7700 11732
rect 7868 11282 7924 11284
rect 7868 11230 7870 11282
rect 7870 11230 7922 11282
rect 7922 11230 7924 11282
rect 7868 11228 7924 11230
rect 7756 11004 7812 11060
rect 7644 10668 7700 10724
rect 6972 9212 7028 9268
rect 7644 9042 7700 9044
rect 7644 8990 7646 9042
rect 7646 8990 7698 9042
rect 7698 8990 7700 9042
rect 7644 8988 7700 8990
rect 7868 10780 7924 10836
rect 8365 11786 8421 11788
rect 8365 11734 8367 11786
rect 8367 11734 8419 11786
rect 8419 11734 8421 11786
rect 8365 11732 8421 11734
rect 8469 11786 8525 11788
rect 8469 11734 8471 11786
rect 8471 11734 8523 11786
rect 8523 11734 8525 11786
rect 8469 11732 8525 11734
rect 8573 11786 8629 11788
rect 8573 11734 8575 11786
rect 8575 11734 8627 11786
rect 8627 11734 8629 11786
rect 8573 11732 8629 11734
rect 9212 12850 9268 12852
rect 9212 12798 9214 12850
rect 9214 12798 9266 12850
rect 9266 12798 9268 12850
rect 9212 12796 9268 12798
rect 9100 11900 9156 11956
rect 8316 11004 8372 11060
rect 8204 10780 8260 10836
rect 8316 10668 8372 10724
rect 8652 10556 8708 10612
rect 8365 10218 8421 10220
rect 8365 10166 8367 10218
rect 8367 10166 8419 10218
rect 8419 10166 8421 10218
rect 8365 10164 8421 10166
rect 8469 10218 8525 10220
rect 8469 10166 8471 10218
rect 8471 10166 8523 10218
rect 8523 10166 8525 10218
rect 8469 10164 8525 10166
rect 8573 10218 8629 10220
rect 8573 10166 8575 10218
rect 8575 10166 8627 10218
rect 8627 10166 8629 10218
rect 8573 10164 8629 10166
rect 8764 9996 8820 10052
rect 5740 8034 5796 8036
rect 5740 7982 5742 8034
rect 5742 7982 5794 8034
rect 5794 7982 5796 8034
rect 5740 7980 5796 7982
rect 5628 7644 5684 7700
rect 5964 7474 6020 7476
rect 5964 7422 5966 7474
rect 5966 7422 6018 7474
rect 6018 7422 6020 7474
rect 5964 7420 6020 7422
rect 6636 7698 6692 7700
rect 6636 7646 6638 7698
rect 6638 7646 6690 7698
rect 6690 7646 6692 7698
rect 6636 7644 6692 7646
rect 7196 7644 7252 7700
rect 5516 7362 5572 7364
rect 5516 7310 5518 7362
rect 5518 7310 5570 7362
rect 5570 7310 5572 7362
rect 5516 7308 5572 7310
rect 6748 7362 6804 7364
rect 6748 7310 6750 7362
rect 6750 7310 6802 7362
rect 6802 7310 6804 7362
rect 6748 7308 6804 7310
rect 5404 7196 5460 7252
rect 7196 7474 7252 7476
rect 7196 7422 7198 7474
rect 7198 7422 7250 7474
rect 7250 7422 7252 7474
rect 7196 7420 7252 7422
rect 7308 7362 7364 7364
rect 7308 7310 7310 7362
rect 7310 7310 7362 7362
rect 7362 7310 7364 7362
rect 7308 7308 7364 7310
rect 6860 7196 6916 7252
rect 4956 6636 5012 6692
rect 3612 5906 3668 5908
rect 3612 5854 3614 5906
rect 3614 5854 3666 5906
rect 3666 5854 3668 5906
rect 3612 5852 3668 5854
rect 3948 5180 4004 5236
rect 4396 3612 4452 3668
rect 5292 6130 5348 6132
rect 5292 6078 5294 6130
rect 5294 6078 5346 6130
rect 5346 6078 5348 6130
rect 5292 6076 5348 6078
rect 5740 6690 5796 6692
rect 5740 6638 5742 6690
rect 5742 6638 5794 6690
rect 5794 6638 5796 6690
rect 5740 6636 5796 6638
rect 6188 6524 6244 6580
rect 5964 6076 6020 6132
rect 6300 5906 6356 5908
rect 6300 5854 6302 5906
rect 6302 5854 6354 5906
rect 6354 5854 6356 5906
rect 6300 5852 6356 5854
rect 7756 7196 7812 7252
rect 6524 6076 6580 6132
rect 6748 5964 6804 6020
rect 6636 5292 6692 5348
rect 6412 4898 6468 4900
rect 6412 4846 6414 4898
rect 6414 4846 6466 4898
rect 6466 4846 6468 4898
rect 6412 4844 6468 4846
rect 6300 3666 6356 3668
rect 6300 3614 6302 3666
rect 6302 3614 6354 3666
rect 6354 3614 6356 3666
rect 6300 3612 6356 3614
rect 7868 6076 7924 6132
rect 7868 5180 7924 5236
rect 7644 3724 7700 3780
rect 7196 3666 7252 3668
rect 7196 3614 7198 3666
rect 7198 3614 7250 3666
rect 7250 3614 7252 3666
rect 7196 3612 7252 3614
rect 5852 3442 5908 3444
rect 5852 3390 5854 3442
rect 5854 3390 5906 3442
rect 5906 3390 5908 3442
rect 5852 3388 5908 3390
rect 8204 9324 8260 9380
rect 8204 8818 8260 8820
rect 8204 8766 8206 8818
rect 8206 8766 8258 8818
rect 8258 8766 8260 8818
rect 8204 8764 8260 8766
rect 8540 8818 8596 8820
rect 8540 8766 8542 8818
rect 8542 8766 8594 8818
rect 8594 8766 8596 8818
rect 8540 8764 8596 8766
rect 8365 8650 8421 8652
rect 8365 8598 8367 8650
rect 8367 8598 8419 8650
rect 8419 8598 8421 8650
rect 8365 8596 8421 8598
rect 8469 8650 8525 8652
rect 8469 8598 8471 8650
rect 8471 8598 8523 8650
rect 8523 8598 8525 8650
rect 8469 8596 8525 8598
rect 8573 8650 8629 8652
rect 8573 8598 8575 8650
rect 8575 8598 8627 8650
rect 8627 8598 8629 8650
rect 8573 8596 8629 8598
rect 8764 8034 8820 8036
rect 8764 7982 8766 8034
rect 8766 7982 8818 8034
rect 8818 7982 8820 8034
rect 8764 7980 8820 7982
rect 8652 7308 8708 7364
rect 8316 7196 8372 7252
rect 8365 7082 8421 7084
rect 8365 7030 8367 7082
rect 8367 7030 8419 7082
rect 8419 7030 8421 7082
rect 8365 7028 8421 7030
rect 8469 7082 8525 7084
rect 8469 7030 8471 7082
rect 8471 7030 8523 7082
rect 8523 7030 8525 7082
rect 8469 7028 8525 7030
rect 8573 7082 8629 7084
rect 8573 7030 8575 7082
rect 8575 7030 8627 7082
rect 8627 7030 8629 7082
rect 8573 7028 8629 7030
rect 9548 16994 9604 16996
rect 9548 16942 9550 16994
rect 9550 16942 9602 16994
rect 9602 16942 9604 16994
rect 9548 16940 9604 16942
rect 9548 16604 9604 16660
rect 9772 17500 9828 17556
rect 9772 16770 9828 16772
rect 9772 16718 9774 16770
rect 9774 16718 9826 16770
rect 9826 16718 9828 16770
rect 9772 16716 9828 16718
rect 10444 19122 10500 19124
rect 10444 19070 10446 19122
rect 10446 19070 10498 19122
rect 10498 19070 10500 19122
rect 10444 19068 10500 19070
rect 10332 18450 10388 18452
rect 10332 18398 10334 18450
rect 10334 18398 10386 18450
rect 10386 18398 10388 18450
rect 10332 18396 10388 18398
rect 10780 19516 10836 19572
rect 10556 18396 10612 18452
rect 10444 18060 10500 18116
rect 10220 17724 10276 17780
rect 10108 17052 10164 17108
rect 9884 16604 9940 16660
rect 9548 15148 9604 15204
rect 9772 15260 9828 15316
rect 9772 15036 9828 15092
rect 10220 15596 10276 15652
rect 10108 15372 10164 15428
rect 9884 14700 9940 14756
rect 9884 14530 9940 14532
rect 9884 14478 9886 14530
rect 9886 14478 9938 14530
rect 9938 14478 9940 14530
rect 9884 14476 9940 14478
rect 10108 14252 10164 14308
rect 10220 14476 10276 14532
rect 9548 13746 9604 13748
rect 9548 13694 9550 13746
rect 9550 13694 9602 13746
rect 9602 13694 9604 13746
rect 9548 13692 9604 13694
rect 10108 13634 10164 13636
rect 10108 13582 10110 13634
rect 10110 13582 10162 13634
rect 10162 13582 10164 13634
rect 10108 13580 10164 13582
rect 9772 13522 9828 13524
rect 9772 13470 9774 13522
rect 9774 13470 9826 13522
rect 9826 13470 9828 13522
rect 9772 13468 9828 13470
rect 9548 12460 9604 12516
rect 9212 11394 9268 11396
rect 9212 11342 9214 11394
rect 9214 11342 9266 11394
rect 9266 11342 9268 11394
rect 9212 11340 9268 11342
rect 8988 10610 9044 10612
rect 8988 10558 8990 10610
rect 8990 10558 9042 10610
rect 9042 10558 9044 10610
rect 8988 10556 9044 10558
rect 8988 9100 9044 9156
rect 10556 16716 10612 16772
rect 11452 20860 11508 20916
rect 11340 20802 11396 20804
rect 11340 20750 11342 20802
rect 11342 20750 11394 20802
rect 11394 20750 11396 20802
rect 11340 20748 11396 20750
rect 12236 23212 12292 23268
rect 12796 23100 12852 23156
rect 12684 23042 12740 23044
rect 12684 22990 12686 23042
rect 12686 22990 12738 23042
rect 12738 22990 12740 23042
rect 12684 22988 12740 22990
rect 13020 22370 13076 22372
rect 13020 22318 13022 22370
rect 13022 22318 13074 22370
rect 13074 22318 13076 22370
rect 13020 22316 13076 22318
rect 12684 22258 12740 22260
rect 12684 22206 12686 22258
rect 12686 22206 12738 22258
rect 12738 22206 12740 22258
rect 12684 22204 12740 22206
rect 11116 20076 11172 20132
rect 11452 20018 11508 20020
rect 11452 19966 11454 20018
rect 11454 19966 11506 20018
rect 11506 19966 11508 20018
rect 11452 19964 11508 19966
rect 11116 19906 11172 19908
rect 11116 19854 11118 19906
rect 11118 19854 11170 19906
rect 11170 19854 11172 19906
rect 11116 19852 11172 19854
rect 11788 20076 11844 20132
rect 11900 19852 11956 19908
rect 12124 20300 12180 20356
rect 11452 19068 11508 19124
rect 11452 18396 11508 18452
rect 10892 18060 10948 18116
rect 10668 17612 10724 17668
rect 11452 17612 11508 17668
rect 12572 20076 12628 20132
rect 12460 19852 12516 19908
rect 12796 19292 12852 19348
rect 12684 19180 12740 19236
rect 12796 19122 12852 19124
rect 12796 19070 12798 19122
rect 12798 19070 12850 19122
rect 12850 19070 12852 19122
rect 12796 19068 12852 19070
rect 12908 18508 12964 18564
rect 12684 18172 12740 18228
rect 12908 18060 12964 18116
rect 11004 17442 11060 17444
rect 11004 17390 11006 17442
rect 11006 17390 11058 17442
rect 11058 17390 11060 17442
rect 11004 17388 11060 17390
rect 10668 16268 10724 16324
rect 10892 16994 10948 16996
rect 10892 16942 10894 16994
rect 10894 16942 10946 16994
rect 10946 16942 10948 16994
rect 10892 16940 10948 16942
rect 11788 17724 11844 17780
rect 10668 15932 10724 15988
rect 10780 15372 10836 15428
rect 10668 15148 10724 15204
rect 10556 14812 10612 14868
rect 10668 14530 10724 14532
rect 10668 14478 10670 14530
rect 10670 14478 10722 14530
rect 10722 14478 10724 14530
rect 10668 14476 10724 14478
rect 10556 13804 10612 13860
rect 11340 16098 11396 16100
rect 11340 16046 11342 16098
rect 11342 16046 11394 16098
rect 11394 16046 11396 16098
rect 11340 16044 11396 16046
rect 11452 15874 11508 15876
rect 11452 15822 11454 15874
rect 11454 15822 11506 15874
rect 11506 15822 11508 15874
rect 11452 15820 11508 15822
rect 11228 14700 11284 14756
rect 11452 15538 11508 15540
rect 11452 15486 11454 15538
rect 11454 15486 11506 15538
rect 11506 15486 11508 15538
rect 11452 15484 11508 15486
rect 11564 15148 11620 15204
rect 11004 14418 11060 14420
rect 11004 14366 11006 14418
rect 11006 14366 11058 14418
rect 11058 14366 11060 14418
rect 11004 14364 11060 14366
rect 10444 11564 10500 11620
rect 10892 13522 10948 13524
rect 10892 13470 10894 13522
rect 10894 13470 10946 13522
rect 10946 13470 10948 13522
rect 10892 13468 10948 13470
rect 10892 12684 10948 12740
rect 9884 11340 9940 11396
rect 9996 10444 10052 10500
rect 9772 9884 9828 9940
rect 9436 9714 9492 9716
rect 9436 9662 9438 9714
rect 9438 9662 9490 9714
rect 9490 9662 9492 9714
rect 9436 9660 9492 9662
rect 9548 9548 9604 9604
rect 9660 9324 9716 9380
rect 9772 9548 9828 9604
rect 9660 8930 9716 8932
rect 9660 8878 9662 8930
rect 9662 8878 9714 8930
rect 9714 8878 9716 8930
rect 9660 8876 9716 8878
rect 10220 9772 10276 9828
rect 10220 9212 10276 9268
rect 9996 8876 10052 8932
rect 10220 8764 10276 8820
rect 8988 6524 9044 6580
rect 8988 6130 9044 6132
rect 8988 6078 8990 6130
rect 8990 6078 9042 6130
rect 9042 6078 9044 6130
rect 8988 6076 9044 6078
rect 8652 6018 8708 6020
rect 8652 5966 8654 6018
rect 8654 5966 8706 6018
rect 8706 5966 8708 6018
rect 8652 5964 8708 5966
rect 8365 5514 8421 5516
rect 8365 5462 8367 5514
rect 8367 5462 8419 5514
rect 8419 5462 8421 5514
rect 8365 5460 8421 5462
rect 8469 5514 8525 5516
rect 8469 5462 8471 5514
rect 8471 5462 8523 5514
rect 8523 5462 8525 5514
rect 8469 5460 8525 5462
rect 8573 5514 8629 5516
rect 8573 5462 8575 5514
rect 8575 5462 8627 5514
rect 8627 5462 8629 5514
rect 8573 5460 8629 5462
rect 8876 5516 8932 5572
rect 9660 6076 9716 6132
rect 10444 9884 10500 9940
rect 10668 10444 10724 10500
rect 10668 9826 10724 9828
rect 10668 9774 10670 9826
rect 10670 9774 10722 9826
rect 10722 9774 10724 9826
rect 10668 9772 10724 9774
rect 10556 9660 10612 9716
rect 10668 9602 10724 9604
rect 10668 9550 10670 9602
rect 10670 9550 10722 9602
rect 10722 9550 10724 9602
rect 10668 9548 10724 9550
rect 11228 13468 11284 13524
rect 11340 14252 11396 14308
rect 11228 13132 11284 13188
rect 11228 12684 11284 12740
rect 11564 14476 11620 14532
rect 11788 14476 11844 14532
rect 11564 13804 11620 13860
rect 11564 13634 11620 13636
rect 11564 13582 11566 13634
rect 11566 13582 11618 13634
rect 11618 13582 11620 13634
rect 11564 13580 11620 13582
rect 11676 12850 11732 12852
rect 11676 12798 11678 12850
rect 11678 12798 11730 12850
rect 11730 12798 11732 12850
rect 11676 12796 11732 12798
rect 12572 17724 12628 17780
rect 12124 17666 12180 17668
rect 12124 17614 12126 17666
rect 12126 17614 12178 17666
rect 12178 17614 12180 17666
rect 12124 17612 12180 17614
rect 13804 29650 13860 29652
rect 13804 29598 13806 29650
rect 13806 29598 13858 29650
rect 13858 29598 13860 29650
rect 13804 29596 13860 29598
rect 13580 29148 13636 29204
rect 14252 31778 14308 31780
rect 14252 31726 14254 31778
rect 14254 31726 14306 31778
rect 14306 31726 14308 31778
rect 14252 31724 14308 31726
rect 14812 31164 14868 31220
rect 15518 32954 15574 32956
rect 15518 32902 15520 32954
rect 15520 32902 15572 32954
rect 15572 32902 15574 32954
rect 15518 32900 15574 32902
rect 15622 32954 15678 32956
rect 15622 32902 15624 32954
rect 15624 32902 15676 32954
rect 15676 32902 15678 32954
rect 15622 32900 15678 32902
rect 15726 32954 15782 32956
rect 15726 32902 15728 32954
rect 15728 32902 15780 32954
rect 15780 32902 15782 32954
rect 15726 32900 15782 32902
rect 16156 32844 16212 32900
rect 16828 32844 16884 32900
rect 16156 32674 16212 32676
rect 16156 32622 16158 32674
rect 16158 32622 16210 32674
rect 16210 32622 16212 32674
rect 16156 32620 16212 32622
rect 15148 32396 15204 32452
rect 15372 32562 15428 32564
rect 15372 32510 15374 32562
rect 15374 32510 15426 32562
rect 15426 32510 15428 32562
rect 15372 32508 15428 32510
rect 15372 32284 15428 32340
rect 15820 32284 15876 32340
rect 15596 32060 15652 32116
rect 14924 31052 14980 31108
rect 16044 32450 16100 32452
rect 16044 32398 16046 32450
rect 16046 32398 16098 32450
rect 16098 32398 16100 32450
rect 16044 32396 16100 32398
rect 17836 34636 17892 34692
rect 22672 36874 22728 36876
rect 22672 36822 22674 36874
rect 22674 36822 22726 36874
rect 22726 36822 22728 36874
rect 22672 36820 22728 36822
rect 22776 36874 22832 36876
rect 22776 36822 22778 36874
rect 22778 36822 22830 36874
rect 22830 36822 22832 36874
rect 22776 36820 22832 36822
rect 22880 36874 22936 36876
rect 22880 36822 22882 36874
rect 22882 36822 22934 36874
rect 22934 36822 22936 36874
rect 22880 36820 22936 36822
rect 27692 37212 27748 37268
rect 21196 36428 21252 36484
rect 18508 36258 18564 36260
rect 18508 36206 18510 36258
rect 18510 36206 18562 36258
rect 18562 36206 18564 36258
rect 18508 36204 18564 36206
rect 18172 35532 18228 35588
rect 20300 35980 20356 36036
rect 18844 35532 18900 35588
rect 18732 34802 18788 34804
rect 18732 34750 18734 34802
rect 18734 34750 18786 34802
rect 18786 34750 18788 34802
rect 18732 34748 18788 34750
rect 18060 32732 18116 32788
rect 18172 34524 18228 34580
rect 16268 32060 16324 32116
rect 15518 31386 15574 31388
rect 15518 31334 15520 31386
rect 15520 31334 15572 31386
rect 15572 31334 15574 31386
rect 15518 31332 15574 31334
rect 15622 31386 15678 31388
rect 15622 31334 15624 31386
rect 15624 31334 15676 31386
rect 15676 31334 15678 31386
rect 15622 31332 15678 31334
rect 15726 31386 15782 31388
rect 15726 31334 15728 31386
rect 15728 31334 15780 31386
rect 15780 31334 15782 31386
rect 15726 31332 15782 31334
rect 16492 31778 16548 31780
rect 16492 31726 16494 31778
rect 16494 31726 16546 31778
rect 16546 31726 16548 31778
rect 16492 31724 16548 31726
rect 16716 32060 16772 32116
rect 14700 29820 14756 29876
rect 14924 30156 14980 30212
rect 15036 29932 15092 29988
rect 15820 31218 15876 31220
rect 15820 31166 15822 31218
rect 15822 31166 15874 31218
rect 15874 31166 15876 31218
rect 15820 31164 15876 31166
rect 16604 31052 16660 31108
rect 15518 29818 15574 29820
rect 15518 29766 15520 29818
rect 15520 29766 15572 29818
rect 15572 29766 15574 29818
rect 15518 29764 15574 29766
rect 15622 29818 15678 29820
rect 15622 29766 15624 29818
rect 15624 29766 15676 29818
rect 15676 29766 15678 29818
rect 15622 29764 15678 29766
rect 15726 29818 15782 29820
rect 15726 29766 15728 29818
rect 15728 29766 15780 29818
rect 15780 29766 15782 29818
rect 15726 29764 15782 29766
rect 14476 28700 14532 28756
rect 13468 26572 13524 26628
rect 13356 25676 13412 25732
rect 13692 25676 13748 25732
rect 13356 24108 13412 24164
rect 13468 24220 13524 24276
rect 13356 23100 13412 23156
rect 13356 22092 13412 22148
rect 13692 23212 13748 23268
rect 13916 27804 13972 27860
rect 14812 27746 14868 27748
rect 14812 27694 14814 27746
rect 14814 27694 14866 27746
rect 14866 27694 14868 27746
rect 14812 27692 14868 27694
rect 14252 27580 14308 27636
rect 15518 28250 15574 28252
rect 15518 28198 15520 28250
rect 15520 28198 15572 28250
rect 15572 28198 15574 28250
rect 15518 28196 15574 28198
rect 15622 28250 15678 28252
rect 15622 28198 15624 28250
rect 15624 28198 15676 28250
rect 15676 28198 15678 28250
rect 15622 28196 15678 28198
rect 15726 28250 15782 28252
rect 15726 28198 15728 28250
rect 15728 28198 15780 28250
rect 15780 28198 15782 28250
rect 15726 28196 15782 28198
rect 14028 26908 14084 26964
rect 15708 27244 15764 27300
rect 15932 27132 15988 27188
rect 15518 26682 15574 26684
rect 15518 26630 15520 26682
rect 15520 26630 15572 26682
rect 15572 26630 15574 26682
rect 15518 26628 15574 26630
rect 15622 26682 15678 26684
rect 15622 26630 15624 26682
rect 15624 26630 15676 26682
rect 15676 26630 15678 26682
rect 15622 26628 15678 26630
rect 15726 26682 15782 26684
rect 15726 26630 15728 26682
rect 15728 26630 15780 26682
rect 15780 26630 15782 26682
rect 15726 26628 15782 26630
rect 14364 25676 14420 25732
rect 15036 25452 15092 25508
rect 15596 26124 15652 26180
rect 15820 25506 15876 25508
rect 15820 25454 15822 25506
rect 15822 25454 15874 25506
rect 15874 25454 15876 25506
rect 15820 25452 15876 25454
rect 14028 25282 14084 25284
rect 14028 25230 14030 25282
rect 14030 25230 14082 25282
rect 14082 25230 14084 25282
rect 14028 25228 14084 25230
rect 15518 25114 15574 25116
rect 15518 25062 15520 25114
rect 15520 25062 15572 25114
rect 15572 25062 15574 25114
rect 15518 25060 15574 25062
rect 15622 25114 15678 25116
rect 15622 25062 15624 25114
rect 15624 25062 15676 25114
rect 15676 25062 15678 25114
rect 15622 25060 15678 25062
rect 15726 25114 15782 25116
rect 15726 25062 15728 25114
rect 15728 25062 15780 25114
rect 15780 25062 15782 25114
rect 15726 25060 15782 25062
rect 15484 24892 15540 24948
rect 15484 24722 15540 24724
rect 15484 24670 15486 24722
rect 15486 24670 15538 24722
rect 15538 24670 15540 24722
rect 15484 24668 15540 24670
rect 16380 26460 16436 26516
rect 16492 26178 16548 26180
rect 16492 26126 16494 26178
rect 16494 26126 16546 26178
rect 16546 26126 16548 26178
rect 16492 26124 16548 26126
rect 16268 25116 16324 25172
rect 16380 25564 16436 25620
rect 15036 24610 15092 24612
rect 15036 24558 15038 24610
rect 15038 24558 15090 24610
rect 15090 24558 15092 24610
rect 15036 24556 15092 24558
rect 13916 23212 13972 23268
rect 14140 23154 14196 23156
rect 14140 23102 14142 23154
rect 14142 23102 14194 23154
rect 14194 23102 14196 23154
rect 14140 23100 14196 23102
rect 13804 22876 13860 22932
rect 14252 22764 14308 22820
rect 14700 22764 14756 22820
rect 13916 22540 13972 22596
rect 13692 22258 13748 22260
rect 13692 22206 13694 22258
rect 13694 22206 13746 22258
rect 13746 22206 13748 22258
rect 14588 22258 14644 22260
rect 13692 22204 13748 22206
rect 13804 22146 13860 22148
rect 13804 22094 13806 22146
rect 13806 22094 13858 22146
rect 13858 22094 13860 22146
rect 13804 22092 13860 22094
rect 14588 22206 14590 22258
rect 14590 22206 14642 22258
rect 14642 22206 14644 22258
rect 14588 22204 14644 22206
rect 14028 21980 14084 22036
rect 13468 21756 13524 21812
rect 13916 21756 13972 21812
rect 13356 21474 13412 21476
rect 13356 21422 13358 21474
rect 13358 21422 13410 21474
rect 13410 21422 13412 21474
rect 13356 21420 13412 21422
rect 13692 20578 13748 20580
rect 13692 20526 13694 20578
rect 13694 20526 13746 20578
rect 13746 20526 13748 20578
rect 13692 20524 13748 20526
rect 13916 20524 13972 20580
rect 14364 22146 14420 22148
rect 14364 22094 14366 22146
rect 14366 22094 14418 22146
rect 14418 22094 14420 22146
rect 14364 22092 14420 22094
rect 14700 21810 14756 21812
rect 14700 21758 14702 21810
rect 14702 21758 14754 21810
rect 14754 21758 14756 21810
rect 14700 21756 14756 21758
rect 14140 21644 14196 21700
rect 14364 21698 14420 21700
rect 14364 21646 14366 21698
rect 14366 21646 14418 21698
rect 14418 21646 14420 21698
rect 14364 21644 14420 21646
rect 15518 23546 15574 23548
rect 15518 23494 15520 23546
rect 15520 23494 15572 23546
rect 15572 23494 15574 23546
rect 15518 23492 15574 23494
rect 15622 23546 15678 23548
rect 15622 23494 15624 23546
rect 15624 23494 15676 23546
rect 15676 23494 15678 23546
rect 15622 23492 15678 23494
rect 15726 23546 15782 23548
rect 15726 23494 15728 23546
rect 15728 23494 15780 23546
rect 15780 23494 15782 23546
rect 15726 23492 15782 23494
rect 15708 23378 15764 23380
rect 15708 23326 15710 23378
rect 15710 23326 15762 23378
rect 15762 23326 15764 23378
rect 15708 23324 15764 23326
rect 15036 22988 15092 23044
rect 15932 23154 15988 23156
rect 15932 23102 15934 23154
rect 15934 23102 15986 23154
rect 15986 23102 15988 23154
rect 15932 23100 15988 23102
rect 14924 22652 14980 22708
rect 15036 22146 15092 22148
rect 15036 22094 15038 22146
rect 15038 22094 15090 22146
rect 15090 22094 15092 22146
rect 15036 22092 15092 22094
rect 15260 22652 15316 22708
rect 15932 22540 15988 22596
rect 15932 22258 15988 22260
rect 15932 22206 15934 22258
rect 15934 22206 15986 22258
rect 15986 22206 15988 22258
rect 15932 22204 15988 22206
rect 16268 22428 16324 22484
rect 15518 21978 15574 21980
rect 15518 21926 15520 21978
rect 15520 21926 15572 21978
rect 15572 21926 15574 21978
rect 15518 21924 15574 21926
rect 15622 21978 15678 21980
rect 15622 21926 15624 21978
rect 15624 21926 15676 21978
rect 15676 21926 15678 21978
rect 15622 21924 15678 21926
rect 15726 21978 15782 21980
rect 15726 21926 15728 21978
rect 15728 21926 15780 21978
rect 15780 21926 15782 21978
rect 15726 21924 15782 21926
rect 15372 21644 15428 21700
rect 15596 21698 15652 21700
rect 15596 21646 15598 21698
rect 15598 21646 15650 21698
rect 15650 21646 15652 21698
rect 15596 21644 15652 21646
rect 16044 21698 16100 21700
rect 16044 21646 16046 21698
rect 16046 21646 16098 21698
rect 16098 21646 16100 21698
rect 16044 21644 16100 21646
rect 15484 21532 15540 21588
rect 15036 21308 15092 21364
rect 15484 21196 15540 21252
rect 14924 20636 14980 20692
rect 14924 20300 14980 20356
rect 13692 19906 13748 19908
rect 13692 19854 13694 19906
rect 13694 19854 13746 19906
rect 13746 19854 13748 19906
rect 13692 19852 13748 19854
rect 14588 19852 14644 19908
rect 13468 19740 13524 19796
rect 13804 18956 13860 19012
rect 14364 19010 14420 19012
rect 14364 18958 14366 19010
rect 14366 18958 14418 19010
rect 14418 18958 14420 19010
rect 14364 18956 14420 18958
rect 13244 18396 13300 18452
rect 12236 15986 12292 15988
rect 12236 15934 12238 15986
rect 12238 15934 12290 15986
rect 12290 15934 12292 15986
rect 12236 15932 12292 15934
rect 12124 15092 12180 15148
rect 12124 14530 12180 14532
rect 12124 14478 12126 14530
rect 12126 14478 12178 14530
rect 12178 14478 12180 14530
rect 12124 14476 12180 14478
rect 12124 13244 12180 13300
rect 11900 12348 11956 12404
rect 12348 15148 12404 15204
rect 12572 16098 12628 16100
rect 12572 16046 12574 16098
rect 12574 16046 12626 16098
rect 12626 16046 12628 16098
rect 12572 16044 12628 16046
rect 13020 17612 13076 17668
rect 13468 18060 13524 18116
rect 13356 17724 13412 17780
rect 13580 17554 13636 17556
rect 13580 17502 13582 17554
rect 13582 17502 13634 17554
rect 13634 17502 13636 17554
rect 13580 17500 13636 17502
rect 13356 17106 13412 17108
rect 13356 17054 13358 17106
rect 13358 17054 13410 17106
rect 13410 17054 13412 17106
rect 13356 17052 13412 17054
rect 13132 16828 13188 16884
rect 12684 15484 12740 15540
rect 13244 16940 13300 16996
rect 12684 15036 12740 15092
rect 12572 14418 12628 14420
rect 12572 14366 12574 14418
rect 12574 14366 12626 14418
rect 12626 14366 12628 14418
rect 12572 14364 12628 14366
rect 12460 13356 12516 13412
rect 12796 13746 12852 13748
rect 12796 13694 12798 13746
rect 12798 13694 12850 13746
rect 12850 13694 12852 13746
rect 12796 13692 12852 13694
rect 13804 16940 13860 16996
rect 14812 17948 14868 18004
rect 15036 17836 15092 17892
rect 14028 17666 14084 17668
rect 14028 17614 14030 17666
rect 14030 17614 14082 17666
rect 14082 17614 14084 17666
rect 14028 17612 14084 17614
rect 14252 17500 14308 17556
rect 14028 17388 14084 17444
rect 14476 17052 14532 17108
rect 14700 16882 14756 16884
rect 14700 16830 14702 16882
rect 14702 16830 14754 16882
rect 14754 16830 14756 16882
rect 14700 16828 14756 16830
rect 16716 25340 16772 25396
rect 16604 23324 16660 23380
rect 16716 21980 16772 22036
rect 16380 21196 16436 21252
rect 16492 21644 16548 21700
rect 16268 21084 16324 21140
rect 16156 20860 16212 20916
rect 16268 20802 16324 20804
rect 16268 20750 16270 20802
rect 16270 20750 16322 20802
rect 16322 20750 16324 20802
rect 16268 20748 16324 20750
rect 15932 20690 15988 20692
rect 15932 20638 15934 20690
rect 15934 20638 15986 20690
rect 15986 20638 15988 20690
rect 15932 20636 15988 20638
rect 15518 20410 15574 20412
rect 15518 20358 15520 20410
rect 15520 20358 15572 20410
rect 15572 20358 15574 20410
rect 15518 20356 15574 20358
rect 15622 20410 15678 20412
rect 15622 20358 15624 20410
rect 15624 20358 15676 20410
rect 15676 20358 15678 20410
rect 15622 20356 15678 20358
rect 15726 20410 15782 20412
rect 15726 20358 15728 20410
rect 15728 20358 15780 20410
rect 15780 20358 15782 20410
rect 15726 20356 15782 20358
rect 15932 20188 15988 20244
rect 15820 19122 15876 19124
rect 15820 19070 15822 19122
rect 15822 19070 15874 19122
rect 15874 19070 15876 19122
rect 15820 19068 15876 19070
rect 15484 19010 15540 19012
rect 15484 18958 15486 19010
rect 15486 18958 15538 19010
rect 15538 18958 15540 19010
rect 15484 18956 15540 18958
rect 15932 19010 15988 19012
rect 15932 18958 15934 19010
rect 15934 18958 15986 19010
rect 15986 18958 15988 19010
rect 15932 18956 15988 18958
rect 15518 18842 15574 18844
rect 15518 18790 15520 18842
rect 15520 18790 15572 18842
rect 15572 18790 15574 18842
rect 15518 18788 15574 18790
rect 15622 18842 15678 18844
rect 15622 18790 15624 18842
rect 15624 18790 15676 18842
rect 15676 18790 15678 18842
rect 15622 18788 15678 18790
rect 15726 18842 15782 18844
rect 15726 18790 15728 18842
rect 15728 18790 15780 18842
rect 15780 18790 15782 18842
rect 15726 18788 15782 18790
rect 15260 17948 15316 18004
rect 15260 17554 15316 17556
rect 15260 17502 15262 17554
rect 15262 17502 15314 17554
rect 15314 17502 15316 17554
rect 15260 17500 15316 17502
rect 15260 16994 15316 16996
rect 15260 16942 15262 16994
rect 15262 16942 15314 16994
rect 15314 16942 15316 16994
rect 15260 16940 15316 16942
rect 16604 21586 16660 21588
rect 16604 21534 16606 21586
rect 16606 21534 16658 21586
rect 16658 21534 16660 21586
rect 16604 21532 16660 21534
rect 16604 20802 16660 20804
rect 16604 20750 16606 20802
rect 16606 20750 16658 20802
rect 16658 20750 16660 20802
rect 16604 20748 16660 20750
rect 16716 19964 16772 20020
rect 15518 17274 15574 17276
rect 15518 17222 15520 17274
rect 15520 17222 15572 17274
rect 15572 17222 15574 17274
rect 15518 17220 15574 17222
rect 15622 17274 15678 17276
rect 15622 17222 15624 17274
rect 15624 17222 15676 17274
rect 15676 17222 15678 17274
rect 15622 17220 15678 17222
rect 15726 17274 15782 17276
rect 15726 17222 15728 17274
rect 15728 17222 15780 17274
rect 15780 17222 15782 17274
rect 16044 17276 16100 17332
rect 15726 17220 15782 17222
rect 15372 16828 15428 16884
rect 15708 16994 15764 16996
rect 15708 16942 15710 16994
rect 15710 16942 15762 16994
rect 15762 16942 15764 16994
rect 15708 16940 15764 16942
rect 14028 16716 14084 16772
rect 14812 16716 14868 16772
rect 14364 16210 14420 16212
rect 14364 16158 14366 16210
rect 14366 16158 14418 16210
rect 14418 16158 14420 16210
rect 14364 16156 14420 16158
rect 14028 15932 14084 15988
rect 13804 15202 13860 15204
rect 13804 15150 13806 15202
rect 13806 15150 13858 15202
rect 13858 15150 13860 15202
rect 13804 15148 13860 15150
rect 13692 14306 13748 14308
rect 13692 14254 13694 14306
rect 13694 14254 13746 14306
rect 13746 14254 13748 14306
rect 13692 14252 13748 14254
rect 13356 13858 13412 13860
rect 13356 13806 13358 13858
rect 13358 13806 13410 13858
rect 13410 13806 13412 13858
rect 13356 13804 13412 13806
rect 12572 13244 12628 13300
rect 12572 12348 12628 12404
rect 11564 11788 11620 11844
rect 12348 11788 12404 11844
rect 11004 10498 11060 10500
rect 11004 10446 11006 10498
rect 11006 10446 11058 10498
rect 11058 10446 11060 10498
rect 11004 10444 11060 10446
rect 12348 11394 12404 11396
rect 12348 11342 12350 11394
rect 12350 11342 12402 11394
rect 12402 11342 12404 11394
rect 12348 11340 12404 11342
rect 13020 12738 13076 12740
rect 13020 12686 13022 12738
rect 13022 12686 13074 12738
rect 13074 12686 13076 12738
rect 13020 12684 13076 12686
rect 13468 12572 13524 12628
rect 11004 10050 11060 10052
rect 11004 9998 11006 10050
rect 11006 9998 11058 10050
rect 11058 9998 11060 10050
rect 11004 9996 11060 9998
rect 11004 9548 11060 9604
rect 10780 7980 10836 8036
rect 10780 6636 10836 6692
rect 11228 8876 11284 8932
rect 10780 6300 10836 6356
rect 10444 6018 10500 6020
rect 10444 5966 10446 6018
rect 10446 5966 10498 6018
rect 10498 5966 10500 6018
rect 10444 5964 10500 5966
rect 10108 5292 10164 5348
rect 8988 5180 9044 5236
rect 9212 5234 9268 5236
rect 9212 5182 9214 5234
rect 9214 5182 9266 5234
rect 9266 5182 9268 5234
rect 9212 5180 9268 5182
rect 9772 5180 9828 5236
rect 8204 5068 8260 5124
rect 9548 5122 9604 5124
rect 9548 5070 9550 5122
rect 9550 5070 9602 5122
rect 9602 5070 9604 5122
rect 9548 5068 9604 5070
rect 8092 4844 8148 4900
rect 8988 4562 9044 4564
rect 8988 4510 8990 4562
rect 8990 4510 9042 4562
rect 9042 4510 9044 4562
rect 8988 4508 9044 4510
rect 10444 5180 10500 5236
rect 8428 4060 8484 4116
rect 8365 3946 8421 3948
rect 8365 3894 8367 3946
rect 8367 3894 8419 3946
rect 8419 3894 8421 3946
rect 8365 3892 8421 3894
rect 8469 3946 8525 3948
rect 8469 3894 8471 3946
rect 8471 3894 8523 3946
rect 8523 3894 8525 3946
rect 8469 3892 8525 3894
rect 8573 3946 8629 3948
rect 8573 3894 8575 3946
rect 8575 3894 8627 3946
rect 8627 3894 8629 3946
rect 8573 3892 8629 3894
rect 10780 5122 10836 5124
rect 10780 5070 10782 5122
rect 10782 5070 10834 5122
rect 10834 5070 10836 5122
rect 10780 5068 10836 5070
rect 11228 6524 11284 6580
rect 13692 13746 13748 13748
rect 13692 13694 13694 13746
rect 13694 13694 13746 13746
rect 13746 13694 13748 13746
rect 13692 13692 13748 13694
rect 13804 13244 13860 13300
rect 14588 15148 14644 15204
rect 14028 15036 14084 15092
rect 16268 17388 16324 17444
rect 14924 15932 14980 15988
rect 15932 16828 15988 16884
rect 15518 15706 15574 15708
rect 15518 15654 15520 15706
rect 15520 15654 15572 15706
rect 15572 15654 15574 15706
rect 15518 15652 15574 15654
rect 15622 15706 15678 15708
rect 15622 15654 15624 15706
rect 15624 15654 15676 15706
rect 15676 15654 15678 15706
rect 15622 15652 15678 15654
rect 15726 15706 15782 15708
rect 15726 15654 15728 15706
rect 15728 15654 15780 15706
rect 15780 15654 15782 15706
rect 15726 15652 15782 15654
rect 15484 15538 15540 15540
rect 15484 15486 15486 15538
rect 15486 15486 15538 15538
rect 15538 15486 15540 15538
rect 15484 15484 15540 15486
rect 16268 16882 16324 16884
rect 16268 16830 16270 16882
rect 16270 16830 16322 16882
rect 16322 16830 16324 16882
rect 16268 16828 16324 16830
rect 16492 18956 16548 19012
rect 16828 18732 16884 18788
rect 16604 17890 16660 17892
rect 16604 17838 16606 17890
rect 16606 17838 16658 17890
rect 16658 17838 16660 17890
rect 16604 17836 16660 17838
rect 16716 17724 16772 17780
rect 16492 17554 16548 17556
rect 16492 17502 16494 17554
rect 16494 17502 16546 17554
rect 16546 17502 16548 17554
rect 16492 17500 16548 17502
rect 17052 31778 17108 31780
rect 17052 31726 17054 31778
rect 17054 31726 17106 31778
rect 17106 31726 17108 31778
rect 17052 31724 17108 31726
rect 17388 31388 17444 31444
rect 17948 31554 18004 31556
rect 17948 31502 17950 31554
rect 17950 31502 18002 31554
rect 18002 31502 18004 31554
rect 17948 31500 18004 31502
rect 18060 31388 18116 31444
rect 17052 30156 17108 30212
rect 17052 29986 17108 29988
rect 17052 29934 17054 29986
rect 17054 29934 17106 29986
rect 17106 29934 17108 29986
rect 17052 29932 17108 29934
rect 17612 29932 17668 29988
rect 17276 27186 17332 27188
rect 17276 27134 17278 27186
rect 17278 27134 17330 27186
rect 17330 27134 17332 27186
rect 17276 27132 17332 27134
rect 16940 18284 16996 18340
rect 16604 16882 16660 16884
rect 16604 16830 16606 16882
rect 16606 16830 16658 16882
rect 16658 16830 16660 16882
rect 16604 16828 16660 16830
rect 15036 15314 15092 15316
rect 15036 15262 15038 15314
rect 15038 15262 15090 15314
rect 15090 15262 15092 15314
rect 15036 15260 15092 15262
rect 14924 15148 14980 15204
rect 14700 15036 14756 15092
rect 14588 14642 14644 14644
rect 14588 14590 14590 14642
rect 14590 14590 14642 14642
rect 14642 14590 14644 14642
rect 14588 14588 14644 14590
rect 14700 14476 14756 14532
rect 14140 14418 14196 14420
rect 14140 14366 14142 14418
rect 14142 14366 14194 14418
rect 14194 14366 14196 14418
rect 14140 14364 14196 14366
rect 15036 14418 15092 14420
rect 15036 14366 15038 14418
rect 15038 14366 15090 14418
rect 15090 14366 15092 14418
rect 15036 14364 15092 14366
rect 15260 14418 15316 14420
rect 15260 14366 15262 14418
rect 15262 14366 15314 14418
rect 15314 14366 15316 14418
rect 15260 14364 15316 14366
rect 15148 13692 15204 13748
rect 16380 15538 16436 15540
rect 16380 15486 16382 15538
rect 16382 15486 16434 15538
rect 16434 15486 16436 15538
rect 16380 15484 16436 15486
rect 15932 14588 15988 14644
rect 15932 14418 15988 14420
rect 15932 14366 15934 14418
rect 15934 14366 15986 14418
rect 15986 14366 15988 14418
rect 15932 14364 15988 14366
rect 15518 14138 15574 14140
rect 15518 14086 15520 14138
rect 15520 14086 15572 14138
rect 15572 14086 15574 14138
rect 15518 14084 15574 14086
rect 15622 14138 15678 14140
rect 15622 14086 15624 14138
rect 15624 14086 15676 14138
rect 15676 14086 15678 14138
rect 15622 14084 15678 14086
rect 15726 14138 15782 14140
rect 15726 14086 15728 14138
rect 15728 14086 15780 14138
rect 15780 14086 15782 14138
rect 15726 14084 15782 14086
rect 14700 13580 14756 13636
rect 14364 13468 14420 13524
rect 17500 26124 17556 26180
rect 17164 25618 17220 25620
rect 17164 25566 17166 25618
rect 17166 25566 17218 25618
rect 17218 25566 17220 25618
rect 17164 25564 17220 25566
rect 17388 23714 17444 23716
rect 17388 23662 17390 23714
rect 17390 23662 17442 23714
rect 17442 23662 17444 23714
rect 17388 23660 17444 23662
rect 17388 23154 17444 23156
rect 17388 23102 17390 23154
rect 17390 23102 17442 23154
rect 17442 23102 17444 23154
rect 17388 23100 17444 23102
rect 17500 21698 17556 21700
rect 17500 21646 17502 21698
rect 17502 21646 17554 21698
rect 17554 21646 17556 21698
rect 17500 21644 17556 21646
rect 17388 20914 17444 20916
rect 17388 20862 17390 20914
rect 17390 20862 17442 20914
rect 17442 20862 17444 20914
rect 17388 20860 17444 20862
rect 17500 20188 17556 20244
rect 19068 34524 19124 34580
rect 18956 34130 19012 34132
rect 18956 34078 18958 34130
rect 18958 34078 19010 34130
rect 19010 34078 19012 34130
rect 18956 34076 19012 34078
rect 18284 33740 18340 33796
rect 18732 33404 18788 33460
rect 18844 33852 18900 33908
rect 18508 32508 18564 32564
rect 18732 32396 18788 32452
rect 18284 31778 18340 31780
rect 18284 31726 18286 31778
rect 18286 31726 18338 31778
rect 18338 31726 18340 31778
rect 18284 31724 18340 31726
rect 20300 34748 20356 34804
rect 20524 34636 20580 34692
rect 25004 36482 25060 36484
rect 25004 36430 25006 36482
rect 25006 36430 25058 36482
rect 25058 36430 25060 36482
rect 25004 36428 25060 36430
rect 21308 35980 21364 36036
rect 21644 35922 21700 35924
rect 21644 35870 21646 35922
rect 21646 35870 21698 35922
rect 21698 35870 21700 35922
rect 21644 35868 21700 35870
rect 20972 34524 21028 34580
rect 21420 34972 21476 35028
rect 21644 35644 21700 35700
rect 22764 35980 22820 36036
rect 22876 35868 22932 35924
rect 22428 35084 22484 35140
rect 22316 34972 22372 35028
rect 21420 34802 21476 34804
rect 21420 34750 21422 34802
rect 21422 34750 21474 34802
rect 21474 34750 21476 34802
rect 21420 34748 21476 34750
rect 21308 34524 21364 34580
rect 19628 34188 19684 34244
rect 19516 33852 19572 33908
rect 19852 33740 19908 33796
rect 20188 33404 20244 33460
rect 20524 33852 20580 33908
rect 21756 34860 21812 34916
rect 22092 34242 22148 34244
rect 22092 34190 22094 34242
rect 22094 34190 22146 34242
rect 22146 34190 22148 34242
rect 22092 34188 22148 34190
rect 21980 33628 22036 33684
rect 21980 33458 22036 33460
rect 21980 33406 21982 33458
rect 21982 33406 22034 33458
rect 22034 33406 22036 33458
rect 21980 33404 22036 33406
rect 19852 33068 19908 33124
rect 19516 32956 19572 33012
rect 19516 32450 19572 32452
rect 19516 32398 19518 32450
rect 19518 32398 19570 32450
rect 19570 32398 19572 32450
rect 19516 32396 19572 32398
rect 18956 31500 19012 31556
rect 19404 31218 19460 31220
rect 19404 31166 19406 31218
rect 19406 31166 19458 31218
rect 19458 31166 19460 31218
rect 19404 31164 19460 31166
rect 18620 30380 18676 30436
rect 18396 30268 18452 30324
rect 18844 30210 18900 30212
rect 18844 30158 18846 30210
rect 18846 30158 18898 30210
rect 18898 30158 18900 30210
rect 18844 30156 18900 30158
rect 18172 29820 18228 29876
rect 19404 29820 19460 29876
rect 18172 28924 18228 28980
rect 19068 28924 19124 28980
rect 17724 28588 17780 28644
rect 18844 28642 18900 28644
rect 18844 28590 18846 28642
rect 18846 28590 18898 28642
rect 18898 28590 18900 28642
rect 18844 28588 18900 28590
rect 18508 28140 18564 28196
rect 18060 27468 18116 27524
rect 18620 27970 18676 27972
rect 18620 27918 18622 27970
rect 18622 27918 18674 27970
rect 18674 27918 18676 27970
rect 18620 27916 18676 27918
rect 18284 27858 18340 27860
rect 18284 27806 18286 27858
rect 18286 27806 18338 27858
rect 18338 27806 18340 27858
rect 18284 27804 18340 27806
rect 18956 27746 19012 27748
rect 18956 27694 18958 27746
rect 18958 27694 19010 27746
rect 19010 27694 19012 27746
rect 18956 27692 19012 27694
rect 18172 27132 18228 27188
rect 19180 27356 19236 27412
rect 18620 27074 18676 27076
rect 18620 27022 18622 27074
rect 18622 27022 18674 27074
rect 18674 27022 18676 27074
rect 18620 27020 18676 27022
rect 18844 26796 18900 26852
rect 17948 26572 18004 26628
rect 17724 24050 17780 24052
rect 17724 23998 17726 24050
rect 17726 23998 17778 24050
rect 17778 23998 17780 24050
rect 17724 23996 17780 23998
rect 18284 24892 18340 24948
rect 19180 24892 19236 24948
rect 18284 24444 18340 24500
rect 18508 23996 18564 24052
rect 18172 22092 18228 22148
rect 18956 22204 19012 22260
rect 17836 21756 17892 21812
rect 18508 21698 18564 21700
rect 18508 21646 18510 21698
rect 18510 21646 18562 21698
rect 18562 21646 18564 21698
rect 18508 21644 18564 21646
rect 18396 21362 18452 21364
rect 18396 21310 18398 21362
rect 18398 21310 18450 21362
rect 18450 21310 18452 21362
rect 18396 21308 18452 21310
rect 18060 20300 18116 20356
rect 19068 21698 19124 21700
rect 19068 21646 19070 21698
rect 19070 21646 19122 21698
rect 19122 21646 19124 21698
rect 19068 21644 19124 21646
rect 18956 20972 19012 21028
rect 19180 21196 19236 21252
rect 18508 20412 18564 20468
rect 18172 20188 18228 20244
rect 17612 20076 17668 20132
rect 19740 29426 19796 29428
rect 19740 29374 19742 29426
rect 19742 29374 19794 29426
rect 19794 29374 19796 29426
rect 19740 29372 19796 29374
rect 22428 34636 22484 34692
rect 22652 35698 22708 35700
rect 22652 35646 22654 35698
rect 22654 35646 22706 35698
rect 22706 35646 22708 35698
rect 22652 35644 22708 35646
rect 22876 35644 22932 35700
rect 24668 36258 24724 36260
rect 24668 36206 24670 36258
rect 24670 36206 24722 36258
rect 24722 36206 24724 36258
rect 24668 36204 24724 36206
rect 24220 35532 24276 35588
rect 24332 35980 24388 36036
rect 22672 35306 22728 35308
rect 22672 35254 22674 35306
rect 22674 35254 22726 35306
rect 22726 35254 22728 35306
rect 22672 35252 22728 35254
rect 22776 35306 22832 35308
rect 22776 35254 22778 35306
rect 22778 35254 22830 35306
rect 22830 35254 22832 35306
rect 22776 35252 22832 35254
rect 22880 35306 22936 35308
rect 22880 35254 22882 35306
rect 22882 35254 22934 35306
rect 22934 35254 22936 35306
rect 22880 35252 22936 35254
rect 23996 35084 24052 35140
rect 22540 34748 22596 34804
rect 22540 34188 22596 34244
rect 23436 34802 23492 34804
rect 23436 34750 23438 34802
rect 23438 34750 23490 34802
rect 23490 34750 23492 34802
rect 23436 34748 23492 34750
rect 24220 34636 24276 34692
rect 26684 36258 26740 36260
rect 26684 36206 26686 36258
rect 26686 36206 26738 36258
rect 26738 36206 26740 36258
rect 26684 36204 26740 36206
rect 24668 35644 24724 35700
rect 24556 35474 24612 35476
rect 24556 35422 24558 35474
rect 24558 35422 24610 35474
rect 24610 35422 24612 35474
rect 24556 35420 24612 35422
rect 24444 35084 24500 35140
rect 26012 35698 26068 35700
rect 26012 35646 26014 35698
rect 26014 35646 26066 35698
rect 26066 35646 26068 35698
rect 26012 35644 26068 35646
rect 26684 35644 26740 35700
rect 25676 35586 25732 35588
rect 25676 35534 25678 35586
rect 25678 35534 25730 35586
rect 25730 35534 25732 35586
rect 25676 35532 25732 35534
rect 22764 33852 22820 33908
rect 22672 33738 22728 33740
rect 22672 33686 22674 33738
rect 22674 33686 22726 33738
rect 22726 33686 22728 33738
rect 22672 33684 22728 33686
rect 22776 33738 22832 33740
rect 22776 33686 22778 33738
rect 22778 33686 22830 33738
rect 22830 33686 22832 33738
rect 22776 33684 22832 33686
rect 22880 33738 22936 33740
rect 22880 33686 22882 33738
rect 22882 33686 22934 33738
rect 22934 33686 22936 33738
rect 22880 33684 22936 33686
rect 20188 32956 20244 33012
rect 21420 32732 21476 32788
rect 21532 32956 21588 33012
rect 20188 31500 20244 31556
rect 20300 31388 20356 31444
rect 20860 30716 20916 30772
rect 19964 30434 20020 30436
rect 19964 30382 19966 30434
rect 19966 30382 20018 30434
rect 20018 30382 20020 30434
rect 19964 30380 20020 30382
rect 20188 30156 20244 30212
rect 20860 29708 20916 29764
rect 21868 32844 21924 32900
rect 21756 32674 21812 32676
rect 21756 32622 21758 32674
rect 21758 32622 21810 32674
rect 21810 32622 21812 32674
rect 21756 32620 21812 32622
rect 21532 31724 21588 31780
rect 21644 31164 21700 31220
rect 21532 30322 21588 30324
rect 21532 30270 21534 30322
rect 21534 30270 21586 30322
rect 21586 30270 21588 30322
rect 21532 30268 21588 30270
rect 20748 29650 20804 29652
rect 20748 29598 20750 29650
rect 20750 29598 20802 29650
rect 20802 29598 20804 29650
rect 20748 29596 20804 29598
rect 19404 27858 19460 27860
rect 19404 27806 19406 27858
rect 19406 27806 19458 27858
rect 19458 27806 19460 27858
rect 19404 27804 19460 27806
rect 19740 28476 19796 28532
rect 19852 27746 19908 27748
rect 19852 27694 19854 27746
rect 19854 27694 19906 27746
rect 19906 27694 19908 27746
rect 19852 27692 19908 27694
rect 19516 27020 19572 27076
rect 19628 26796 19684 26852
rect 19628 26236 19684 26292
rect 19628 24722 19684 24724
rect 19628 24670 19630 24722
rect 19630 24670 19682 24722
rect 19682 24670 19684 24722
rect 19628 24668 19684 24670
rect 19740 24444 19796 24500
rect 19628 24050 19684 24052
rect 19628 23998 19630 24050
rect 19630 23998 19682 24050
rect 19682 23998 19684 24050
rect 19628 23996 19684 23998
rect 19740 23660 19796 23716
rect 19404 22258 19460 22260
rect 19404 22206 19406 22258
rect 19406 22206 19458 22258
rect 19458 22206 19460 22258
rect 19404 22204 19460 22206
rect 19516 20972 19572 21028
rect 20076 28924 20132 28980
rect 21196 29596 21252 29652
rect 20188 28700 20244 28756
rect 21308 29260 21364 29316
rect 20636 28924 20692 28980
rect 20524 28476 20580 28532
rect 20188 27916 20244 27972
rect 20076 27804 20132 27860
rect 20412 27746 20468 27748
rect 20412 27694 20414 27746
rect 20414 27694 20466 27746
rect 20466 27694 20468 27746
rect 20412 27692 20468 27694
rect 20300 27356 20356 27412
rect 21868 29932 21924 29988
rect 21868 29708 21924 29764
rect 21756 29596 21812 29652
rect 22316 29260 22372 29316
rect 23324 34018 23380 34020
rect 23324 33966 23326 34018
rect 23326 33966 23378 34018
rect 23378 33966 23380 34018
rect 23324 33964 23380 33966
rect 23996 33852 24052 33908
rect 23100 32844 23156 32900
rect 24444 33740 24500 33796
rect 23884 32844 23940 32900
rect 22672 32170 22728 32172
rect 22672 32118 22674 32170
rect 22674 32118 22726 32170
rect 22726 32118 22728 32170
rect 22672 32116 22728 32118
rect 22776 32170 22832 32172
rect 22776 32118 22778 32170
rect 22778 32118 22830 32170
rect 22830 32118 22832 32170
rect 22776 32116 22832 32118
rect 22880 32170 22936 32172
rect 22880 32118 22882 32170
rect 22882 32118 22934 32170
rect 22934 32118 22936 32170
rect 22880 32116 22936 32118
rect 24332 31948 24388 32004
rect 22428 30716 22484 30772
rect 21980 28700 22036 28756
rect 20860 27858 20916 27860
rect 20860 27806 20862 27858
rect 20862 27806 20914 27858
rect 20914 27806 20916 27858
rect 20860 27804 20916 27806
rect 21420 28418 21476 28420
rect 21420 28366 21422 28418
rect 21422 28366 21474 28418
rect 21474 28366 21476 28418
rect 21420 28364 21476 28366
rect 22092 28530 22148 28532
rect 22092 28478 22094 28530
rect 22094 28478 22146 28530
rect 22146 28478 22148 28530
rect 22092 28476 22148 28478
rect 22316 28364 22372 28420
rect 22316 27692 22372 27748
rect 22092 27244 22148 27300
rect 20188 26572 20244 26628
rect 20300 26290 20356 26292
rect 20300 26238 20302 26290
rect 20302 26238 20354 26290
rect 20354 26238 20356 26290
rect 20300 26236 20356 26238
rect 20300 23660 20356 23716
rect 19964 21196 20020 21252
rect 20076 22092 20132 22148
rect 19740 20860 19796 20916
rect 19516 20300 19572 20356
rect 19292 20242 19348 20244
rect 19292 20190 19294 20242
rect 19294 20190 19346 20242
rect 19346 20190 19348 20242
rect 19292 20188 19348 20190
rect 18956 19852 19012 19908
rect 17836 19794 17892 19796
rect 17836 19742 17838 19794
rect 17838 19742 17890 19794
rect 17890 19742 17892 19794
rect 17836 19740 17892 19742
rect 17052 16828 17108 16884
rect 17164 19292 17220 19348
rect 17276 19234 17332 19236
rect 17276 19182 17278 19234
rect 17278 19182 17330 19234
rect 17330 19182 17332 19234
rect 17276 19180 17332 19182
rect 17164 18956 17220 19012
rect 17612 19122 17668 19124
rect 17612 19070 17614 19122
rect 17614 19070 17666 19122
rect 17666 19070 17668 19122
rect 17612 19068 17668 19070
rect 17500 18732 17556 18788
rect 17724 19010 17780 19012
rect 17724 18958 17726 19010
rect 17726 18958 17778 19010
rect 17778 18958 17780 19010
rect 17724 18956 17780 18958
rect 16940 15932 16996 15988
rect 17948 18450 18004 18452
rect 17948 18398 17950 18450
rect 17950 18398 18002 18450
rect 18002 18398 18004 18450
rect 17948 18396 18004 18398
rect 18060 18284 18116 18340
rect 18060 17442 18116 17444
rect 18060 17390 18062 17442
rect 18062 17390 18114 17442
rect 18114 17390 18116 17442
rect 18060 17388 18116 17390
rect 17836 16940 17892 16996
rect 18172 17052 18228 17108
rect 17164 15484 17220 15540
rect 16716 15372 16772 15428
rect 16268 14418 16324 14420
rect 16268 14366 16270 14418
rect 16270 14366 16322 14418
rect 16322 14366 16324 14418
rect 16268 14364 16324 14366
rect 16380 14306 16436 14308
rect 16380 14254 16382 14306
rect 16382 14254 16434 14306
rect 16434 14254 16436 14306
rect 16380 14252 16436 14254
rect 16156 14140 16212 14196
rect 15372 13132 15428 13188
rect 14252 12738 14308 12740
rect 14252 12686 14254 12738
rect 14254 12686 14306 12738
rect 14306 12686 14308 12738
rect 14252 12684 14308 12686
rect 14140 11564 14196 11620
rect 14364 11676 14420 11732
rect 14364 11394 14420 11396
rect 14364 11342 14366 11394
rect 14366 11342 14418 11394
rect 14418 11342 14420 11394
rect 14364 11340 14420 11342
rect 12012 9602 12068 9604
rect 12012 9550 12014 9602
rect 12014 9550 12066 9602
rect 12066 9550 12068 9602
rect 12012 9548 12068 9550
rect 12460 8428 12516 8484
rect 11900 8204 11956 8260
rect 11116 6076 11172 6132
rect 11228 6018 11284 6020
rect 11228 5966 11230 6018
rect 11230 5966 11282 6018
rect 11282 5966 11284 6018
rect 11228 5964 11284 5966
rect 11116 5852 11172 5908
rect 11004 4844 11060 4900
rect 10668 4396 10724 4452
rect 10892 3948 10948 4004
rect 10556 3724 10612 3780
rect 8092 3388 8148 3444
rect 7756 3276 7812 3332
rect 8876 3442 8932 3444
rect 8876 3390 8878 3442
rect 8878 3390 8930 3442
rect 8930 3390 8932 3442
rect 8876 3388 8932 3390
rect 11340 5010 11396 5012
rect 11340 4958 11342 5010
rect 11342 4958 11394 5010
rect 11394 4958 11396 5010
rect 11340 4956 11396 4958
rect 11340 4732 11396 4788
rect 11452 4338 11508 4340
rect 11452 4286 11454 4338
rect 11454 4286 11506 4338
rect 11506 4286 11508 4338
rect 11452 4284 11508 4286
rect 11452 4060 11508 4116
rect 11564 3948 11620 4004
rect 11228 3388 11284 3444
rect 11228 2940 11284 2996
rect 11900 6018 11956 6020
rect 11900 5966 11902 6018
rect 11902 5966 11954 6018
rect 11954 5966 11956 6018
rect 11900 5964 11956 5966
rect 11788 4620 11844 4676
rect 12572 10108 12628 10164
rect 12796 9938 12852 9940
rect 12796 9886 12798 9938
rect 12798 9886 12850 9938
rect 12850 9886 12852 9938
rect 12796 9884 12852 9886
rect 13132 8988 13188 9044
rect 13020 8764 13076 8820
rect 13356 8316 13412 8372
rect 12684 8146 12740 8148
rect 12684 8094 12686 8146
rect 12686 8094 12738 8146
rect 12738 8094 12740 8146
rect 12684 8092 12740 8094
rect 12796 8034 12852 8036
rect 12796 7982 12798 8034
rect 12798 7982 12850 8034
rect 12850 7982 12852 8034
rect 12796 7980 12852 7982
rect 13356 7868 13412 7924
rect 12124 6690 12180 6692
rect 12124 6638 12126 6690
rect 12126 6638 12178 6690
rect 12178 6638 12180 6690
rect 12124 6636 12180 6638
rect 14812 12012 14868 12068
rect 15596 12850 15652 12852
rect 15596 12798 15598 12850
rect 15598 12798 15650 12850
rect 15650 12798 15652 12850
rect 15596 12796 15652 12798
rect 15820 13356 15876 13412
rect 16268 13692 16324 13748
rect 16156 13020 16212 13076
rect 16380 13356 16436 13412
rect 16604 13916 16660 13972
rect 16604 13746 16660 13748
rect 16604 13694 16606 13746
rect 16606 13694 16658 13746
rect 16658 13694 16660 13746
rect 16604 13692 16660 13694
rect 16604 13020 16660 13076
rect 15708 12684 15764 12740
rect 16492 12796 16548 12852
rect 15518 12570 15574 12572
rect 15518 12518 15520 12570
rect 15520 12518 15572 12570
rect 15572 12518 15574 12570
rect 15518 12516 15574 12518
rect 15622 12570 15678 12572
rect 15622 12518 15624 12570
rect 15624 12518 15676 12570
rect 15676 12518 15678 12570
rect 15622 12516 15678 12518
rect 15726 12570 15782 12572
rect 15726 12518 15728 12570
rect 15728 12518 15780 12570
rect 15780 12518 15782 12570
rect 15726 12516 15782 12518
rect 16492 12572 16548 12628
rect 15820 12348 15876 12404
rect 15596 12290 15652 12292
rect 15596 12238 15598 12290
rect 15598 12238 15650 12290
rect 15650 12238 15652 12290
rect 15596 12236 15652 12238
rect 15260 12124 15316 12180
rect 16604 12066 16660 12068
rect 16604 12014 16606 12066
rect 16606 12014 16658 12066
rect 16658 12014 16660 12066
rect 16604 12012 16660 12014
rect 13580 10556 13636 10612
rect 15518 11002 15574 11004
rect 15518 10950 15520 11002
rect 15520 10950 15572 11002
rect 15572 10950 15574 11002
rect 15518 10948 15574 10950
rect 15622 11002 15678 11004
rect 15622 10950 15624 11002
rect 15624 10950 15676 11002
rect 15676 10950 15678 11002
rect 15622 10948 15678 10950
rect 15726 11002 15782 11004
rect 15726 10950 15728 11002
rect 15728 10950 15780 11002
rect 15780 10950 15782 11002
rect 15726 10948 15782 10950
rect 15932 10780 15988 10836
rect 13916 9884 13972 9940
rect 14476 10332 14532 10388
rect 14252 9548 14308 9604
rect 13916 9042 13972 9044
rect 13916 8990 13918 9042
rect 13918 8990 13970 9042
rect 13970 8990 13972 9042
rect 13916 8988 13972 8990
rect 14252 8652 14308 8708
rect 14364 10108 14420 10164
rect 13804 8540 13860 8596
rect 14700 8988 14756 9044
rect 15260 10498 15316 10500
rect 15260 10446 15262 10498
rect 15262 10446 15314 10498
rect 15314 10446 15316 10498
rect 15260 10444 15316 10446
rect 15036 9660 15092 9716
rect 16380 10834 16436 10836
rect 16380 10782 16382 10834
rect 16382 10782 16434 10834
rect 16434 10782 16436 10834
rect 16380 10780 16436 10782
rect 16380 10220 16436 10276
rect 16828 13468 16884 13524
rect 17052 14642 17108 14644
rect 17052 14590 17054 14642
rect 17054 14590 17106 14642
rect 17106 14590 17108 14642
rect 17052 14588 17108 14590
rect 18060 16828 18116 16884
rect 17724 16210 17780 16212
rect 17724 16158 17726 16210
rect 17726 16158 17778 16210
rect 17778 16158 17780 16210
rect 17724 16156 17780 16158
rect 17612 15538 17668 15540
rect 17612 15486 17614 15538
rect 17614 15486 17666 15538
rect 17666 15486 17668 15538
rect 17612 15484 17668 15486
rect 19180 19794 19236 19796
rect 19180 19742 19182 19794
rect 19182 19742 19234 19794
rect 19234 19742 19236 19794
rect 19180 19740 19236 19742
rect 18956 19180 19012 19236
rect 18732 19010 18788 19012
rect 18732 18958 18734 19010
rect 18734 18958 18786 19010
rect 18786 18958 18788 19010
rect 18732 18956 18788 18958
rect 19068 18732 19124 18788
rect 19404 18956 19460 19012
rect 19516 18844 19572 18900
rect 19740 20412 19796 20468
rect 19852 19516 19908 19572
rect 18620 16492 18676 16548
rect 18396 15820 18452 15876
rect 17724 15148 17780 15204
rect 18396 15372 18452 15428
rect 18620 15036 18676 15092
rect 18284 14476 18340 14532
rect 17612 14252 17668 14308
rect 17948 13580 18004 13636
rect 17500 13356 17556 13412
rect 17164 13074 17220 13076
rect 17164 13022 17166 13074
rect 17166 13022 17218 13074
rect 17218 13022 17220 13074
rect 17164 13020 17220 13022
rect 17612 12684 17668 12740
rect 16828 12124 16884 12180
rect 17388 12178 17444 12180
rect 17388 12126 17390 12178
rect 17390 12126 17442 12178
rect 17442 12126 17444 12178
rect 17388 12124 17444 12126
rect 16940 11676 16996 11732
rect 16940 11340 16996 11396
rect 16828 10220 16884 10276
rect 16380 9826 16436 9828
rect 16380 9774 16382 9826
rect 16382 9774 16434 9826
rect 16434 9774 16436 9826
rect 16380 9772 16436 9774
rect 15518 9434 15574 9436
rect 15518 9382 15520 9434
rect 15520 9382 15572 9434
rect 15572 9382 15574 9434
rect 15518 9380 15574 9382
rect 15622 9434 15678 9436
rect 15622 9382 15624 9434
rect 15624 9382 15676 9434
rect 15676 9382 15678 9434
rect 15622 9380 15678 9382
rect 15726 9434 15782 9436
rect 15726 9382 15728 9434
rect 15728 9382 15780 9434
rect 15780 9382 15782 9434
rect 15726 9380 15782 9382
rect 15484 8930 15540 8932
rect 15484 8878 15486 8930
rect 15486 8878 15538 8930
rect 15538 8878 15540 8930
rect 15484 8876 15540 8878
rect 15148 8764 15204 8820
rect 13692 8316 13748 8372
rect 13580 8258 13636 8260
rect 13580 8206 13582 8258
rect 13582 8206 13634 8258
rect 13634 8206 13636 8258
rect 13580 8204 13636 8206
rect 14028 8034 14084 8036
rect 14028 7982 14030 8034
rect 14030 7982 14082 8034
rect 14082 7982 14084 8034
rect 14028 7980 14084 7982
rect 14364 7868 14420 7924
rect 14476 7980 14532 8036
rect 14028 7586 14084 7588
rect 14028 7534 14030 7586
rect 14030 7534 14082 7586
rect 14082 7534 14084 7586
rect 14028 7532 14084 7534
rect 13468 6860 13524 6916
rect 12796 6748 12852 6804
rect 12124 5964 12180 6020
rect 12348 6018 12404 6020
rect 12348 5966 12350 6018
rect 12350 5966 12402 6018
rect 12402 5966 12404 6018
rect 12348 5964 12404 5966
rect 12572 5906 12628 5908
rect 12572 5854 12574 5906
rect 12574 5854 12626 5906
rect 12626 5854 12628 5906
rect 12572 5852 12628 5854
rect 12908 5964 12964 6020
rect 11900 4338 11956 4340
rect 11900 4286 11902 4338
rect 11902 4286 11954 4338
rect 11954 4286 11956 4338
rect 11900 4284 11956 4286
rect 13356 5906 13412 5908
rect 13356 5854 13358 5906
rect 13358 5854 13410 5906
rect 13410 5854 13412 5906
rect 13356 5852 13412 5854
rect 13132 5794 13188 5796
rect 13132 5742 13134 5794
rect 13134 5742 13186 5794
rect 13186 5742 13188 5794
rect 13132 5740 13188 5742
rect 13132 5404 13188 5460
rect 12908 5346 12964 5348
rect 12908 5294 12910 5346
rect 12910 5294 12962 5346
rect 12962 5294 12964 5346
rect 12908 5292 12964 5294
rect 12460 5234 12516 5236
rect 12460 5182 12462 5234
rect 12462 5182 12514 5234
rect 12514 5182 12516 5234
rect 12460 5180 12516 5182
rect 14924 8316 14980 8372
rect 14700 6748 14756 6804
rect 14476 6130 14532 6132
rect 14476 6078 14478 6130
rect 14478 6078 14530 6130
rect 14530 6078 14532 6130
rect 14476 6076 14532 6078
rect 15708 8204 15764 8260
rect 16044 8876 16100 8932
rect 15260 8146 15316 8148
rect 15260 8094 15262 8146
rect 15262 8094 15314 8146
rect 15314 8094 15316 8146
rect 15260 8092 15316 8094
rect 15596 8146 15652 8148
rect 15596 8094 15598 8146
rect 15598 8094 15650 8146
rect 15650 8094 15652 8146
rect 15596 8092 15652 8094
rect 15932 8146 15988 8148
rect 15932 8094 15934 8146
rect 15934 8094 15986 8146
rect 15986 8094 15988 8146
rect 15932 8092 15988 8094
rect 15036 7698 15092 7700
rect 15036 7646 15038 7698
rect 15038 7646 15090 7698
rect 15090 7646 15092 7698
rect 15036 7644 15092 7646
rect 15518 7866 15574 7868
rect 15518 7814 15520 7866
rect 15520 7814 15572 7866
rect 15572 7814 15574 7866
rect 15518 7812 15574 7814
rect 15622 7866 15678 7868
rect 15622 7814 15624 7866
rect 15624 7814 15676 7866
rect 15676 7814 15678 7866
rect 15622 7812 15678 7814
rect 15726 7866 15782 7868
rect 15726 7814 15728 7866
rect 15728 7814 15780 7866
rect 15780 7814 15782 7866
rect 15726 7812 15782 7814
rect 15372 7532 15428 7588
rect 15932 7532 15988 7588
rect 15260 7084 15316 7140
rect 15708 7250 15764 7252
rect 15708 7198 15710 7250
rect 15710 7198 15762 7250
rect 15762 7198 15764 7250
rect 15708 7196 15764 7198
rect 15372 6972 15428 7028
rect 14924 6300 14980 6356
rect 15148 6748 15204 6804
rect 15484 6748 15540 6804
rect 14812 6130 14868 6132
rect 14812 6078 14814 6130
rect 14814 6078 14866 6130
rect 14866 6078 14868 6130
rect 14812 6076 14868 6078
rect 12796 5010 12852 5012
rect 12796 4958 12798 5010
rect 12798 4958 12850 5010
rect 12850 4958 12852 5010
rect 12796 4956 12852 4958
rect 12684 4844 12740 4900
rect 12124 4450 12180 4452
rect 12124 4398 12126 4450
rect 12126 4398 12178 4450
rect 12178 4398 12180 4450
rect 12124 4396 12180 4398
rect 14028 5740 14084 5796
rect 14700 5516 14756 5572
rect 13580 4898 13636 4900
rect 13580 4846 13582 4898
rect 13582 4846 13634 4898
rect 13634 4846 13636 4898
rect 13580 4844 13636 4846
rect 13468 4732 13524 4788
rect 12908 4450 12964 4452
rect 12908 4398 12910 4450
rect 12910 4398 12962 4450
rect 12962 4398 12964 4450
rect 12908 4396 12964 4398
rect 13468 4396 13524 4452
rect 14028 4450 14084 4452
rect 14028 4398 14030 4450
rect 14030 4398 14082 4450
rect 14082 4398 14084 4450
rect 14028 4396 14084 4398
rect 13804 4172 13860 4228
rect 13468 3948 13524 4004
rect 12012 3612 12068 3668
rect 12236 3500 12292 3556
rect 12572 3724 12628 3780
rect 11676 2716 11732 2772
rect 11116 2492 11172 2548
rect 11116 2268 11172 2324
rect 15036 5180 15092 5236
rect 15518 6298 15574 6300
rect 15518 6246 15520 6298
rect 15520 6246 15572 6298
rect 15572 6246 15574 6298
rect 15518 6244 15574 6246
rect 15622 6298 15678 6300
rect 15622 6246 15624 6298
rect 15624 6246 15676 6298
rect 15676 6246 15678 6298
rect 15622 6244 15678 6246
rect 15726 6298 15782 6300
rect 15726 6246 15728 6298
rect 15728 6246 15780 6298
rect 15780 6246 15782 6298
rect 15726 6244 15782 6246
rect 15820 6076 15876 6132
rect 15596 5180 15652 5236
rect 16268 8930 16324 8932
rect 16268 8878 16270 8930
rect 16270 8878 16322 8930
rect 16322 8878 16324 8930
rect 16268 8876 16324 8878
rect 16492 7644 16548 7700
rect 16380 6636 16436 6692
rect 16156 5740 16212 5796
rect 15932 5628 15988 5684
rect 15820 5068 15876 5124
rect 15148 4844 15204 4900
rect 14700 3554 14756 3556
rect 14700 3502 14702 3554
rect 14702 3502 14754 3554
rect 14754 3502 14756 3554
rect 14700 3500 14756 3502
rect 15036 4450 15092 4452
rect 15036 4398 15038 4450
rect 15038 4398 15090 4450
rect 15090 4398 15092 4450
rect 15036 4396 15092 4398
rect 15518 4730 15574 4732
rect 15518 4678 15520 4730
rect 15520 4678 15572 4730
rect 15572 4678 15574 4730
rect 15518 4676 15574 4678
rect 15622 4730 15678 4732
rect 15622 4678 15624 4730
rect 15624 4678 15676 4730
rect 15676 4678 15678 4730
rect 15622 4676 15678 4678
rect 15726 4730 15782 4732
rect 15726 4678 15728 4730
rect 15728 4678 15780 4730
rect 15780 4678 15782 4730
rect 15726 4676 15782 4678
rect 15932 4620 15988 4676
rect 16044 4396 16100 4452
rect 15820 3948 15876 4004
rect 16268 4226 16324 4228
rect 16268 4174 16270 4226
rect 16270 4174 16322 4226
rect 16322 4174 16324 4226
rect 16268 4172 16324 4174
rect 16380 3778 16436 3780
rect 16380 3726 16382 3778
rect 16382 3726 16434 3778
rect 16434 3726 16436 3778
rect 16380 3724 16436 3726
rect 14812 3388 14868 3444
rect 15518 3162 15574 3164
rect 15518 3110 15520 3162
rect 15520 3110 15572 3162
rect 15572 3110 15574 3162
rect 15518 3108 15574 3110
rect 15622 3162 15678 3164
rect 15622 3110 15624 3162
rect 15624 3110 15676 3162
rect 15676 3110 15678 3162
rect 15622 3108 15678 3110
rect 15726 3162 15782 3164
rect 15726 3110 15728 3162
rect 15728 3110 15780 3162
rect 15780 3110 15782 3162
rect 15726 3108 15782 3110
rect 16492 2828 16548 2884
rect 15260 2380 15316 2436
rect 17164 9436 17220 9492
rect 17388 10220 17444 10276
rect 16828 9154 16884 9156
rect 16828 9102 16830 9154
rect 16830 9102 16882 9154
rect 16882 9102 16884 9154
rect 16828 9100 16884 9102
rect 16828 8316 16884 8372
rect 17164 8258 17220 8260
rect 17164 8206 17166 8258
rect 17166 8206 17218 8258
rect 17218 8206 17220 8258
rect 17164 8204 17220 8206
rect 17836 12236 17892 12292
rect 18060 12236 18116 12292
rect 18172 13468 18228 13524
rect 19292 17724 19348 17780
rect 19628 17724 19684 17780
rect 18956 15874 19012 15876
rect 18956 15822 18958 15874
rect 18958 15822 19010 15874
rect 19010 15822 19012 15874
rect 18956 15820 19012 15822
rect 19516 15820 19572 15876
rect 19740 16492 19796 16548
rect 19628 15484 19684 15540
rect 18956 13692 19012 13748
rect 18620 13468 18676 13524
rect 18844 12066 18900 12068
rect 18844 12014 18846 12066
rect 18846 12014 18898 12066
rect 18898 12014 18900 12066
rect 18844 12012 18900 12014
rect 18172 11900 18228 11956
rect 17948 11452 18004 11508
rect 17836 11394 17892 11396
rect 17836 11342 17838 11394
rect 17838 11342 17890 11394
rect 17890 11342 17892 11394
rect 17836 11340 17892 11342
rect 18620 11788 18676 11844
rect 18956 11788 19012 11844
rect 19068 11676 19124 11732
rect 18284 11116 18340 11172
rect 17836 10220 17892 10276
rect 18172 10108 18228 10164
rect 18060 9100 18116 9156
rect 17836 8876 17892 8932
rect 17500 8428 17556 8484
rect 18172 8764 18228 8820
rect 17724 8316 17780 8372
rect 17500 8204 17556 8260
rect 17836 7756 17892 7812
rect 17500 6860 17556 6916
rect 16828 6748 16884 6804
rect 17836 6636 17892 6692
rect 17500 6578 17556 6580
rect 17500 6526 17502 6578
rect 17502 6526 17554 6578
rect 17554 6526 17556 6578
rect 17500 6524 17556 6526
rect 16716 6300 16772 6356
rect 17052 6076 17108 6132
rect 16716 5852 16772 5908
rect 17388 5122 17444 5124
rect 17388 5070 17390 5122
rect 17390 5070 17442 5122
rect 17442 5070 17444 5122
rect 17388 5068 17444 5070
rect 16828 4956 16884 5012
rect 17724 4732 17780 4788
rect 16716 4172 16772 4228
rect 17500 4338 17556 4340
rect 17500 4286 17502 4338
rect 17502 4286 17554 4338
rect 17554 4286 17556 4338
rect 17500 4284 17556 4286
rect 17500 3948 17556 4004
rect 16604 2156 16660 2212
rect 17500 3388 17556 3444
rect 18060 5292 18116 5348
rect 18732 11116 18788 11172
rect 20524 26796 20580 26852
rect 20748 26572 20804 26628
rect 20524 25340 20580 25396
rect 21084 23884 21140 23940
rect 20412 22316 20468 22372
rect 20188 21868 20244 21924
rect 20300 21084 20356 21140
rect 21308 25452 21364 25508
rect 21532 26124 21588 26180
rect 21868 26572 21924 26628
rect 21532 25788 21588 25844
rect 21644 25394 21700 25396
rect 21644 25342 21646 25394
rect 21646 25342 21698 25394
rect 21698 25342 21700 25394
rect 21644 25340 21700 25342
rect 21420 24050 21476 24052
rect 21420 23998 21422 24050
rect 21422 23998 21474 24050
rect 21474 23998 21476 24050
rect 21420 23996 21476 23998
rect 21420 23772 21476 23828
rect 21196 22540 21252 22596
rect 21308 23660 21364 23716
rect 21084 22204 21140 22260
rect 20972 20860 21028 20916
rect 20188 19906 20244 19908
rect 20188 19854 20190 19906
rect 20190 19854 20242 19906
rect 20242 19854 20244 19906
rect 20188 19852 20244 19854
rect 20188 19516 20244 19572
rect 20076 19234 20132 19236
rect 20076 19182 20078 19234
rect 20078 19182 20130 19234
rect 20130 19182 20132 19234
rect 20076 19180 20132 19182
rect 20188 17778 20244 17780
rect 20188 17726 20190 17778
rect 20190 17726 20242 17778
rect 20242 17726 20244 17778
rect 20188 17724 20244 17726
rect 22316 27468 22372 27524
rect 22204 27132 22260 27188
rect 22672 30602 22728 30604
rect 22672 30550 22674 30602
rect 22674 30550 22726 30602
rect 22726 30550 22728 30602
rect 22672 30548 22728 30550
rect 22776 30602 22832 30604
rect 22776 30550 22778 30602
rect 22778 30550 22830 30602
rect 22830 30550 22832 30602
rect 22776 30548 22832 30550
rect 22880 30602 22936 30604
rect 22880 30550 22882 30602
rect 22882 30550 22934 30602
rect 22934 30550 22936 30602
rect 22880 30548 22936 30550
rect 23996 30940 24052 30996
rect 23324 30716 23380 30772
rect 23548 30604 23604 30660
rect 24444 30716 24500 30772
rect 24556 30604 24612 30660
rect 23548 30156 23604 30212
rect 23996 29986 24052 29988
rect 23996 29934 23998 29986
rect 23998 29934 24050 29986
rect 24050 29934 24052 29986
rect 23996 29932 24052 29934
rect 24332 29596 24388 29652
rect 23548 29372 23604 29428
rect 23772 29426 23828 29428
rect 23772 29374 23774 29426
rect 23774 29374 23826 29426
rect 23826 29374 23828 29426
rect 23772 29372 23828 29374
rect 24780 29932 24836 29988
rect 24220 29260 24276 29316
rect 22672 29034 22728 29036
rect 22672 28982 22674 29034
rect 22674 28982 22726 29034
rect 22726 28982 22728 29034
rect 22672 28980 22728 28982
rect 22776 29034 22832 29036
rect 22776 28982 22778 29034
rect 22778 28982 22830 29034
rect 22830 28982 22832 29034
rect 22776 28980 22832 28982
rect 22880 29034 22936 29036
rect 22880 28982 22882 29034
rect 22882 28982 22934 29034
rect 22934 28982 22936 29034
rect 22880 28980 22936 28982
rect 23324 29036 23380 29092
rect 22988 28700 23044 28756
rect 22540 28588 22596 28644
rect 23436 28924 23492 28980
rect 23324 28642 23380 28644
rect 23324 28590 23326 28642
rect 23326 28590 23378 28642
rect 23378 28590 23380 28642
rect 23324 28588 23380 28590
rect 23996 28642 24052 28644
rect 23996 28590 23998 28642
rect 23998 28590 24050 28642
rect 24050 28590 24052 28642
rect 23996 28588 24052 28590
rect 24892 28754 24948 28756
rect 24892 28702 24894 28754
rect 24894 28702 24946 28754
rect 24946 28702 24948 28754
rect 24892 28700 24948 28702
rect 23324 28140 23380 28196
rect 22876 27746 22932 27748
rect 22876 27694 22878 27746
rect 22878 27694 22930 27746
rect 22930 27694 22932 27746
rect 22876 27692 22932 27694
rect 22672 27466 22728 27468
rect 22672 27414 22674 27466
rect 22674 27414 22726 27466
rect 22726 27414 22728 27466
rect 22672 27412 22728 27414
rect 22776 27466 22832 27468
rect 22776 27414 22778 27466
rect 22778 27414 22830 27466
rect 22830 27414 22832 27466
rect 22776 27412 22832 27414
rect 22880 27466 22936 27468
rect 22880 27414 22882 27466
rect 22882 27414 22934 27466
rect 22934 27414 22936 27466
rect 22880 27412 22936 27414
rect 22876 27244 22932 27300
rect 22540 27074 22596 27076
rect 22540 27022 22542 27074
rect 22542 27022 22594 27074
rect 22594 27022 22596 27074
rect 22540 27020 22596 27022
rect 22652 26962 22708 26964
rect 22652 26910 22654 26962
rect 22654 26910 22706 26962
rect 22706 26910 22708 26962
rect 22652 26908 22708 26910
rect 22316 26850 22372 26852
rect 22316 26798 22318 26850
rect 22318 26798 22370 26850
rect 22370 26798 22372 26850
rect 22316 26796 22372 26798
rect 22316 26572 22372 26628
rect 22428 25788 22484 25844
rect 22428 25340 22484 25396
rect 22316 25004 22372 25060
rect 21980 24892 22036 24948
rect 21532 22370 21588 22372
rect 21532 22318 21534 22370
rect 21534 22318 21586 22370
rect 21586 22318 21588 22370
rect 21532 22316 21588 22318
rect 21644 21980 21700 22036
rect 21644 21756 21700 21812
rect 21308 20636 21364 20692
rect 21420 20748 21476 20804
rect 20636 19852 20692 19908
rect 20972 19180 21028 19236
rect 20636 18396 20692 18452
rect 20524 17666 20580 17668
rect 20524 17614 20526 17666
rect 20526 17614 20578 17666
rect 20578 17614 20580 17666
rect 20524 17612 20580 17614
rect 20076 15874 20132 15876
rect 20076 15822 20078 15874
rect 20078 15822 20130 15874
rect 20130 15822 20132 15874
rect 20076 15820 20132 15822
rect 20412 17500 20468 17556
rect 20300 16770 20356 16772
rect 20300 16718 20302 16770
rect 20302 16718 20354 16770
rect 20354 16718 20356 16770
rect 20300 16716 20356 16718
rect 20188 14924 20244 14980
rect 20188 14140 20244 14196
rect 20300 16492 20356 16548
rect 19740 12572 19796 12628
rect 19740 12348 19796 12404
rect 19852 12290 19908 12292
rect 19852 12238 19854 12290
rect 19854 12238 19906 12290
rect 19906 12238 19908 12290
rect 19852 12236 19908 12238
rect 19964 11900 20020 11956
rect 20076 11788 20132 11844
rect 20860 17106 20916 17108
rect 20860 17054 20862 17106
rect 20862 17054 20914 17106
rect 20914 17054 20916 17106
rect 20860 17052 20916 17054
rect 20188 12124 20244 12180
rect 20300 11900 20356 11956
rect 20300 11676 20356 11732
rect 20188 11564 20244 11620
rect 19740 11452 19796 11508
rect 19964 11394 20020 11396
rect 19964 11342 19966 11394
rect 19966 11342 20018 11394
rect 20018 11342 20020 11394
rect 19964 11340 20020 11342
rect 19292 11116 19348 11172
rect 19740 10668 19796 10724
rect 19292 10610 19348 10612
rect 19292 10558 19294 10610
rect 19294 10558 19346 10610
rect 19346 10558 19348 10610
rect 19292 10556 19348 10558
rect 19180 10498 19236 10500
rect 19180 10446 19182 10498
rect 19182 10446 19234 10498
rect 19234 10446 19236 10498
rect 19180 10444 19236 10446
rect 18620 8652 18676 8708
rect 18396 8316 18452 8372
rect 18284 5794 18340 5796
rect 18284 5742 18286 5794
rect 18286 5742 18338 5794
rect 18338 5742 18340 5794
rect 18284 5740 18340 5742
rect 18284 4508 18340 4564
rect 18060 4338 18116 4340
rect 18060 4286 18062 4338
rect 18062 4286 18114 4338
rect 18114 4286 18116 4338
rect 18060 4284 18116 4286
rect 17836 3276 17892 3332
rect 18508 5180 18564 5236
rect 19628 10332 19684 10388
rect 19068 9324 19124 9380
rect 19740 9548 19796 9604
rect 20972 16994 21028 16996
rect 20972 16942 20974 16994
rect 20974 16942 21026 16994
rect 21026 16942 21028 16994
rect 20972 16940 21028 16942
rect 21532 19516 21588 19572
rect 22092 22316 22148 22372
rect 22428 22370 22484 22372
rect 22428 22318 22430 22370
rect 22430 22318 22482 22370
rect 22482 22318 22484 22370
rect 22428 22316 22484 22318
rect 22092 21980 22148 22036
rect 21980 20802 22036 20804
rect 21980 20750 21982 20802
rect 21982 20750 22034 20802
rect 22034 20750 22036 20802
rect 21980 20748 22036 20750
rect 22428 21644 22484 21700
rect 22092 20076 22148 20132
rect 22204 18450 22260 18452
rect 22204 18398 22206 18450
rect 22206 18398 22258 18450
rect 22258 18398 22260 18450
rect 22204 18396 22260 18398
rect 21308 18284 21364 18340
rect 21980 18338 22036 18340
rect 21980 18286 21982 18338
rect 21982 18286 22034 18338
rect 22034 18286 22036 18338
rect 21980 18284 22036 18286
rect 22316 17836 22372 17892
rect 21308 17612 21364 17668
rect 21532 17554 21588 17556
rect 21532 17502 21534 17554
rect 21534 17502 21586 17554
rect 21586 17502 21588 17554
rect 21532 17500 21588 17502
rect 22988 27132 23044 27188
rect 24556 28418 24612 28420
rect 24556 28366 24558 28418
rect 24558 28366 24610 28418
rect 24610 28366 24612 28418
rect 24556 28364 24612 28366
rect 23324 27356 23380 27412
rect 23884 27132 23940 27188
rect 23212 26572 23268 26628
rect 23548 26908 23604 26964
rect 22876 26290 22932 26292
rect 22876 26238 22878 26290
rect 22878 26238 22930 26290
rect 22930 26238 22932 26290
rect 22876 26236 22932 26238
rect 23772 26290 23828 26292
rect 23772 26238 23774 26290
rect 23774 26238 23826 26290
rect 23826 26238 23828 26290
rect 23772 26236 23828 26238
rect 22672 25898 22728 25900
rect 22672 25846 22674 25898
rect 22674 25846 22726 25898
rect 22726 25846 22728 25898
rect 22672 25844 22728 25846
rect 22776 25898 22832 25900
rect 22776 25846 22778 25898
rect 22778 25846 22830 25898
rect 22830 25846 22832 25898
rect 22776 25844 22832 25846
rect 22880 25898 22936 25900
rect 22880 25846 22882 25898
rect 22882 25846 22934 25898
rect 22934 25846 22936 25898
rect 22880 25844 22936 25846
rect 22876 25116 22932 25172
rect 24668 27746 24724 27748
rect 24668 27694 24670 27746
rect 24670 27694 24722 27746
rect 24722 27694 24724 27746
rect 24668 27692 24724 27694
rect 25228 34972 25284 35028
rect 25900 35420 25956 35476
rect 26348 34972 26404 35028
rect 26460 34914 26516 34916
rect 26460 34862 26462 34914
rect 26462 34862 26514 34914
rect 26514 34862 26516 34914
rect 26460 34860 26516 34862
rect 26124 34690 26180 34692
rect 26124 34638 26126 34690
rect 26126 34638 26178 34690
rect 26178 34638 26180 34690
rect 26124 34636 26180 34638
rect 25228 34076 25284 34132
rect 25340 33906 25396 33908
rect 25340 33854 25342 33906
rect 25342 33854 25394 33906
rect 25394 33854 25396 33906
rect 25340 33852 25396 33854
rect 26012 34076 26068 34132
rect 25676 33852 25732 33908
rect 27580 34300 27636 34356
rect 26908 33852 26964 33908
rect 27580 33852 27636 33908
rect 27356 33628 27412 33684
rect 27244 33346 27300 33348
rect 27244 33294 27246 33346
rect 27246 33294 27298 33346
rect 27298 33294 27300 33346
rect 27244 33292 27300 33294
rect 28812 37100 28868 37156
rect 28364 36316 28420 36372
rect 27804 35532 27860 35588
rect 28476 36204 28532 36260
rect 28476 35308 28532 35364
rect 29148 36370 29204 36372
rect 29148 36318 29150 36370
rect 29150 36318 29202 36370
rect 29202 36318 29204 36370
rect 29148 36316 29204 36318
rect 33292 36988 33348 37044
rect 32060 36876 32116 36932
rect 29825 36090 29881 36092
rect 29825 36038 29827 36090
rect 29827 36038 29879 36090
rect 29879 36038 29881 36090
rect 29825 36036 29881 36038
rect 29929 36090 29985 36092
rect 29929 36038 29931 36090
rect 29931 36038 29983 36090
rect 29983 36038 29985 36090
rect 29929 36036 29985 36038
rect 30033 36090 30089 36092
rect 30033 36038 30035 36090
rect 30035 36038 30087 36090
rect 30087 36038 30089 36090
rect 30033 36036 30089 36038
rect 28924 35586 28980 35588
rect 28924 35534 28926 35586
rect 28926 35534 28978 35586
rect 28978 35534 28980 35586
rect 28924 35532 28980 35534
rect 29596 35308 29652 35364
rect 30156 35308 30212 35364
rect 32620 36482 32676 36484
rect 32620 36430 32622 36482
rect 32622 36430 32674 36482
rect 32674 36430 32676 36482
rect 32620 36428 32676 36430
rect 31836 36092 31892 36148
rect 31724 34860 31780 34916
rect 29372 34524 29428 34580
rect 29825 34522 29881 34524
rect 29825 34470 29827 34522
rect 29827 34470 29879 34522
rect 29879 34470 29881 34522
rect 29825 34468 29881 34470
rect 29929 34522 29985 34524
rect 29929 34470 29931 34522
rect 29931 34470 29983 34522
rect 29983 34470 29985 34522
rect 29929 34468 29985 34470
rect 30033 34522 30089 34524
rect 30033 34470 30035 34522
rect 30035 34470 30087 34522
rect 30087 34470 30089 34522
rect 30033 34468 30089 34470
rect 31612 34524 31668 34580
rect 27580 33404 27636 33460
rect 28476 33852 28532 33908
rect 26572 33122 26628 33124
rect 26572 33070 26574 33122
rect 26574 33070 26626 33122
rect 26626 33070 26628 33122
rect 26572 33068 26628 33070
rect 27692 33346 27748 33348
rect 27692 33294 27694 33346
rect 27694 33294 27746 33346
rect 27746 33294 27748 33346
rect 27692 33292 27748 33294
rect 25676 32284 25732 32340
rect 25676 31948 25732 32004
rect 26124 31724 26180 31780
rect 25676 31554 25732 31556
rect 25676 31502 25678 31554
rect 25678 31502 25730 31554
rect 25730 31502 25732 31554
rect 25676 31500 25732 31502
rect 27132 32508 27188 32564
rect 26348 31724 26404 31780
rect 26460 31948 26516 32004
rect 26012 30210 26068 30212
rect 26012 30158 26014 30210
rect 26014 30158 26066 30210
rect 26066 30158 26068 30210
rect 26012 30156 26068 30158
rect 25676 29650 25732 29652
rect 25676 29598 25678 29650
rect 25678 29598 25730 29650
rect 25730 29598 25732 29650
rect 25676 29596 25732 29598
rect 25116 29036 25172 29092
rect 25788 28700 25844 28756
rect 25900 28924 25956 28980
rect 25452 28588 25508 28644
rect 25788 28418 25844 28420
rect 25788 28366 25790 28418
rect 25790 28366 25842 28418
rect 25842 28366 25844 28418
rect 25788 28364 25844 28366
rect 25228 27746 25284 27748
rect 25228 27694 25230 27746
rect 25230 27694 25282 27746
rect 25282 27694 25284 27746
rect 25228 27692 25284 27694
rect 26012 27692 26068 27748
rect 25900 27634 25956 27636
rect 25900 27582 25902 27634
rect 25902 27582 25954 27634
rect 25954 27582 25956 27634
rect 25900 27580 25956 27582
rect 25452 27468 25508 27524
rect 24892 27132 24948 27188
rect 26236 27634 26292 27636
rect 26236 27582 26238 27634
rect 26238 27582 26290 27634
rect 26290 27582 26292 27634
rect 26236 27580 26292 27582
rect 24332 26962 24388 26964
rect 24332 26910 24334 26962
rect 24334 26910 24386 26962
rect 24386 26910 24388 26962
rect 24332 26908 24388 26910
rect 26236 26962 26292 26964
rect 26236 26910 26238 26962
rect 26238 26910 26290 26962
rect 26290 26910 26292 26962
rect 26236 26908 26292 26910
rect 28588 33458 28644 33460
rect 28588 33406 28590 33458
rect 28590 33406 28642 33458
rect 28642 33406 28644 33458
rect 28588 33404 28644 33406
rect 29372 34354 29428 34356
rect 29372 34302 29374 34354
rect 29374 34302 29426 34354
rect 29426 34302 29428 34354
rect 29372 34300 29428 34302
rect 29932 34300 29988 34356
rect 30940 34354 30996 34356
rect 30940 34302 30942 34354
rect 30942 34302 30994 34354
rect 30994 34302 30996 34354
rect 30940 34300 30996 34302
rect 31500 34130 31556 34132
rect 31500 34078 31502 34130
rect 31502 34078 31554 34130
rect 31554 34078 31556 34130
rect 31500 34076 31556 34078
rect 29596 33458 29652 33460
rect 29596 33406 29598 33458
rect 29598 33406 29650 33458
rect 29650 33406 29652 33458
rect 29596 33404 29652 33406
rect 28812 33292 28868 33348
rect 29148 33292 29204 33348
rect 27692 32396 27748 32452
rect 28028 32732 28084 32788
rect 28252 32450 28308 32452
rect 28252 32398 28254 32450
rect 28254 32398 28306 32450
rect 28306 32398 28308 32450
rect 28252 32396 28308 32398
rect 27916 31836 27972 31892
rect 27356 31778 27412 31780
rect 27356 31726 27358 31778
rect 27358 31726 27410 31778
rect 27410 31726 27412 31778
rect 27356 31724 27412 31726
rect 26572 31500 26628 31556
rect 26684 31164 26740 31220
rect 26908 31052 26964 31108
rect 26908 28476 26964 28532
rect 27580 31554 27636 31556
rect 27580 31502 27582 31554
rect 27582 31502 27634 31554
rect 27634 31502 27636 31554
rect 27580 31500 27636 31502
rect 29484 33346 29540 33348
rect 29484 33294 29486 33346
rect 29486 33294 29538 33346
rect 29538 33294 29540 33346
rect 29484 33292 29540 33294
rect 29372 33068 29428 33124
rect 29148 32338 29204 32340
rect 29148 32286 29150 32338
rect 29150 32286 29202 32338
rect 29202 32286 29204 32338
rect 29148 32284 29204 32286
rect 29825 32954 29881 32956
rect 29825 32902 29827 32954
rect 29827 32902 29879 32954
rect 29879 32902 29881 32954
rect 29825 32900 29881 32902
rect 29929 32954 29985 32956
rect 29929 32902 29931 32954
rect 29931 32902 29983 32954
rect 29983 32902 29985 32954
rect 29929 32900 29985 32902
rect 30033 32954 30089 32956
rect 30033 32902 30035 32954
rect 30035 32902 30087 32954
rect 30087 32902 30089 32954
rect 30033 32900 30089 32902
rect 29596 32284 29652 32340
rect 30492 33068 30548 33124
rect 30940 33122 30996 33124
rect 30940 33070 30942 33122
rect 30942 33070 30994 33122
rect 30994 33070 30996 33122
rect 30940 33068 30996 33070
rect 30604 32956 30660 33012
rect 30380 32674 30436 32676
rect 30380 32622 30382 32674
rect 30382 32622 30434 32674
rect 30434 32622 30436 32674
rect 30380 32620 30436 32622
rect 30268 32562 30324 32564
rect 30268 32510 30270 32562
rect 30270 32510 30322 32562
rect 30322 32510 30324 32562
rect 30268 32508 30324 32510
rect 30828 32562 30884 32564
rect 30828 32510 30830 32562
rect 30830 32510 30882 32562
rect 30882 32510 30884 32562
rect 30828 32508 30884 32510
rect 31388 32450 31444 32452
rect 31388 32398 31390 32450
rect 31390 32398 31442 32450
rect 31442 32398 31444 32450
rect 31388 32396 31444 32398
rect 30156 31948 30212 32004
rect 27692 31052 27748 31108
rect 28364 30882 28420 30884
rect 28364 30830 28366 30882
rect 28366 30830 28418 30882
rect 28418 30830 28420 30882
rect 28364 30828 28420 30830
rect 28252 30492 28308 30548
rect 28476 30380 28532 30436
rect 27580 29372 27636 29428
rect 27132 28530 27188 28532
rect 27132 28478 27134 28530
rect 27134 28478 27186 28530
rect 27186 28478 27188 28530
rect 27132 28476 27188 28478
rect 27020 27916 27076 27972
rect 24220 26236 24276 26292
rect 24892 26572 24948 26628
rect 24668 26290 24724 26292
rect 24668 26238 24670 26290
rect 24670 26238 24722 26290
rect 24722 26238 24724 26290
rect 24668 26236 24724 26238
rect 24556 25900 24612 25956
rect 24556 25564 24612 25620
rect 24332 24892 24388 24948
rect 22672 24330 22728 24332
rect 22672 24278 22674 24330
rect 22674 24278 22726 24330
rect 22726 24278 22728 24330
rect 22672 24276 22728 24278
rect 22776 24330 22832 24332
rect 22776 24278 22778 24330
rect 22778 24278 22830 24330
rect 22830 24278 22832 24330
rect 22776 24276 22832 24278
rect 22880 24330 22936 24332
rect 22880 24278 22882 24330
rect 22882 24278 22934 24330
rect 22934 24278 22936 24330
rect 22880 24276 22936 24278
rect 23772 24722 23828 24724
rect 23772 24670 23774 24722
rect 23774 24670 23826 24722
rect 23826 24670 23828 24722
rect 23772 24668 23828 24670
rect 23212 24220 23268 24276
rect 23212 23884 23268 23940
rect 24668 24556 24724 24612
rect 24556 23714 24612 23716
rect 24556 23662 24558 23714
rect 24558 23662 24610 23714
rect 24610 23662 24612 23714
rect 24556 23660 24612 23662
rect 24444 23548 24500 23604
rect 23100 23100 23156 23156
rect 22672 22762 22728 22764
rect 22672 22710 22674 22762
rect 22674 22710 22726 22762
rect 22726 22710 22728 22762
rect 22672 22708 22728 22710
rect 22776 22762 22832 22764
rect 22776 22710 22778 22762
rect 22778 22710 22830 22762
rect 22830 22710 22832 22762
rect 22776 22708 22832 22710
rect 22880 22762 22936 22764
rect 22880 22710 22882 22762
rect 22882 22710 22934 22762
rect 22934 22710 22936 22762
rect 22880 22708 22936 22710
rect 23100 22540 23156 22596
rect 22876 22370 22932 22372
rect 22876 22318 22878 22370
rect 22878 22318 22930 22370
rect 22930 22318 22932 22370
rect 22876 22316 22932 22318
rect 24332 23100 24388 23156
rect 24220 22540 24276 22596
rect 23996 22258 24052 22260
rect 23996 22206 23998 22258
rect 23998 22206 24050 22258
rect 24050 22206 24052 22258
rect 23996 22204 24052 22206
rect 24220 22146 24276 22148
rect 24220 22094 24222 22146
rect 24222 22094 24274 22146
rect 24274 22094 24276 22146
rect 24220 22092 24276 22094
rect 24444 22146 24500 22148
rect 24444 22094 24446 22146
rect 24446 22094 24498 22146
rect 24498 22094 24500 22146
rect 24444 22092 24500 22094
rect 22764 21810 22820 21812
rect 22764 21758 22766 21810
rect 22766 21758 22818 21810
rect 22818 21758 22820 21810
rect 22764 21756 22820 21758
rect 22672 21194 22728 21196
rect 22672 21142 22674 21194
rect 22674 21142 22726 21194
rect 22726 21142 22728 21194
rect 22672 21140 22728 21142
rect 22776 21194 22832 21196
rect 22776 21142 22778 21194
rect 22778 21142 22830 21194
rect 22830 21142 22832 21194
rect 22776 21140 22832 21142
rect 22880 21194 22936 21196
rect 22880 21142 22882 21194
rect 22882 21142 22934 21194
rect 22934 21142 22936 21194
rect 22880 21140 22936 21142
rect 23100 20076 23156 20132
rect 22672 19626 22728 19628
rect 22672 19574 22674 19626
rect 22674 19574 22726 19626
rect 22726 19574 22728 19626
rect 22672 19572 22728 19574
rect 22776 19626 22832 19628
rect 22776 19574 22778 19626
rect 22778 19574 22830 19626
rect 22830 19574 22832 19626
rect 22776 19572 22832 19574
rect 22880 19626 22936 19628
rect 22880 19574 22882 19626
rect 22882 19574 22934 19626
rect 22934 19574 22936 19626
rect 22880 19572 22936 19574
rect 22764 19180 22820 19236
rect 22876 19292 22932 19348
rect 23772 20636 23828 20692
rect 24332 19852 24388 19908
rect 23996 19346 24052 19348
rect 23996 19294 23998 19346
rect 23998 19294 24050 19346
rect 24050 19294 24052 19346
rect 23996 19292 24052 19294
rect 24668 20130 24724 20132
rect 24668 20078 24670 20130
rect 24670 20078 24722 20130
rect 24722 20078 24724 20130
rect 24668 20076 24724 20078
rect 25228 26572 25284 26628
rect 25564 26290 25620 26292
rect 25564 26238 25566 26290
rect 25566 26238 25618 26290
rect 25618 26238 25620 26290
rect 25564 26236 25620 26238
rect 25228 25452 25284 25508
rect 25788 25340 25844 25396
rect 25340 24556 25396 24612
rect 25004 24444 25060 24500
rect 25228 23714 25284 23716
rect 25228 23662 25230 23714
rect 25230 23662 25282 23714
rect 25282 23662 25284 23714
rect 25228 23660 25284 23662
rect 26124 24556 26180 24612
rect 25340 22988 25396 23044
rect 25228 22652 25284 22708
rect 25228 22316 25284 22372
rect 24892 22258 24948 22260
rect 24892 22206 24894 22258
rect 24894 22206 24946 22258
rect 24946 22206 24948 22258
rect 24892 22204 24948 22206
rect 25116 21868 25172 21924
rect 25340 22146 25396 22148
rect 25340 22094 25342 22146
rect 25342 22094 25394 22146
rect 25394 22094 25396 22146
rect 25340 22092 25396 22094
rect 25228 21420 25284 21476
rect 25228 20860 25284 20916
rect 26012 22204 26068 22260
rect 25788 21980 25844 22036
rect 26124 21980 26180 22036
rect 25900 21868 25956 21924
rect 26236 21420 26292 21476
rect 26348 21196 26404 21252
rect 26012 20188 26068 20244
rect 27356 27804 27412 27860
rect 27356 27468 27412 27524
rect 27580 28924 27636 28980
rect 28588 30210 28644 30212
rect 28588 30158 28590 30210
rect 28590 30158 28642 30210
rect 28642 30158 28644 30210
rect 28588 30156 28644 30158
rect 28252 29708 28308 29764
rect 27916 29260 27972 29316
rect 29148 31666 29204 31668
rect 29148 31614 29150 31666
rect 29150 31614 29202 31666
rect 29202 31614 29204 31666
rect 29148 31612 29204 31614
rect 29825 31386 29881 31388
rect 29825 31334 29827 31386
rect 29827 31334 29879 31386
rect 29879 31334 29881 31386
rect 29825 31332 29881 31334
rect 29929 31386 29985 31388
rect 29929 31334 29931 31386
rect 29931 31334 29983 31386
rect 29983 31334 29985 31386
rect 29929 31332 29985 31334
rect 30033 31386 30089 31388
rect 30033 31334 30035 31386
rect 30035 31334 30087 31386
rect 30087 31334 30089 31386
rect 30033 31332 30089 31334
rect 29372 31164 29428 31220
rect 28924 30716 28980 30772
rect 29372 30882 29428 30884
rect 29372 30830 29374 30882
rect 29374 30830 29426 30882
rect 29426 30830 29428 30882
rect 29372 30828 29428 30830
rect 29820 30828 29876 30884
rect 29372 30492 29428 30548
rect 29484 30380 29540 30436
rect 30604 30882 30660 30884
rect 30604 30830 30606 30882
rect 30606 30830 30658 30882
rect 30658 30830 30660 30882
rect 30604 30828 30660 30830
rect 30156 30380 30212 30436
rect 32172 35308 32228 35364
rect 31836 34748 31892 34804
rect 32172 34130 32228 34132
rect 32172 34078 32174 34130
rect 32174 34078 32226 34130
rect 32226 34078 32228 34130
rect 32172 34076 32228 34078
rect 32396 34018 32452 34020
rect 32396 33966 32398 34018
rect 32398 33966 32450 34018
rect 32450 33966 32452 34018
rect 32396 33964 32452 33966
rect 32732 33964 32788 34020
rect 32956 34636 33012 34692
rect 32956 34076 33012 34132
rect 32844 33852 32900 33908
rect 33740 36876 33796 36932
rect 33964 35420 34020 35476
rect 33740 34972 33796 35028
rect 34524 36988 34580 37044
rect 35308 36540 35364 36596
rect 35532 35756 35588 35812
rect 34524 35420 34580 35476
rect 34300 35196 34356 35252
rect 35084 35196 35140 35252
rect 35308 35084 35364 35140
rect 33852 34690 33908 34692
rect 33852 34638 33854 34690
rect 33854 34638 33906 34690
rect 33906 34638 33908 34690
rect 33852 34636 33908 34638
rect 34188 34690 34244 34692
rect 34188 34638 34190 34690
rect 34190 34638 34242 34690
rect 34242 34638 34244 34690
rect 34188 34636 34244 34638
rect 33516 34300 33572 34356
rect 34860 34300 34916 34356
rect 33964 34018 34020 34020
rect 33964 33966 33966 34018
rect 33966 33966 34018 34018
rect 34018 33966 34020 34018
rect 33964 33964 34020 33966
rect 33292 33404 33348 33460
rect 31836 32956 31892 33012
rect 32620 32956 32676 33012
rect 33180 32562 33236 32564
rect 33180 32510 33182 32562
rect 33182 32510 33234 32562
rect 33234 32510 33236 32562
rect 33180 32508 33236 32510
rect 36979 36874 37035 36876
rect 36979 36822 36981 36874
rect 36981 36822 37033 36874
rect 37033 36822 37035 36874
rect 36979 36820 37035 36822
rect 37083 36874 37139 36876
rect 37083 36822 37085 36874
rect 37085 36822 37137 36874
rect 37137 36822 37139 36874
rect 37083 36820 37139 36822
rect 37187 36874 37243 36876
rect 37187 36822 37189 36874
rect 37189 36822 37241 36874
rect 37241 36822 37243 36874
rect 37187 36820 37243 36822
rect 37212 36540 37268 36596
rect 35868 35756 35924 35812
rect 36428 35756 36484 35812
rect 37772 35644 37828 35700
rect 37436 35586 37492 35588
rect 37436 35534 37438 35586
rect 37438 35534 37490 35586
rect 37490 35534 37492 35586
rect 37436 35532 37492 35534
rect 36428 35420 36484 35476
rect 38556 36316 38612 36372
rect 37996 35420 38052 35476
rect 36979 35306 37035 35308
rect 36979 35254 36981 35306
rect 36981 35254 37033 35306
rect 37033 35254 37035 35306
rect 36979 35252 37035 35254
rect 37083 35306 37139 35308
rect 37083 35254 37085 35306
rect 37085 35254 37137 35306
rect 37137 35254 37139 35306
rect 37083 35252 37139 35254
rect 37187 35306 37243 35308
rect 37187 35254 37189 35306
rect 37189 35254 37241 35306
rect 37241 35254 37243 35306
rect 37187 35252 37243 35254
rect 37660 35308 37716 35364
rect 36988 35026 37044 35028
rect 36988 34974 36990 35026
rect 36990 34974 37042 35026
rect 37042 34974 37044 35026
rect 36988 34972 37044 34974
rect 37212 34972 37268 35028
rect 35980 34300 36036 34356
rect 34636 33404 34692 33460
rect 34524 33234 34580 33236
rect 34524 33182 34526 33234
rect 34526 33182 34578 33234
rect 34578 33182 34580 33234
rect 34524 33180 34580 33182
rect 34860 33404 34916 33460
rect 34972 33346 35028 33348
rect 34972 33294 34974 33346
rect 34974 33294 35026 33346
rect 35026 33294 35028 33346
rect 34972 33292 35028 33294
rect 33292 32396 33348 32452
rect 33516 32508 33572 32564
rect 34300 32562 34356 32564
rect 34300 32510 34302 32562
rect 34302 32510 34354 32562
rect 34354 32510 34356 32562
rect 34300 32508 34356 32510
rect 31724 31724 31780 31780
rect 31724 31500 31780 31556
rect 31500 30828 31556 30884
rect 29596 29708 29652 29764
rect 29708 29932 29764 29988
rect 29036 29426 29092 29428
rect 29036 29374 29038 29426
rect 29038 29374 29090 29426
rect 29090 29374 29092 29426
rect 29036 29372 29092 29374
rect 28812 29260 28868 29316
rect 29596 29260 29652 29316
rect 28476 28476 28532 28532
rect 28812 28028 28868 28084
rect 27692 27858 27748 27860
rect 27692 27806 27694 27858
rect 27694 27806 27746 27858
rect 27746 27806 27748 27858
rect 27692 27804 27748 27806
rect 28028 27692 28084 27748
rect 28588 27746 28644 27748
rect 28588 27694 28590 27746
rect 28590 27694 28642 27746
rect 28642 27694 28644 27746
rect 28588 27692 28644 27694
rect 28028 27468 28084 27524
rect 27916 26962 27972 26964
rect 27916 26910 27918 26962
rect 27918 26910 27970 26962
rect 27970 26910 27972 26962
rect 27916 26908 27972 26910
rect 27580 25340 27636 25396
rect 27132 25228 27188 25284
rect 28140 25676 28196 25732
rect 27916 25506 27972 25508
rect 27916 25454 27918 25506
rect 27918 25454 27970 25506
rect 27970 25454 27972 25506
rect 27916 25452 27972 25454
rect 27804 25394 27860 25396
rect 27804 25342 27806 25394
rect 27806 25342 27858 25394
rect 27858 25342 27860 25394
rect 27804 25340 27860 25342
rect 27692 24892 27748 24948
rect 27916 25228 27972 25284
rect 27020 24780 27076 24836
rect 27580 24780 27636 24836
rect 27020 24050 27076 24052
rect 27020 23998 27022 24050
rect 27022 23998 27074 24050
rect 27074 23998 27076 24050
rect 27020 23996 27076 23998
rect 28588 25676 28644 25732
rect 28812 25116 28868 25172
rect 28476 24892 28532 24948
rect 28028 24668 28084 24724
rect 27580 23996 27636 24052
rect 27020 23324 27076 23380
rect 26684 21868 26740 21924
rect 26796 22428 26852 22484
rect 26348 20076 26404 20132
rect 25676 19852 25732 19908
rect 23772 19234 23828 19236
rect 23772 19182 23774 19234
rect 23774 19182 23826 19234
rect 23826 19182 23828 19234
rect 23772 19180 23828 19182
rect 23772 18956 23828 19012
rect 23212 18508 23268 18564
rect 22672 18058 22728 18060
rect 22672 18006 22674 18058
rect 22674 18006 22726 18058
rect 22726 18006 22728 18058
rect 22672 18004 22728 18006
rect 22776 18058 22832 18060
rect 22776 18006 22778 18058
rect 22778 18006 22830 18058
rect 22830 18006 22832 18058
rect 22776 18004 22832 18006
rect 22880 18058 22936 18060
rect 22880 18006 22882 18058
rect 22882 18006 22934 18058
rect 22934 18006 22936 18058
rect 22880 18004 22936 18006
rect 21196 16828 21252 16884
rect 21756 16604 21812 16660
rect 21868 16828 21924 16884
rect 20860 16098 20916 16100
rect 20860 16046 20862 16098
rect 20862 16046 20914 16098
rect 20914 16046 20916 16098
rect 20860 16044 20916 16046
rect 21756 16044 21812 16100
rect 21084 15820 21140 15876
rect 20636 14252 20692 14308
rect 20524 13580 20580 13636
rect 20972 13634 21028 13636
rect 20972 13582 20974 13634
rect 20974 13582 21026 13634
rect 21026 13582 21028 13634
rect 20972 13580 21028 13582
rect 21644 15708 21700 15764
rect 21420 15372 21476 15428
rect 22092 16604 22148 16660
rect 22204 15986 22260 15988
rect 22204 15934 22206 15986
rect 22206 15934 22258 15986
rect 22258 15934 22260 15986
rect 22204 15932 22260 15934
rect 23100 17052 23156 17108
rect 21644 14924 21700 14980
rect 21308 14530 21364 14532
rect 21308 14478 21310 14530
rect 21310 14478 21362 14530
rect 21362 14478 21364 14530
rect 21308 14476 21364 14478
rect 21756 14588 21812 14644
rect 21084 13020 21140 13076
rect 21196 14364 21252 14420
rect 20636 12684 20692 12740
rect 20636 12348 20692 12404
rect 20524 11506 20580 11508
rect 20524 11454 20526 11506
rect 20526 11454 20578 11506
rect 20578 11454 20580 11506
rect 20524 11452 20580 11454
rect 20860 12012 20916 12068
rect 20748 11618 20804 11620
rect 20748 11566 20750 11618
rect 20750 11566 20802 11618
rect 20802 11566 20804 11618
rect 20748 11564 20804 11566
rect 20860 11452 20916 11508
rect 20524 10108 20580 10164
rect 20636 10780 20692 10836
rect 22204 13804 22260 13860
rect 21420 13580 21476 13636
rect 21868 13468 21924 13524
rect 21756 12908 21812 12964
rect 21308 11394 21364 11396
rect 21308 11342 21310 11394
rect 21310 11342 21362 11394
rect 21362 11342 21364 11394
rect 21308 11340 21364 11342
rect 20188 9602 20244 9604
rect 20188 9550 20190 9602
rect 20190 9550 20242 9602
rect 20242 9550 20244 9602
rect 20188 9548 20244 9550
rect 19628 9212 19684 9268
rect 20412 9100 20468 9156
rect 19740 8428 19796 8484
rect 19292 8092 19348 8148
rect 19180 7532 19236 7588
rect 18844 7474 18900 7476
rect 18844 7422 18846 7474
rect 18846 7422 18898 7474
rect 18898 7422 18900 7474
rect 18844 7420 18900 7422
rect 18732 7196 18788 7252
rect 18620 5068 18676 5124
rect 18508 4620 18564 4676
rect 19292 5068 19348 5124
rect 19180 4620 19236 4676
rect 19404 4396 19460 4452
rect 19068 4060 19124 4116
rect 20412 8428 20468 8484
rect 23548 17836 23604 17892
rect 23324 17052 23380 17108
rect 23324 16716 23380 16772
rect 23436 16940 23492 16996
rect 22672 16490 22728 16492
rect 22672 16438 22674 16490
rect 22674 16438 22726 16490
rect 22726 16438 22728 16490
rect 22672 16436 22728 16438
rect 22776 16490 22832 16492
rect 22776 16438 22778 16490
rect 22778 16438 22830 16490
rect 22830 16438 22832 16490
rect 22776 16436 22832 16438
rect 22880 16490 22936 16492
rect 22880 16438 22882 16490
rect 22882 16438 22934 16490
rect 22934 16438 22936 16490
rect 22880 16436 22936 16438
rect 23324 16098 23380 16100
rect 23324 16046 23326 16098
rect 23326 16046 23378 16098
rect 23378 16046 23380 16098
rect 23324 16044 23380 16046
rect 22540 15372 22596 15428
rect 22764 15148 22820 15204
rect 22672 14922 22728 14924
rect 22672 14870 22674 14922
rect 22674 14870 22726 14922
rect 22726 14870 22728 14922
rect 22672 14868 22728 14870
rect 22776 14922 22832 14924
rect 22776 14870 22778 14922
rect 22778 14870 22830 14922
rect 22830 14870 22832 14922
rect 22776 14868 22832 14870
rect 22880 14922 22936 14924
rect 22880 14870 22882 14922
rect 22882 14870 22934 14922
rect 22934 14870 22936 14922
rect 22880 14868 22936 14870
rect 22652 14530 22708 14532
rect 22652 14478 22654 14530
rect 22654 14478 22706 14530
rect 22706 14478 22708 14530
rect 22652 14476 22708 14478
rect 23212 15314 23268 15316
rect 23212 15262 23214 15314
rect 23214 15262 23266 15314
rect 23266 15262 23268 15314
rect 23212 15260 23268 15262
rect 23100 14476 23156 14532
rect 23660 17724 23716 17780
rect 23660 15932 23716 15988
rect 23436 14924 23492 14980
rect 22988 14306 23044 14308
rect 22988 14254 22990 14306
rect 22990 14254 23042 14306
rect 23042 14254 23044 14306
rect 22988 14252 23044 14254
rect 22092 13132 22148 13188
rect 22672 13354 22728 13356
rect 22672 13302 22674 13354
rect 22674 13302 22726 13354
rect 22726 13302 22728 13354
rect 22672 13300 22728 13302
rect 22776 13354 22832 13356
rect 22776 13302 22778 13354
rect 22778 13302 22830 13354
rect 22830 13302 22832 13354
rect 22776 13300 22832 13302
rect 22880 13354 22936 13356
rect 22880 13302 22882 13354
rect 22882 13302 22934 13354
rect 22934 13302 22936 13354
rect 22880 13300 22936 13302
rect 23548 13916 23604 13972
rect 23436 13746 23492 13748
rect 23436 13694 23438 13746
rect 23438 13694 23490 13746
rect 23490 13694 23492 13746
rect 23436 13692 23492 13694
rect 21868 12572 21924 12628
rect 22204 12738 22260 12740
rect 22204 12686 22206 12738
rect 22206 12686 22258 12738
rect 22258 12686 22260 12738
rect 22204 12684 22260 12686
rect 21980 12236 22036 12292
rect 21756 11900 21812 11956
rect 21980 11394 22036 11396
rect 21980 11342 21982 11394
rect 21982 11342 22034 11394
rect 22034 11342 22036 11394
rect 21980 11340 22036 11342
rect 22428 12684 22484 12740
rect 22428 12290 22484 12292
rect 22428 12238 22430 12290
rect 22430 12238 22482 12290
rect 22482 12238 22484 12290
rect 22428 12236 22484 12238
rect 23436 12572 23492 12628
rect 23212 11954 23268 11956
rect 23212 11902 23214 11954
rect 23214 11902 23266 11954
rect 23266 11902 23268 11954
rect 23212 11900 23268 11902
rect 22540 11788 22596 11844
rect 22672 11786 22728 11788
rect 22672 11734 22674 11786
rect 22674 11734 22726 11786
rect 22726 11734 22728 11786
rect 22672 11732 22728 11734
rect 22776 11786 22832 11788
rect 22776 11734 22778 11786
rect 22778 11734 22830 11786
rect 22830 11734 22832 11786
rect 22776 11732 22832 11734
rect 22880 11786 22936 11788
rect 22880 11734 22882 11786
rect 22882 11734 22934 11786
rect 22934 11734 22936 11786
rect 22880 11732 22936 11734
rect 22764 11340 22820 11396
rect 22204 11228 22260 11284
rect 22876 11282 22932 11284
rect 22876 11230 22878 11282
rect 22878 11230 22930 11282
rect 22930 11230 22932 11282
rect 22876 11228 22932 11230
rect 22764 10722 22820 10724
rect 22764 10670 22766 10722
rect 22766 10670 22818 10722
rect 22818 10670 22820 10722
rect 22764 10668 22820 10670
rect 20748 10220 20804 10276
rect 21644 10220 21700 10276
rect 21980 10444 22036 10500
rect 21532 9714 21588 9716
rect 21532 9662 21534 9714
rect 21534 9662 21586 9714
rect 21586 9662 21588 9714
rect 21532 9660 21588 9662
rect 20860 9324 20916 9380
rect 20860 7868 20916 7924
rect 20076 7420 20132 7476
rect 19852 7362 19908 7364
rect 19852 7310 19854 7362
rect 19854 7310 19906 7362
rect 19906 7310 19908 7362
rect 19852 7308 19908 7310
rect 19964 7084 20020 7140
rect 20188 7644 20244 7700
rect 20860 7644 20916 7700
rect 20188 7196 20244 7252
rect 20860 7362 20916 7364
rect 20860 7310 20862 7362
rect 20862 7310 20914 7362
rect 20914 7310 20916 7362
rect 20860 7308 20916 7310
rect 20524 6690 20580 6692
rect 20524 6638 20526 6690
rect 20526 6638 20578 6690
rect 20578 6638 20580 6690
rect 20524 6636 20580 6638
rect 22316 10444 22372 10500
rect 22876 10444 22932 10500
rect 22988 10892 23044 10948
rect 22988 10332 23044 10388
rect 23324 10892 23380 10948
rect 23548 12178 23604 12180
rect 23548 12126 23550 12178
rect 23550 12126 23602 12178
rect 23602 12126 23604 12178
rect 23548 12124 23604 12126
rect 23436 10780 23492 10836
rect 23212 10332 23268 10388
rect 22672 10218 22728 10220
rect 22672 10166 22674 10218
rect 22674 10166 22726 10218
rect 22726 10166 22728 10218
rect 22672 10164 22728 10166
rect 22776 10218 22832 10220
rect 22776 10166 22778 10218
rect 22778 10166 22830 10218
rect 22830 10166 22832 10218
rect 22776 10164 22832 10166
rect 22880 10218 22936 10220
rect 22880 10166 22882 10218
rect 22882 10166 22934 10218
rect 22934 10166 22936 10218
rect 22880 10164 22936 10166
rect 22988 9772 23044 9828
rect 21644 8764 21700 8820
rect 21308 6972 21364 7028
rect 21084 6860 21140 6916
rect 20636 6412 20692 6468
rect 20412 6076 20468 6132
rect 20300 5234 20356 5236
rect 20300 5182 20302 5234
rect 20302 5182 20354 5234
rect 20354 5182 20356 5234
rect 20300 5180 20356 5182
rect 19852 4284 19908 4340
rect 20412 4284 20468 4340
rect 19852 3554 19908 3556
rect 19852 3502 19854 3554
rect 19854 3502 19906 3554
rect 19906 3502 19908 3554
rect 19852 3500 19908 3502
rect 18396 2604 18452 2660
rect 21084 4844 21140 4900
rect 20972 4450 21028 4452
rect 20972 4398 20974 4450
rect 20974 4398 21026 4450
rect 21026 4398 21028 4450
rect 20972 4396 21028 4398
rect 20860 4338 20916 4340
rect 20860 4286 20862 4338
rect 20862 4286 20914 4338
rect 20914 4286 20916 4338
rect 20860 4284 20916 4286
rect 20972 4226 21028 4228
rect 20972 4174 20974 4226
rect 20974 4174 21026 4226
rect 21026 4174 21028 4226
rect 20972 4172 21028 4174
rect 21756 8034 21812 8036
rect 21756 7982 21758 8034
rect 21758 7982 21810 8034
rect 21810 7982 21812 8034
rect 21756 7980 21812 7982
rect 21644 7420 21700 7476
rect 22876 9660 22932 9716
rect 25452 18956 25508 19012
rect 24668 18674 24724 18676
rect 24668 18622 24670 18674
rect 24670 18622 24722 18674
rect 24722 18622 24724 18674
rect 24668 18620 24724 18622
rect 24780 18508 24836 18564
rect 24220 17724 24276 17780
rect 24556 17500 24612 17556
rect 25788 18620 25844 18676
rect 26348 19010 26404 19012
rect 26348 18958 26350 19010
rect 26350 18958 26402 19010
rect 26402 18958 26404 19010
rect 26348 18956 26404 18958
rect 26684 19068 26740 19124
rect 26908 19122 26964 19124
rect 26908 19070 26910 19122
rect 26910 19070 26962 19122
rect 26962 19070 26964 19122
rect 26908 19068 26964 19070
rect 26684 18562 26740 18564
rect 26684 18510 26686 18562
rect 26686 18510 26738 18562
rect 26738 18510 26740 18562
rect 26684 18508 26740 18510
rect 26796 17500 26852 17556
rect 25900 17388 25956 17444
rect 24108 16492 24164 16548
rect 24444 16268 24500 16324
rect 24332 16156 24388 16212
rect 24108 15314 24164 15316
rect 24108 15262 24110 15314
rect 24110 15262 24162 15314
rect 24162 15262 24164 15314
rect 24108 15260 24164 15262
rect 23884 13858 23940 13860
rect 23884 13806 23886 13858
rect 23886 13806 23938 13858
rect 23938 13806 23940 13858
rect 23884 13804 23940 13806
rect 24220 13692 24276 13748
rect 23884 12738 23940 12740
rect 23884 12686 23886 12738
rect 23886 12686 23938 12738
rect 23938 12686 23940 12738
rect 23884 12684 23940 12686
rect 25340 16940 25396 16996
rect 24780 16882 24836 16884
rect 24780 16830 24782 16882
rect 24782 16830 24834 16882
rect 24834 16830 24836 16882
rect 24780 16828 24836 16830
rect 25676 16882 25732 16884
rect 25676 16830 25678 16882
rect 25678 16830 25730 16882
rect 25730 16830 25732 16882
rect 25676 16828 25732 16830
rect 25452 16716 25508 16772
rect 25340 16492 25396 16548
rect 25116 16210 25172 16212
rect 25116 16158 25118 16210
rect 25118 16158 25170 16210
rect 25170 16158 25172 16210
rect 25116 16156 25172 16158
rect 24780 15820 24836 15876
rect 24444 13468 24500 13524
rect 24556 14476 24612 14532
rect 24332 12178 24388 12180
rect 24332 12126 24334 12178
rect 24334 12126 24386 12178
rect 24386 12126 24388 12178
rect 24332 12124 24388 12126
rect 24668 14252 24724 14308
rect 25116 15148 25172 15204
rect 25340 15820 25396 15876
rect 25452 15314 25508 15316
rect 25452 15262 25454 15314
rect 25454 15262 25506 15314
rect 25506 15262 25508 15314
rect 25452 15260 25508 15262
rect 25452 14530 25508 14532
rect 25452 14478 25454 14530
rect 25454 14478 25506 14530
rect 25506 14478 25508 14530
rect 25452 14476 25508 14478
rect 25228 14306 25284 14308
rect 25228 14254 25230 14306
rect 25230 14254 25282 14306
rect 25282 14254 25284 14306
rect 25228 14252 25284 14254
rect 26908 16044 26964 16100
rect 26012 15148 26068 15204
rect 26348 15874 26404 15876
rect 26348 15822 26350 15874
rect 26350 15822 26402 15874
rect 26402 15822 26404 15874
rect 26348 15820 26404 15822
rect 26124 15484 26180 15540
rect 25900 14812 25956 14868
rect 26124 14588 26180 14644
rect 26572 14588 26628 14644
rect 26460 14306 26516 14308
rect 26460 14254 26462 14306
rect 26462 14254 26514 14306
rect 26514 14254 26516 14306
rect 26460 14252 26516 14254
rect 26572 14364 26628 14420
rect 25788 14028 25844 14084
rect 26348 14028 26404 14084
rect 25228 13970 25284 13972
rect 25228 13918 25230 13970
rect 25230 13918 25282 13970
rect 25282 13918 25284 13970
rect 25228 13916 25284 13918
rect 24668 13804 24724 13860
rect 24668 12962 24724 12964
rect 24668 12910 24670 12962
rect 24670 12910 24722 12962
rect 24722 12910 24724 12962
rect 24668 12908 24724 12910
rect 24780 13468 24836 13524
rect 24892 13356 24948 13412
rect 25676 12962 25732 12964
rect 25676 12910 25678 12962
rect 25678 12910 25730 12962
rect 25730 12910 25732 12962
rect 25676 12908 25732 12910
rect 24556 12290 24612 12292
rect 24556 12238 24558 12290
rect 24558 12238 24610 12290
rect 24610 12238 24612 12290
rect 24556 12236 24612 12238
rect 24444 12012 24500 12068
rect 23772 10610 23828 10612
rect 23772 10558 23774 10610
rect 23774 10558 23826 10610
rect 23826 10558 23828 10610
rect 23772 10556 23828 10558
rect 23660 9996 23716 10052
rect 23660 9826 23716 9828
rect 23660 9774 23662 9826
rect 23662 9774 23714 9826
rect 23714 9774 23716 9826
rect 23660 9772 23716 9774
rect 23324 9548 23380 9604
rect 23100 9154 23156 9156
rect 23100 9102 23102 9154
rect 23102 9102 23154 9154
rect 23154 9102 23156 9154
rect 23100 9100 23156 9102
rect 23436 8930 23492 8932
rect 23436 8878 23438 8930
rect 23438 8878 23490 8930
rect 23490 8878 23492 8930
rect 23436 8876 23492 8878
rect 22672 8650 22728 8652
rect 22672 8598 22674 8650
rect 22674 8598 22726 8650
rect 22726 8598 22728 8650
rect 22672 8596 22728 8598
rect 22776 8650 22832 8652
rect 22776 8598 22778 8650
rect 22778 8598 22830 8650
rect 22830 8598 22832 8650
rect 22776 8596 22832 8598
rect 22880 8650 22936 8652
rect 22880 8598 22882 8650
rect 22882 8598 22934 8650
rect 22934 8598 22936 8650
rect 22880 8596 22936 8598
rect 22764 8258 22820 8260
rect 22764 8206 22766 8258
rect 22766 8206 22818 8258
rect 22818 8206 22820 8258
rect 22764 8204 22820 8206
rect 23100 8092 23156 8148
rect 23324 8428 23380 8484
rect 23100 7644 23156 7700
rect 22988 7474 23044 7476
rect 22988 7422 22990 7474
rect 22990 7422 23042 7474
rect 23042 7422 23044 7474
rect 22988 7420 23044 7422
rect 22672 7082 22728 7084
rect 21868 6972 21924 7028
rect 22672 7030 22674 7082
rect 22674 7030 22726 7082
rect 22726 7030 22728 7082
rect 22672 7028 22728 7030
rect 22776 7082 22832 7084
rect 22776 7030 22778 7082
rect 22778 7030 22830 7082
rect 22830 7030 22832 7082
rect 22776 7028 22832 7030
rect 22880 7082 22936 7084
rect 22880 7030 22882 7082
rect 22882 7030 22934 7082
rect 22934 7030 22936 7082
rect 22880 7028 22936 7030
rect 22764 6860 22820 6916
rect 22428 6412 22484 6468
rect 21420 3724 21476 3780
rect 22316 4620 22372 4676
rect 21980 4338 22036 4340
rect 21980 4286 21982 4338
rect 21982 4286 22034 4338
rect 22034 4286 22036 4338
rect 21980 4284 22036 4286
rect 22316 3948 22372 4004
rect 20748 2492 20804 2548
rect 22652 6076 22708 6132
rect 22672 5514 22728 5516
rect 22672 5462 22674 5514
rect 22674 5462 22726 5514
rect 22726 5462 22728 5514
rect 22672 5460 22728 5462
rect 22776 5514 22832 5516
rect 22776 5462 22778 5514
rect 22778 5462 22830 5514
rect 22830 5462 22832 5514
rect 22776 5460 22832 5462
rect 22880 5514 22936 5516
rect 22880 5462 22882 5514
rect 22882 5462 22934 5514
rect 22934 5462 22936 5514
rect 22880 5460 22936 5462
rect 22540 5180 22596 5236
rect 22764 5292 22820 5348
rect 22652 4508 22708 4564
rect 23100 5068 23156 5124
rect 22876 4226 22932 4228
rect 22876 4174 22878 4226
rect 22878 4174 22930 4226
rect 22930 4174 22932 4226
rect 22876 4172 22932 4174
rect 22672 3946 22728 3948
rect 22672 3894 22674 3946
rect 22674 3894 22726 3946
rect 22726 3894 22728 3946
rect 22672 3892 22728 3894
rect 22776 3946 22832 3948
rect 22776 3894 22778 3946
rect 22778 3894 22830 3946
rect 22830 3894 22832 3946
rect 22776 3892 22832 3894
rect 22880 3946 22936 3948
rect 22880 3894 22882 3946
rect 22882 3894 22934 3946
rect 22934 3894 22936 3946
rect 22880 3892 22936 3894
rect 23772 8092 23828 8148
rect 23436 6076 23492 6132
rect 23548 6524 23604 6580
rect 23324 5516 23380 5572
rect 24556 11394 24612 11396
rect 24556 11342 24558 11394
rect 24558 11342 24610 11394
rect 24610 11342 24612 11394
rect 24556 11340 24612 11342
rect 24332 9884 24388 9940
rect 24556 9154 24612 9156
rect 24556 9102 24558 9154
rect 24558 9102 24610 9154
rect 24610 9102 24612 9154
rect 24556 9100 24612 9102
rect 24108 9042 24164 9044
rect 24108 8990 24110 9042
rect 24110 8990 24162 9042
rect 24162 8990 24164 9042
rect 24108 8988 24164 8990
rect 23996 8764 24052 8820
rect 24108 8428 24164 8484
rect 23884 7532 23940 7588
rect 24668 6130 24724 6132
rect 24668 6078 24670 6130
rect 24670 6078 24722 6130
rect 24722 6078 24724 6130
rect 24668 6076 24724 6078
rect 24332 5068 24388 5124
rect 24780 5852 24836 5908
rect 23212 4956 23268 5012
rect 23996 4844 24052 4900
rect 24332 4562 24388 4564
rect 24332 4510 24334 4562
rect 24334 4510 24386 4562
rect 24386 4510 24388 4562
rect 24332 4508 24388 4510
rect 25116 12850 25172 12852
rect 25116 12798 25118 12850
rect 25118 12798 25170 12850
rect 25170 12798 25172 12850
rect 25116 12796 25172 12798
rect 25340 12236 25396 12292
rect 25900 12796 25956 12852
rect 25900 12124 25956 12180
rect 25228 11394 25284 11396
rect 25228 11342 25230 11394
rect 25230 11342 25282 11394
rect 25282 11342 25284 11394
rect 25228 11340 25284 11342
rect 25340 10834 25396 10836
rect 25340 10782 25342 10834
rect 25342 10782 25394 10834
rect 25394 10782 25396 10834
rect 25340 10780 25396 10782
rect 25228 9996 25284 10052
rect 25676 11282 25732 11284
rect 25676 11230 25678 11282
rect 25678 11230 25730 11282
rect 25730 11230 25732 11282
rect 25676 11228 25732 11230
rect 26236 12962 26292 12964
rect 26236 12910 26238 12962
rect 26238 12910 26290 12962
rect 26290 12910 26292 12962
rect 26236 12908 26292 12910
rect 26684 14140 26740 14196
rect 26908 13132 26964 13188
rect 26796 12460 26852 12516
rect 26012 11452 26068 11508
rect 26124 12066 26180 12068
rect 26124 12014 26126 12066
rect 26126 12014 26178 12066
rect 26178 12014 26180 12066
rect 26124 12012 26180 12014
rect 26236 11900 26292 11956
rect 26460 12012 26516 12068
rect 26124 10834 26180 10836
rect 26124 10782 26126 10834
rect 26126 10782 26178 10834
rect 26178 10782 26180 10834
rect 26124 10780 26180 10782
rect 26124 9996 26180 10052
rect 26012 9938 26068 9940
rect 26012 9886 26014 9938
rect 26014 9886 26066 9938
rect 26066 9886 26068 9938
rect 26012 9884 26068 9886
rect 25900 9436 25956 9492
rect 26124 8988 26180 9044
rect 25900 8876 25956 8932
rect 26348 10892 26404 10948
rect 26684 11452 26740 11508
rect 25788 8764 25844 8820
rect 25676 8652 25732 8708
rect 25228 8316 25284 8372
rect 25228 6300 25284 6356
rect 24892 4508 24948 4564
rect 25004 5068 25060 5124
rect 23996 3666 24052 3668
rect 23996 3614 23998 3666
rect 23998 3614 24050 3666
rect 24050 3614 24052 3666
rect 23996 3612 24052 3614
rect 25116 4844 25172 4900
rect 25228 5404 25284 5460
rect 25564 8370 25620 8372
rect 25564 8318 25566 8370
rect 25566 8318 25618 8370
rect 25618 8318 25620 8370
rect 25564 8316 25620 8318
rect 25900 8258 25956 8260
rect 25900 8206 25902 8258
rect 25902 8206 25954 8258
rect 25954 8206 25956 8258
rect 25900 8204 25956 8206
rect 26348 8652 26404 8708
rect 27020 12460 27076 12516
rect 27692 23714 27748 23716
rect 27692 23662 27694 23714
rect 27694 23662 27746 23714
rect 27746 23662 27748 23714
rect 27692 23660 27748 23662
rect 28028 23714 28084 23716
rect 28028 23662 28030 23714
rect 28030 23662 28082 23714
rect 28082 23662 28084 23714
rect 28028 23660 28084 23662
rect 27916 23548 27972 23604
rect 28028 23324 28084 23380
rect 28588 23938 28644 23940
rect 28588 23886 28590 23938
rect 28590 23886 28642 23938
rect 28642 23886 28644 23938
rect 28588 23884 28644 23886
rect 27804 23042 27860 23044
rect 27804 22990 27806 23042
rect 27806 22990 27858 23042
rect 27858 22990 27860 23042
rect 27804 22988 27860 22990
rect 27244 22652 27300 22708
rect 27356 22876 27412 22932
rect 27356 22540 27412 22596
rect 27580 22204 27636 22260
rect 28028 21420 28084 21476
rect 28028 21084 28084 21140
rect 28140 20076 28196 20132
rect 28028 19964 28084 20020
rect 28588 22370 28644 22372
rect 28588 22318 28590 22370
rect 28590 22318 28642 22370
rect 28642 22318 28644 22370
rect 28588 22316 28644 22318
rect 28588 22092 28644 22148
rect 28812 23772 28868 23828
rect 29260 28476 29316 28532
rect 29260 26962 29316 26964
rect 29260 26910 29262 26962
rect 29262 26910 29314 26962
rect 29314 26910 29316 26962
rect 29260 26908 29316 26910
rect 29148 25506 29204 25508
rect 29148 25454 29150 25506
rect 29150 25454 29202 25506
rect 29202 25454 29204 25506
rect 29148 25452 29204 25454
rect 29148 25004 29204 25060
rect 29372 27468 29428 27524
rect 29825 29818 29881 29820
rect 29825 29766 29827 29818
rect 29827 29766 29879 29818
rect 29879 29766 29881 29818
rect 29825 29764 29881 29766
rect 29929 29818 29985 29820
rect 29929 29766 29931 29818
rect 29931 29766 29983 29818
rect 29983 29766 29985 29818
rect 29929 29764 29985 29766
rect 30033 29818 30089 29820
rect 30033 29766 30035 29818
rect 30035 29766 30087 29818
rect 30087 29766 30089 29818
rect 30033 29764 30089 29766
rect 31388 30210 31444 30212
rect 31388 30158 31390 30210
rect 31390 30158 31442 30210
rect 31442 30158 31444 30210
rect 31388 30156 31444 30158
rect 30604 29426 30660 29428
rect 30604 29374 30606 29426
rect 30606 29374 30658 29426
rect 30658 29374 30660 29426
rect 30604 29372 30660 29374
rect 29825 28250 29881 28252
rect 29825 28198 29827 28250
rect 29827 28198 29879 28250
rect 29879 28198 29881 28250
rect 29825 28196 29881 28198
rect 29929 28250 29985 28252
rect 29929 28198 29931 28250
rect 29931 28198 29983 28250
rect 29983 28198 29985 28250
rect 29929 28196 29985 28198
rect 30033 28250 30089 28252
rect 30033 28198 30035 28250
rect 30035 28198 30087 28250
rect 30087 28198 30089 28250
rect 30033 28196 30089 28198
rect 33292 31778 33348 31780
rect 33292 31726 33294 31778
rect 33294 31726 33346 31778
rect 33346 31726 33348 31778
rect 33292 31724 33348 31726
rect 32508 31554 32564 31556
rect 32508 31502 32510 31554
rect 32510 31502 32562 31554
rect 32562 31502 32564 31554
rect 32508 31500 32564 31502
rect 31836 31164 31892 31220
rect 33404 31666 33460 31668
rect 33404 31614 33406 31666
rect 33406 31614 33458 31666
rect 33458 31614 33460 31666
rect 33404 31612 33460 31614
rect 33292 31106 33348 31108
rect 33292 31054 33294 31106
rect 33294 31054 33346 31106
rect 33346 31054 33348 31106
rect 33292 31052 33348 31054
rect 31836 30492 31892 30548
rect 31612 30268 31668 30324
rect 31948 30156 32004 30212
rect 32396 30604 32452 30660
rect 32060 30044 32116 30100
rect 31948 29708 32004 29764
rect 33068 29708 33124 29764
rect 32396 29650 32452 29652
rect 32396 29598 32398 29650
rect 32398 29598 32450 29650
rect 32450 29598 32452 29650
rect 32396 29596 32452 29598
rect 32956 29596 33012 29652
rect 31612 29426 31668 29428
rect 31612 29374 31614 29426
rect 31614 29374 31666 29426
rect 31666 29374 31668 29426
rect 31612 29372 31668 29374
rect 32172 29426 32228 29428
rect 32172 29374 32174 29426
rect 32174 29374 32226 29426
rect 32226 29374 32228 29426
rect 32172 29372 32228 29374
rect 31612 28812 31668 28868
rect 31276 27692 31332 27748
rect 30044 26850 30100 26852
rect 30044 26798 30046 26850
rect 30046 26798 30098 26850
rect 30098 26798 30100 26850
rect 30044 26796 30100 26798
rect 29825 26682 29881 26684
rect 29825 26630 29827 26682
rect 29827 26630 29879 26682
rect 29879 26630 29881 26682
rect 29825 26628 29881 26630
rect 29929 26682 29985 26684
rect 29929 26630 29931 26682
rect 29931 26630 29983 26682
rect 29983 26630 29985 26682
rect 29929 26628 29985 26630
rect 30033 26682 30089 26684
rect 30033 26630 30035 26682
rect 30035 26630 30087 26682
rect 30087 26630 30089 26682
rect 30033 26628 30089 26630
rect 30044 25228 30100 25284
rect 30156 25452 30212 25508
rect 29596 25116 29652 25172
rect 29260 24722 29316 24724
rect 29260 24670 29262 24722
rect 29262 24670 29314 24722
rect 29314 24670 29316 24722
rect 29260 24668 29316 24670
rect 29825 25114 29881 25116
rect 29825 25062 29827 25114
rect 29827 25062 29879 25114
rect 29879 25062 29881 25114
rect 29825 25060 29881 25062
rect 29929 25114 29985 25116
rect 29929 25062 29931 25114
rect 29931 25062 29983 25114
rect 29983 25062 29985 25114
rect 29929 25060 29985 25062
rect 30033 25114 30089 25116
rect 30033 25062 30035 25114
rect 30035 25062 30087 25114
rect 30087 25062 30089 25114
rect 30033 25060 30089 25062
rect 29708 24668 29764 24724
rect 29820 24444 29876 24500
rect 29260 23548 29316 23604
rect 28476 20802 28532 20804
rect 28476 20750 28478 20802
rect 28478 20750 28530 20802
rect 28530 20750 28532 20802
rect 28476 20748 28532 20750
rect 28364 19964 28420 20020
rect 28140 19906 28196 19908
rect 28140 19854 28142 19906
rect 28142 19854 28194 19906
rect 28194 19854 28196 19906
rect 28140 19852 28196 19854
rect 28700 20018 28756 20020
rect 28700 19966 28702 20018
rect 28702 19966 28754 20018
rect 28754 19966 28756 20018
rect 28700 19964 28756 19966
rect 28140 19068 28196 19124
rect 28476 19234 28532 19236
rect 28476 19182 28478 19234
rect 28478 19182 28530 19234
rect 28530 19182 28532 19234
rect 28476 19180 28532 19182
rect 27916 18172 27972 18228
rect 28028 18284 28084 18340
rect 28476 18284 28532 18340
rect 27916 17666 27972 17668
rect 27916 17614 27918 17666
rect 27918 17614 27970 17666
rect 27970 17614 27972 17666
rect 27916 17612 27972 17614
rect 27356 16658 27412 16660
rect 27356 16606 27358 16658
rect 27358 16606 27410 16658
rect 27410 16606 27412 16658
rect 27356 16604 27412 16606
rect 28476 16604 28532 16660
rect 27244 15820 27300 15876
rect 27580 16044 27636 16100
rect 28252 16098 28308 16100
rect 28252 16046 28254 16098
rect 28254 16046 28306 16098
rect 28306 16046 28308 16098
rect 28252 16044 28308 16046
rect 27356 15148 27412 15204
rect 27580 15426 27636 15428
rect 27580 15374 27582 15426
rect 27582 15374 27634 15426
rect 27634 15374 27636 15426
rect 27580 15372 27636 15374
rect 27356 14028 27412 14084
rect 27132 12908 27188 12964
rect 27132 12290 27188 12292
rect 27132 12238 27134 12290
rect 27134 12238 27186 12290
rect 27186 12238 27188 12290
rect 27132 12236 27188 12238
rect 27020 12012 27076 12068
rect 26908 11788 26964 11844
rect 27020 11564 27076 11620
rect 26908 11394 26964 11396
rect 26908 11342 26910 11394
rect 26910 11342 26962 11394
rect 26962 11342 26964 11394
rect 26908 11340 26964 11342
rect 27132 11394 27188 11396
rect 27132 11342 27134 11394
rect 27134 11342 27186 11394
rect 27186 11342 27188 11394
rect 27132 11340 27188 11342
rect 27468 12684 27524 12740
rect 27580 12066 27636 12068
rect 27580 12014 27582 12066
rect 27582 12014 27634 12066
rect 27634 12014 27636 12066
rect 27580 12012 27636 12014
rect 28140 15596 28196 15652
rect 28028 15426 28084 15428
rect 28028 15374 28030 15426
rect 28030 15374 28082 15426
rect 28082 15374 28084 15426
rect 28028 15372 28084 15374
rect 27916 15314 27972 15316
rect 27916 15262 27918 15314
rect 27918 15262 27970 15314
rect 27970 15262 27972 15314
rect 27916 15260 27972 15262
rect 27804 15036 27860 15092
rect 27804 14700 27860 14756
rect 27916 14418 27972 14420
rect 27916 14366 27918 14418
rect 27918 14366 27970 14418
rect 27970 14366 27972 14418
rect 27916 14364 27972 14366
rect 28028 12738 28084 12740
rect 28028 12686 28030 12738
rect 28030 12686 28082 12738
rect 28082 12686 28084 12738
rect 28028 12684 28084 12686
rect 27692 11788 27748 11844
rect 27804 12236 27860 12292
rect 27916 12178 27972 12180
rect 27916 12126 27918 12178
rect 27918 12126 27970 12178
rect 27970 12126 27972 12178
rect 27916 12124 27972 12126
rect 27356 11170 27412 11172
rect 27356 11118 27358 11170
rect 27358 11118 27410 11170
rect 27410 11118 27412 11170
rect 27356 11116 27412 11118
rect 27244 10892 27300 10948
rect 27020 10668 27076 10724
rect 27132 10780 27188 10836
rect 27020 9826 27076 9828
rect 27020 9774 27022 9826
rect 27022 9774 27074 9826
rect 27074 9774 27076 9826
rect 27020 9772 27076 9774
rect 26460 9660 26516 9716
rect 26124 8092 26180 8148
rect 25564 7196 25620 7252
rect 26236 7196 26292 7252
rect 25788 6636 25844 6692
rect 26124 6524 26180 6580
rect 26012 5906 26068 5908
rect 26012 5854 26014 5906
rect 26014 5854 26066 5906
rect 26066 5854 26068 5906
rect 26012 5852 26068 5854
rect 25788 5404 25844 5460
rect 26236 5628 26292 5684
rect 25676 5292 25732 5348
rect 25452 4844 25508 4900
rect 25452 4620 25508 4676
rect 25564 4396 25620 4452
rect 25676 4620 25732 4676
rect 25004 3554 25060 3556
rect 25004 3502 25006 3554
rect 25006 3502 25058 3554
rect 25058 3502 25060 3554
rect 25004 3500 25060 3502
rect 25676 3442 25732 3444
rect 25676 3390 25678 3442
rect 25678 3390 25730 3442
rect 25730 3390 25732 3442
rect 25676 3388 25732 3390
rect 27356 10722 27412 10724
rect 27356 10670 27358 10722
rect 27358 10670 27410 10722
rect 27410 10670 27412 10722
rect 27356 10668 27412 10670
rect 27356 10108 27412 10164
rect 27020 9548 27076 9604
rect 26684 9100 26740 9156
rect 26460 5964 26516 6020
rect 26572 7756 26628 7812
rect 26908 9324 26964 9380
rect 26796 8818 26852 8820
rect 26796 8766 26798 8818
rect 26798 8766 26850 8818
rect 26850 8766 26852 8818
rect 26796 8764 26852 8766
rect 27132 9212 27188 9268
rect 27132 7980 27188 8036
rect 27916 9548 27972 9604
rect 27804 9436 27860 9492
rect 29596 23884 29652 23940
rect 28924 23378 28980 23380
rect 28924 23326 28926 23378
rect 28926 23326 28978 23378
rect 28978 23326 28980 23378
rect 28924 23324 28980 23326
rect 29260 22930 29316 22932
rect 29260 22878 29262 22930
rect 29262 22878 29314 22930
rect 29314 22878 29316 22930
rect 29260 22876 29316 22878
rect 29260 22316 29316 22372
rect 29036 22092 29092 22148
rect 29148 21420 29204 21476
rect 30828 26908 30884 26964
rect 30492 26236 30548 26292
rect 30268 25340 30324 25396
rect 30268 24444 30324 24500
rect 30492 26012 30548 26068
rect 29825 23546 29881 23548
rect 29825 23494 29827 23546
rect 29827 23494 29879 23546
rect 29879 23494 29881 23546
rect 29825 23492 29881 23494
rect 29929 23546 29985 23548
rect 29929 23494 29931 23546
rect 29931 23494 29983 23546
rect 29983 23494 29985 23546
rect 29929 23492 29985 23494
rect 30033 23546 30089 23548
rect 30033 23494 30035 23546
rect 30035 23494 30087 23546
rect 30087 23494 30089 23546
rect 30033 23492 30089 23494
rect 30156 23100 30212 23156
rect 30268 23042 30324 23044
rect 30268 22990 30270 23042
rect 30270 22990 30322 23042
rect 30322 22990 30324 23042
rect 30268 22988 30324 22990
rect 29372 21532 29428 21588
rect 29596 21420 29652 21476
rect 29825 21978 29881 21980
rect 29825 21926 29827 21978
rect 29827 21926 29879 21978
rect 29879 21926 29881 21978
rect 29825 21924 29881 21926
rect 29929 21978 29985 21980
rect 29929 21926 29931 21978
rect 29931 21926 29983 21978
rect 29983 21926 29985 21978
rect 29929 21924 29985 21926
rect 30033 21978 30089 21980
rect 30033 21926 30035 21978
rect 30035 21926 30087 21978
rect 30087 21926 30089 21978
rect 30033 21924 30089 21926
rect 29260 20690 29316 20692
rect 29260 20638 29262 20690
rect 29262 20638 29314 20690
rect 29314 20638 29316 20690
rect 29260 20636 29316 20638
rect 30268 21532 30324 21588
rect 30940 26402 30996 26404
rect 30940 26350 30942 26402
rect 30942 26350 30994 26402
rect 30994 26350 30996 26402
rect 30940 26348 30996 26350
rect 32172 27692 32228 27748
rect 32060 26962 32116 26964
rect 32060 26910 32062 26962
rect 32062 26910 32114 26962
rect 32114 26910 32116 26962
rect 32060 26908 32116 26910
rect 30716 25506 30772 25508
rect 30716 25454 30718 25506
rect 30718 25454 30770 25506
rect 30770 25454 30772 25506
rect 30716 25452 30772 25454
rect 30604 25116 30660 25172
rect 30492 24834 30548 24836
rect 30492 24782 30494 24834
rect 30494 24782 30546 24834
rect 30546 24782 30548 24834
rect 30492 24780 30548 24782
rect 30940 24668 30996 24724
rect 30716 24556 30772 24612
rect 30604 23324 30660 23380
rect 30492 23266 30548 23268
rect 30492 23214 30494 23266
rect 30494 23214 30546 23266
rect 30546 23214 30548 23266
rect 30492 23212 30548 23214
rect 30604 22652 30660 22708
rect 30604 22258 30660 22260
rect 30604 22206 30606 22258
rect 30606 22206 30658 22258
rect 30658 22206 30660 22258
rect 30604 22204 30660 22206
rect 30492 21420 30548 21476
rect 30492 20860 30548 20916
rect 30828 23154 30884 23156
rect 30828 23102 30830 23154
rect 30830 23102 30882 23154
rect 30882 23102 30884 23154
rect 30828 23100 30884 23102
rect 30940 22540 30996 22596
rect 30828 22428 30884 22484
rect 30940 21532 30996 21588
rect 30156 20748 30212 20804
rect 29825 20410 29881 20412
rect 29825 20358 29827 20410
rect 29827 20358 29879 20410
rect 29879 20358 29881 20410
rect 29825 20356 29881 20358
rect 29929 20410 29985 20412
rect 29929 20358 29931 20410
rect 29931 20358 29983 20410
rect 29983 20358 29985 20410
rect 29929 20356 29985 20358
rect 30033 20410 30089 20412
rect 30033 20358 30035 20410
rect 30035 20358 30087 20410
rect 30087 20358 30089 20410
rect 30033 20356 30089 20358
rect 29708 20188 29764 20244
rect 30716 20636 30772 20692
rect 30156 20018 30212 20020
rect 30156 19966 30158 20018
rect 30158 19966 30210 20018
rect 30210 19966 30212 20018
rect 30156 19964 30212 19966
rect 29932 19404 29988 19460
rect 29260 19346 29316 19348
rect 29260 19294 29262 19346
rect 29262 19294 29314 19346
rect 29314 19294 29316 19346
rect 29260 19292 29316 19294
rect 30716 20076 30772 20132
rect 29036 19234 29092 19236
rect 29036 19182 29038 19234
rect 29038 19182 29090 19234
rect 29090 19182 29092 19234
rect 29036 19180 29092 19182
rect 29484 19122 29540 19124
rect 29484 19070 29486 19122
rect 29486 19070 29538 19122
rect 29538 19070 29540 19122
rect 29484 19068 29540 19070
rect 29825 18842 29881 18844
rect 29825 18790 29827 18842
rect 29827 18790 29879 18842
rect 29879 18790 29881 18842
rect 29825 18788 29881 18790
rect 29929 18842 29985 18844
rect 29929 18790 29931 18842
rect 29931 18790 29983 18842
rect 29983 18790 29985 18842
rect 29929 18788 29985 18790
rect 30033 18842 30089 18844
rect 30033 18790 30035 18842
rect 30035 18790 30087 18842
rect 30087 18790 30089 18842
rect 30033 18788 30089 18790
rect 30268 18844 30324 18900
rect 29260 18450 29316 18452
rect 29260 18398 29262 18450
rect 29262 18398 29314 18450
rect 29314 18398 29316 18450
rect 29260 18396 29316 18398
rect 29148 17836 29204 17892
rect 29148 17666 29204 17668
rect 29148 17614 29150 17666
rect 29150 17614 29202 17666
rect 29202 17614 29204 17666
rect 29148 17612 29204 17614
rect 29820 18450 29876 18452
rect 29820 18398 29822 18450
rect 29822 18398 29874 18450
rect 29874 18398 29876 18450
rect 29820 18396 29876 18398
rect 30380 18338 30436 18340
rect 30380 18286 30382 18338
rect 30382 18286 30434 18338
rect 30434 18286 30436 18338
rect 30380 18284 30436 18286
rect 30156 18060 30212 18116
rect 30044 17836 30100 17892
rect 29825 17274 29881 17276
rect 29825 17222 29827 17274
rect 29827 17222 29879 17274
rect 29879 17222 29881 17274
rect 29825 17220 29881 17222
rect 29929 17274 29985 17276
rect 29929 17222 29931 17274
rect 29931 17222 29983 17274
rect 29983 17222 29985 17274
rect 29929 17220 29985 17222
rect 30033 17274 30089 17276
rect 30033 17222 30035 17274
rect 30035 17222 30087 17274
rect 30087 17222 30089 17274
rect 30033 17220 30089 17222
rect 30604 18956 30660 19012
rect 30716 18396 30772 18452
rect 30604 18172 30660 18228
rect 31612 26290 31668 26292
rect 31612 26238 31614 26290
rect 31614 26238 31666 26290
rect 31666 26238 31668 26290
rect 31612 26236 31668 26238
rect 32060 26236 32116 26292
rect 31164 25506 31220 25508
rect 31164 25454 31166 25506
rect 31166 25454 31218 25506
rect 31218 25454 31220 25506
rect 31164 25452 31220 25454
rect 32284 26236 32340 26292
rect 32172 25452 32228 25508
rect 32956 28588 33012 28644
rect 33180 29372 33236 29428
rect 33292 28754 33348 28756
rect 33292 28702 33294 28754
rect 33294 28702 33346 28754
rect 33346 28702 33348 28754
rect 33292 28700 33348 28702
rect 33180 28642 33236 28644
rect 33180 28590 33182 28642
rect 33182 28590 33234 28642
rect 33234 28590 33236 28642
rect 33180 28588 33236 28590
rect 33852 31890 33908 31892
rect 33852 31838 33854 31890
rect 33854 31838 33906 31890
rect 33906 31838 33908 31890
rect 33852 31836 33908 31838
rect 33740 31724 33796 31780
rect 34972 31836 35028 31892
rect 34524 31612 34580 31668
rect 34412 31388 34468 31444
rect 34076 30994 34132 30996
rect 34076 30942 34078 30994
rect 34078 30942 34130 30994
rect 34130 30942 34132 30994
rect 34076 30940 34132 30942
rect 34636 29596 34692 29652
rect 33740 29148 33796 29204
rect 34524 29202 34580 29204
rect 34524 29150 34526 29202
rect 34526 29150 34578 29202
rect 34578 29150 34580 29202
rect 34524 29148 34580 29150
rect 33180 26572 33236 26628
rect 33292 26460 33348 26516
rect 33740 28642 33796 28644
rect 33740 28590 33742 28642
rect 33742 28590 33794 28642
rect 33794 28590 33796 28642
rect 33740 28588 33796 28590
rect 33740 27020 33796 27076
rect 34076 27074 34132 27076
rect 34076 27022 34078 27074
rect 34078 27022 34130 27074
rect 34130 27022 34132 27074
rect 34076 27020 34132 27022
rect 34636 27858 34692 27860
rect 34636 27806 34638 27858
rect 34638 27806 34690 27858
rect 34690 27806 34692 27858
rect 34636 27804 34692 27806
rect 34524 27580 34580 27636
rect 34860 27356 34916 27412
rect 34972 26962 35028 26964
rect 34972 26910 34974 26962
rect 34974 26910 35026 26962
rect 35026 26910 35028 26962
rect 34972 26908 35028 26910
rect 33964 26572 34020 26628
rect 33852 26460 33908 26516
rect 32844 25788 32900 25844
rect 33740 26402 33796 26404
rect 33740 26350 33742 26402
rect 33742 26350 33794 26402
rect 33794 26350 33796 26402
rect 33740 26348 33796 26350
rect 33180 25788 33236 25844
rect 34300 26402 34356 26404
rect 34300 26350 34302 26402
rect 34302 26350 34354 26402
rect 34354 26350 34356 26402
rect 34300 26348 34356 26350
rect 33180 25394 33236 25396
rect 33180 25342 33182 25394
rect 33182 25342 33234 25394
rect 33234 25342 33236 25394
rect 33180 25340 33236 25342
rect 32956 25228 33012 25284
rect 31500 24610 31556 24612
rect 31500 24558 31502 24610
rect 31502 24558 31554 24610
rect 31554 24558 31556 24610
rect 31500 24556 31556 24558
rect 32172 24722 32228 24724
rect 32172 24670 32174 24722
rect 32174 24670 32226 24722
rect 32226 24670 32228 24722
rect 32172 24668 32228 24670
rect 31724 23884 31780 23940
rect 31948 24220 32004 24276
rect 31388 23660 31444 23716
rect 31724 23324 31780 23380
rect 31164 22876 31220 22932
rect 31276 22652 31332 22708
rect 31500 23212 31556 23268
rect 31612 22876 31668 22932
rect 31836 22988 31892 23044
rect 31388 22258 31444 22260
rect 31388 22206 31390 22258
rect 31390 22206 31442 22258
rect 31442 22206 31444 22258
rect 31388 22204 31444 22206
rect 31612 21980 31668 22036
rect 31500 21532 31556 21588
rect 31164 21196 31220 21252
rect 32060 23772 32116 23828
rect 33404 24722 33460 24724
rect 33404 24670 33406 24722
rect 33406 24670 33458 24722
rect 33458 24670 33460 24722
rect 33404 24668 33460 24670
rect 33628 24892 33684 24948
rect 32396 23938 32452 23940
rect 32396 23886 32398 23938
rect 32398 23886 32450 23938
rect 32450 23886 32452 23938
rect 32396 23884 32452 23886
rect 32956 23938 33012 23940
rect 32956 23886 32958 23938
rect 32958 23886 33010 23938
rect 33010 23886 33012 23938
rect 32956 23884 33012 23886
rect 33068 23826 33124 23828
rect 33068 23774 33070 23826
rect 33070 23774 33122 23826
rect 33122 23774 33124 23826
rect 33068 23772 33124 23774
rect 32284 23660 32340 23716
rect 33292 23436 33348 23492
rect 32060 22876 32116 22932
rect 31948 22428 32004 22484
rect 31948 22092 32004 22148
rect 32508 22428 32564 22484
rect 32396 22316 32452 22372
rect 32620 22092 32676 22148
rect 32508 21756 32564 21812
rect 31948 21586 32004 21588
rect 31948 21534 31950 21586
rect 31950 21534 32002 21586
rect 32002 21534 32004 21586
rect 31948 21532 32004 21534
rect 32060 21420 32116 21476
rect 32508 21420 32564 21476
rect 32620 21532 32676 21588
rect 32844 21756 32900 21812
rect 32844 21532 32900 21588
rect 33852 25116 33908 25172
rect 34076 25004 34132 25060
rect 34524 26514 34580 26516
rect 34524 26462 34526 26514
rect 34526 26462 34578 26514
rect 34578 26462 34580 26514
rect 34524 26460 34580 26462
rect 34860 26402 34916 26404
rect 34860 26350 34862 26402
rect 34862 26350 34914 26402
rect 34914 26350 34916 26402
rect 34860 26348 34916 26350
rect 34972 26236 35028 26292
rect 34412 25228 34468 25284
rect 34860 25506 34916 25508
rect 34860 25454 34862 25506
rect 34862 25454 34914 25506
rect 34914 25454 34916 25506
rect 34860 25452 34916 25454
rect 34972 25340 35028 25396
rect 33852 23436 33908 23492
rect 33292 22652 33348 22708
rect 33516 23324 33572 23380
rect 34076 23436 34132 23492
rect 33404 22370 33460 22372
rect 33404 22318 33406 22370
rect 33406 22318 33458 22370
rect 33458 22318 33460 22370
rect 33404 22316 33460 22318
rect 32172 21084 32228 21140
rect 34300 23154 34356 23156
rect 34300 23102 34302 23154
rect 34302 23102 34354 23154
rect 34354 23102 34356 23154
rect 34300 23100 34356 23102
rect 34636 23324 34692 23380
rect 34860 23266 34916 23268
rect 34860 23214 34862 23266
rect 34862 23214 34914 23266
rect 34914 23214 34916 23266
rect 34860 23212 34916 23214
rect 33516 21756 33572 21812
rect 33964 22204 34020 22260
rect 33740 21868 33796 21924
rect 33628 21532 33684 21588
rect 33852 21810 33908 21812
rect 33852 21758 33854 21810
rect 33854 21758 33906 21810
rect 33906 21758 33908 21810
rect 33852 21756 33908 21758
rect 33180 21196 33236 21252
rect 32732 20802 32788 20804
rect 32732 20750 32734 20802
rect 32734 20750 32786 20802
rect 32786 20750 32788 20802
rect 32732 20748 32788 20750
rect 33516 20802 33572 20804
rect 33516 20750 33518 20802
rect 33518 20750 33570 20802
rect 33570 20750 33572 20802
rect 33516 20748 33572 20750
rect 33852 21084 33908 21140
rect 31052 20636 31108 20692
rect 32172 20690 32228 20692
rect 32172 20638 32174 20690
rect 32174 20638 32226 20690
rect 32226 20638 32228 20690
rect 32172 20636 32228 20638
rect 33852 20636 33908 20692
rect 32508 20578 32564 20580
rect 32508 20526 32510 20578
rect 32510 20526 32562 20578
rect 32562 20526 32564 20578
rect 32508 20524 32564 20526
rect 31388 20188 31444 20244
rect 32508 20076 32564 20132
rect 31948 19964 32004 20020
rect 33180 20018 33236 20020
rect 33180 19966 33182 20018
rect 33182 19966 33234 20018
rect 33234 19966 33236 20018
rect 33180 19964 33236 19966
rect 32284 19794 32340 19796
rect 32284 19742 32286 19794
rect 32286 19742 32338 19794
rect 32338 19742 32340 19794
rect 32284 19740 32340 19742
rect 33068 19794 33124 19796
rect 33068 19742 33070 19794
rect 33070 19742 33122 19794
rect 33122 19742 33124 19794
rect 33068 19740 33124 19742
rect 32732 19628 32788 19684
rect 31948 19516 32004 19572
rect 32844 19516 32900 19572
rect 32732 19458 32788 19460
rect 32732 19406 32734 19458
rect 32734 19406 32786 19458
rect 32786 19406 32788 19458
rect 32732 19404 32788 19406
rect 33068 19404 33124 19460
rect 33068 19234 33124 19236
rect 33068 19182 33070 19234
rect 33070 19182 33122 19234
rect 33122 19182 33124 19234
rect 33068 19180 33124 19182
rect 33180 19068 33236 19124
rect 32284 18620 32340 18676
rect 30604 17164 30660 17220
rect 29484 16882 29540 16884
rect 29484 16830 29486 16882
rect 29486 16830 29538 16882
rect 29538 16830 29540 16882
rect 29484 16828 29540 16830
rect 29372 16380 29428 16436
rect 28812 16156 28868 16212
rect 29372 15314 29428 15316
rect 29372 15262 29374 15314
rect 29374 15262 29426 15314
rect 29426 15262 29428 15314
rect 29372 15260 29428 15262
rect 29932 16770 29988 16772
rect 29932 16718 29934 16770
rect 29934 16718 29986 16770
rect 29986 16718 29988 16770
rect 29932 16716 29988 16718
rect 30492 16994 30548 16996
rect 30492 16942 30494 16994
rect 30494 16942 30546 16994
rect 30546 16942 30548 16994
rect 30492 16940 30548 16942
rect 30828 17276 30884 17332
rect 31276 18172 31332 18228
rect 30716 16828 30772 16884
rect 30044 16268 30100 16324
rect 29708 16098 29764 16100
rect 29708 16046 29710 16098
rect 29710 16046 29762 16098
rect 29762 16046 29764 16098
rect 29708 16044 29764 16046
rect 30380 16098 30436 16100
rect 30380 16046 30382 16098
rect 30382 16046 30434 16098
rect 30434 16046 30436 16098
rect 30380 16044 30436 16046
rect 29820 15874 29876 15876
rect 29820 15822 29822 15874
rect 29822 15822 29874 15874
rect 29874 15822 29876 15874
rect 29820 15820 29876 15822
rect 29825 15706 29881 15708
rect 29825 15654 29827 15706
rect 29827 15654 29879 15706
rect 29879 15654 29881 15706
rect 29825 15652 29881 15654
rect 29929 15706 29985 15708
rect 29929 15654 29931 15706
rect 29931 15654 29983 15706
rect 29983 15654 29985 15706
rect 29929 15652 29985 15654
rect 30033 15706 30089 15708
rect 30033 15654 30035 15706
rect 30035 15654 30087 15706
rect 30087 15654 30089 15706
rect 30033 15652 30089 15654
rect 29596 15372 29652 15428
rect 28588 14812 28644 14868
rect 28476 14364 28532 14420
rect 28252 14252 28308 14308
rect 28252 12178 28308 12180
rect 28252 12126 28254 12178
rect 28254 12126 28306 12178
rect 28306 12126 28308 12178
rect 28252 12124 28308 12126
rect 28588 14252 28644 14308
rect 29148 13916 29204 13972
rect 30716 16156 30772 16212
rect 32396 18450 32452 18452
rect 32396 18398 32398 18450
rect 32398 18398 32450 18450
rect 32450 18398 32452 18450
rect 32396 18396 32452 18398
rect 33068 18450 33124 18452
rect 33068 18398 33070 18450
rect 33070 18398 33122 18450
rect 33122 18398 33124 18450
rect 33068 18396 33124 18398
rect 34188 18732 34244 18788
rect 33292 18674 33348 18676
rect 33292 18622 33294 18674
rect 33294 18622 33346 18674
rect 33346 18622 33348 18674
rect 33292 18620 33348 18622
rect 32732 17666 32788 17668
rect 32732 17614 32734 17666
rect 32734 17614 32786 17666
rect 32786 17614 32788 17666
rect 32732 17612 32788 17614
rect 31052 17442 31108 17444
rect 31052 17390 31054 17442
rect 31054 17390 31106 17442
rect 31106 17390 31108 17442
rect 31052 17388 31108 17390
rect 31388 17276 31444 17332
rect 31724 17276 31780 17332
rect 32172 17164 32228 17220
rect 31724 16994 31780 16996
rect 31724 16942 31726 16994
rect 31726 16942 31778 16994
rect 31778 16942 31780 16994
rect 31724 16940 31780 16942
rect 32396 16882 32452 16884
rect 32396 16830 32398 16882
rect 32398 16830 32450 16882
rect 32450 16830 32452 16882
rect 32396 16828 32452 16830
rect 31500 16268 31556 16324
rect 32284 16716 32340 16772
rect 30716 15372 30772 15428
rect 31724 15986 31780 15988
rect 31724 15934 31726 15986
rect 31726 15934 31778 15986
rect 31778 15934 31780 15986
rect 31724 15932 31780 15934
rect 32060 15986 32116 15988
rect 32060 15934 32062 15986
rect 32062 15934 32114 15986
rect 32114 15934 32116 15986
rect 32060 15932 32116 15934
rect 30828 15820 30884 15876
rect 31948 15874 32004 15876
rect 31948 15822 31950 15874
rect 31950 15822 32002 15874
rect 32002 15822 32004 15874
rect 31948 15820 32004 15822
rect 32284 15596 32340 15652
rect 31276 15372 31332 15428
rect 30492 14476 30548 14532
rect 29372 13804 29428 13860
rect 29932 14306 29988 14308
rect 29932 14254 29934 14306
rect 29934 14254 29986 14306
rect 29986 14254 29988 14306
rect 29932 14252 29988 14254
rect 29825 14138 29881 14140
rect 29825 14086 29827 14138
rect 29827 14086 29879 14138
rect 29879 14086 29881 14138
rect 29825 14084 29881 14086
rect 29929 14138 29985 14140
rect 29929 14086 29931 14138
rect 29931 14086 29983 14138
rect 29983 14086 29985 14138
rect 29929 14084 29985 14086
rect 30033 14138 30089 14140
rect 30033 14086 30035 14138
rect 30035 14086 30087 14138
rect 30087 14086 30089 14138
rect 30033 14084 30089 14086
rect 30268 13916 30324 13972
rect 30716 13970 30772 13972
rect 30716 13918 30718 13970
rect 30718 13918 30770 13970
rect 30770 13918 30772 13970
rect 30716 13916 30772 13918
rect 30156 13804 30212 13860
rect 30940 13858 30996 13860
rect 30940 13806 30942 13858
rect 30942 13806 30994 13858
rect 30994 13806 30996 13858
rect 30940 13804 30996 13806
rect 30380 13356 30436 13412
rect 30156 13132 30212 13188
rect 29596 12738 29652 12740
rect 29596 12686 29598 12738
rect 29598 12686 29650 12738
rect 29650 12686 29652 12738
rect 29596 12684 29652 12686
rect 29372 12572 29428 12628
rect 28924 12402 28980 12404
rect 28924 12350 28926 12402
rect 28926 12350 28978 12402
rect 28978 12350 28980 12402
rect 28924 12348 28980 12350
rect 28364 12012 28420 12068
rect 28588 11564 28644 11620
rect 28140 11340 28196 11396
rect 28476 11228 28532 11284
rect 28140 10556 28196 10612
rect 28364 11170 28420 11172
rect 28364 11118 28366 11170
rect 28366 11118 28418 11170
rect 28418 11118 28420 11170
rect 28364 11116 28420 11118
rect 29825 12570 29881 12572
rect 29825 12518 29827 12570
rect 29827 12518 29879 12570
rect 29879 12518 29881 12570
rect 29825 12516 29881 12518
rect 29929 12570 29985 12572
rect 29929 12518 29931 12570
rect 29931 12518 29983 12570
rect 29983 12518 29985 12570
rect 29929 12516 29985 12518
rect 30033 12570 30089 12572
rect 30033 12518 30035 12570
rect 30035 12518 30087 12570
rect 30087 12518 30089 12570
rect 30033 12516 30089 12518
rect 29484 12124 29540 12180
rect 29820 11564 29876 11620
rect 29596 11452 29652 11508
rect 30940 13580 30996 13636
rect 31612 14252 31668 14308
rect 31500 13522 31556 13524
rect 31500 13470 31502 13522
rect 31502 13470 31554 13522
rect 31554 13470 31556 13522
rect 31500 13468 31556 13470
rect 31388 13132 31444 13188
rect 31164 12962 31220 12964
rect 31164 12910 31166 12962
rect 31166 12910 31218 12962
rect 31218 12910 31220 12962
rect 31164 12908 31220 12910
rect 30940 12850 30996 12852
rect 30940 12798 30942 12850
rect 30942 12798 30994 12850
rect 30994 12798 30996 12850
rect 30940 12796 30996 12798
rect 30604 12684 30660 12740
rect 30380 11452 30436 11508
rect 29708 11282 29764 11284
rect 29708 11230 29710 11282
rect 29710 11230 29762 11282
rect 29762 11230 29764 11282
rect 29708 11228 29764 11230
rect 29484 11116 29540 11172
rect 29372 10780 29428 10836
rect 28476 10220 28532 10276
rect 28364 10108 28420 10164
rect 28028 9212 28084 9268
rect 27804 9154 27860 9156
rect 27804 9102 27806 9154
rect 27806 9102 27858 9154
rect 27858 9102 27860 9154
rect 27804 9100 27860 9102
rect 27580 8876 27636 8932
rect 27244 8204 27300 8260
rect 27020 7644 27076 7700
rect 26684 6972 26740 7028
rect 26684 6300 26740 6356
rect 26348 5292 26404 5348
rect 26572 4956 26628 5012
rect 26572 4172 26628 4228
rect 29825 11002 29881 11004
rect 29825 10950 29827 11002
rect 29827 10950 29879 11002
rect 29879 10950 29881 11002
rect 29825 10948 29881 10950
rect 29929 11002 29985 11004
rect 29929 10950 29931 11002
rect 29931 10950 29983 11002
rect 29983 10950 29985 11002
rect 29929 10948 29985 10950
rect 30033 11002 30089 11004
rect 30033 10950 30035 11002
rect 30035 10950 30087 11002
rect 30087 10950 30089 11002
rect 30380 11004 30436 11060
rect 30033 10948 30089 10950
rect 29708 10610 29764 10612
rect 29708 10558 29710 10610
rect 29710 10558 29762 10610
rect 29762 10558 29764 10610
rect 29708 10556 29764 10558
rect 29820 10220 29876 10276
rect 28812 9212 28868 9268
rect 29372 9548 29428 9604
rect 29825 9434 29881 9436
rect 29825 9382 29827 9434
rect 29827 9382 29879 9434
rect 29879 9382 29881 9434
rect 29825 9380 29881 9382
rect 29929 9434 29985 9436
rect 29929 9382 29931 9434
rect 29931 9382 29983 9434
rect 29983 9382 29985 9434
rect 29929 9380 29985 9382
rect 30033 9434 30089 9436
rect 30033 9382 30035 9434
rect 30035 9382 30087 9434
rect 30087 9382 30089 9434
rect 30033 9380 30089 9382
rect 30044 9212 30100 9268
rect 27804 8652 27860 8708
rect 27692 8540 27748 8596
rect 27804 8428 27860 8484
rect 27692 7868 27748 7924
rect 27356 6636 27412 6692
rect 27580 6412 27636 6468
rect 27468 5906 27524 5908
rect 27468 5854 27470 5906
rect 27470 5854 27522 5906
rect 27522 5854 27524 5906
rect 27468 5852 27524 5854
rect 27468 5516 27524 5572
rect 27132 4450 27188 4452
rect 27132 4398 27134 4450
rect 27134 4398 27186 4450
rect 27186 4398 27188 4450
rect 27132 4396 27188 4398
rect 27580 4226 27636 4228
rect 27580 4174 27582 4226
rect 27582 4174 27634 4226
rect 27634 4174 27636 4226
rect 27580 4172 27636 4174
rect 28140 8428 28196 8484
rect 28252 8652 28308 8708
rect 28028 7644 28084 7700
rect 28476 8540 28532 8596
rect 29932 9100 29988 9156
rect 29036 8930 29092 8932
rect 29036 8878 29038 8930
rect 29038 8878 29090 8930
rect 29090 8878 29092 8930
rect 29036 8876 29092 8878
rect 29596 8204 29652 8260
rect 28700 7644 28756 7700
rect 28700 6076 28756 6132
rect 27804 6018 27860 6020
rect 27804 5966 27806 6018
rect 27806 5966 27858 6018
rect 27858 5966 27860 6018
rect 27804 5964 27860 5966
rect 30268 8540 30324 8596
rect 30492 8988 30548 9044
rect 30716 12124 30772 12180
rect 31388 12178 31444 12180
rect 31388 12126 31390 12178
rect 31390 12126 31442 12178
rect 31442 12126 31444 12178
rect 31388 12124 31444 12126
rect 30940 11452 30996 11508
rect 31500 11564 31556 11620
rect 31164 11394 31220 11396
rect 31164 11342 31166 11394
rect 31166 11342 31218 11394
rect 31218 11342 31220 11394
rect 31164 11340 31220 11342
rect 30716 11282 30772 11284
rect 30716 11230 30718 11282
rect 30718 11230 30770 11282
rect 30770 11230 30772 11282
rect 30716 11228 30772 11230
rect 30940 11170 30996 11172
rect 30940 11118 30942 11170
rect 30942 11118 30994 11170
rect 30994 11118 30996 11170
rect 30940 11116 30996 11118
rect 31276 10780 31332 10836
rect 31724 13356 31780 13412
rect 32284 15314 32340 15316
rect 32284 15262 32286 15314
rect 32286 15262 32338 15314
rect 32338 15262 32340 15314
rect 32284 15260 32340 15262
rect 32508 15874 32564 15876
rect 32508 15822 32510 15874
rect 32510 15822 32562 15874
rect 32562 15822 32564 15874
rect 32508 15820 32564 15822
rect 32620 15596 32676 15652
rect 33740 18060 33796 18116
rect 33740 17724 33796 17780
rect 33068 17388 33124 17444
rect 33180 17052 33236 17108
rect 33852 17948 33908 18004
rect 34748 22540 34804 22596
rect 34524 22316 34580 22372
rect 34412 21868 34468 21924
rect 36204 34018 36260 34020
rect 36204 33966 36206 34018
rect 36206 33966 36258 34018
rect 36258 33966 36260 34018
rect 36204 33964 36260 33966
rect 35532 33852 35588 33908
rect 35420 33404 35476 33460
rect 36540 34636 36596 34692
rect 36764 34354 36820 34356
rect 36764 34302 36766 34354
rect 36766 34302 36818 34354
rect 36818 34302 36820 34354
rect 36764 34300 36820 34302
rect 36876 33964 36932 34020
rect 37324 33964 37380 34020
rect 36428 33628 36484 33684
rect 36979 33738 37035 33740
rect 36979 33686 36981 33738
rect 36981 33686 37033 33738
rect 37033 33686 37035 33738
rect 36979 33684 37035 33686
rect 37083 33738 37139 33740
rect 37083 33686 37085 33738
rect 37085 33686 37137 33738
rect 37137 33686 37139 33738
rect 37083 33684 37139 33686
rect 37187 33738 37243 33740
rect 37187 33686 37189 33738
rect 37189 33686 37241 33738
rect 37241 33686 37243 33738
rect 37187 33684 37243 33686
rect 35532 33346 35588 33348
rect 35532 33294 35534 33346
rect 35534 33294 35586 33346
rect 35586 33294 35588 33346
rect 35532 33292 35588 33294
rect 36428 33292 36484 33348
rect 35420 33234 35476 33236
rect 35420 33182 35422 33234
rect 35422 33182 35474 33234
rect 35474 33182 35476 33234
rect 35420 33180 35476 33182
rect 37100 33346 37156 33348
rect 37100 33294 37102 33346
rect 37102 33294 37154 33346
rect 37154 33294 37156 33346
rect 37100 33292 37156 33294
rect 37436 33292 37492 33348
rect 36316 32674 36372 32676
rect 36316 32622 36318 32674
rect 36318 32622 36370 32674
rect 36370 32622 36372 32674
rect 36316 32620 36372 32622
rect 36988 32956 37044 33012
rect 35532 31778 35588 31780
rect 35532 31726 35534 31778
rect 35534 31726 35586 31778
rect 35586 31726 35588 31778
rect 35532 31724 35588 31726
rect 35980 31612 36036 31668
rect 36428 31890 36484 31892
rect 36428 31838 36430 31890
rect 36430 31838 36482 31890
rect 36482 31838 36484 31890
rect 36428 31836 36484 31838
rect 36316 31106 36372 31108
rect 36316 31054 36318 31106
rect 36318 31054 36370 31106
rect 36370 31054 36372 31106
rect 36316 31052 36372 31054
rect 35196 30716 35252 30772
rect 35980 30268 36036 30324
rect 35532 30044 35588 30100
rect 35420 29372 35476 29428
rect 36204 29596 36260 29652
rect 35308 29260 35364 29316
rect 35420 28140 35476 28196
rect 35868 28700 35924 28756
rect 35756 28418 35812 28420
rect 35756 28366 35758 28418
rect 35758 28366 35810 28418
rect 35810 28366 35812 28418
rect 35756 28364 35812 28366
rect 35756 27916 35812 27972
rect 35644 27858 35700 27860
rect 35644 27806 35646 27858
rect 35646 27806 35698 27858
rect 35698 27806 35700 27858
rect 35644 27804 35700 27806
rect 35756 26908 35812 26964
rect 35308 26402 35364 26404
rect 35308 26350 35310 26402
rect 35310 26350 35362 26402
rect 35362 26350 35364 26402
rect 35308 26348 35364 26350
rect 36540 31612 36596 31668
rect 41020 36876 41076 36932
rect 42252 36876 42308 36932
rect 41916 36764 41972 36820
rect 40796 36652 40852 36708
rect 41356 36652 41412 36708
rect 43036 36876 43092 36932
rect 39228 35420 39284 35476
rect 38780 35196 38836 35252
rect 37884 34802 37940 34804
rect 37884 34750 37886 34802
rect 37886 34750 37938 34802
rect 37938 34750 37940 34802
rect 37884 34748 37940 34750
rect 38780 34748 38836 34804
rect 39788 35532 39844 35588
rect 40908 35810 40964 35812
rect 40908 35758 40910 35810
rect 40910 35758 40962 35810
rect 40962 35758 40964 35810
rect 40908 35756 40964 35758
rect 40236 35474 40292 35476
rect 40236 35422 40238 35474
rect 40238 35422 40290 35474
rect 40290 35422 40292 35474
rect 40236 35420 40292 35422
rect 41020 35420 41076 35476
rect 39564 34802 39620 34804
rect 39564 34750 39566 34802
rect 39566 34750 39618 34802
rect 39618 34750 39620 34802
rect 39564 34748 39620 34750
rect 41132 35196 41188 35252
rect 42140 35420 42196 35476
rect 38444 34524 38500 34580
rect 39004 34636 39060 34692
rect 37996 33740 38052 33796
rect 40012 34242 40068 34244
rect 40012 34190 40014 34242
rect 40014 34190 40066 34242
rect 40066 34190 40068 34242
rect 40012 34188 40068 34190
rect 41580 34188 41636 34244
rect 38220 33292 38276 33348
rect 39564 34130 39620 34132
rect 39564 34078 39566 34130
rect 39566 34078 39618 34130
rect 39618 34078 39620 34130
rect 39564 34076 39620 34078
rect 40124 34130 40180 34132
rect 40124 34078 40126 34130
rect 40126 34078 40178 34130
rect 40178 34078 40180 34130
rect 40124 34076 40180 34078
rect 41020 34130 41076 34132
rect 41020 34078 41022 34130
rect 41022 34078 41074 34130
rect 41074 34078 41076 34130
rect 41020 34076 41076 34078
rect 40908 34018 40964 34020
rect 40908 33966 40910 34018
rect 40910 33966 40962 34018
rect 40962 33966 40964 34018
rect 40908 33964 40964 33966
rect 40012 33906 40068 33908
rect 40012 33854 40014 33906
rect 40014 33854 40066 33906
rect 40066 33854 40068 33906
rect 40012 33852 40068 33854
rect 37548 33180 37604 33236
rect 38780 32844 38836 32900
rect 39452 33346 39508 33348
rect 39452 33294 39454 33346
rect 39454 33294 39506 33346
rect 39506 33294 39508 33346
rect 39452 33292 39508 33294
rect 40236 33292 40292 33348
rect 38668 32674 38724 32676
rect 38668 32622 38670 32674
rect 38670 32622 38722 32674
rect 38722 32622 38724 32674
rect 38668 32620 38724 32622
rect 36979 32170 37035 32172
rect 36979 32118 36981 32170
rect 36981 32118 37033 32170
rect 37033 32118 37035 32170
rect 36979 32116 37035 32118
rect 37083 32170 37139 32172
rect 37083 32118 37085 32170
rect 37085 32118 37137 32170
rect 37137 32118 37139 32170
rect 37083 32116 37139 32118
rect 37187 32170 37243 32172
rect 37187 32118 37189 32170
rect 37189 32118 37241 32170
rect 37241 32118 37243 32170
rect 37187 32116 37243 32118
rect 38444 32562 38500 32564
rect 38444 32510 38446 32562
rect 38446 32510 38498 32562
rect 38498 32510 38500 32562
rect 38444 32508 38500 32510
rect 37772 32450 37828 32452
rect 37772 32398 37774 32450
rect 37774 32398 37826 32450
rect 37826 32398 37828 32450
rect 37772 32396 37828 32398
rect 38668 32396 38724 32452
rect 37884 32060 37940 32116
rect 37772 31890 37828 31892
rect 37772 31838 37774 31890
rect 37774 31838 37826 31890
rect 37826 31838 37828 31890
rect 37772 31836 37828 31838
rect 36652 31500 36708 31556
rect 38108 31500 38164 31556
rect 37548 31164 37604 31220
rect 37324 31052 37380 31108
rect 36979 30602 37035 30604
rect 36979 30550 36981 30602
rect 36981 30550 37033 30602
rect 37033 30550 37035 30602
rect 36979 30548 37035 30550
rect 37083 30602 37139 30604
rect 37083 30550 37085 30602
rect 37085 30550 37137 30602
rect 37137 30550 37139 30602
rect 37083 30548 37139 30550
rect 37187 30602 37243 30604
rect 37187 30550 37189 30602
rect 37189 30550 37241 30602
rect 37241 30550 37243 30602
rect 37187 30548 37243 30550
rect 36988 30098 37044 30100
rect 36988 30046 36990 30098
rect 36990 30046 37042 30098
rect 37042 30046 37044 30098
rect 36988 30044 37044 30046
rect 37100 29932 37156 29988
rect 36428 28924 36484 28980
rect 36540 29426 36596 29428
rect 36540 29374 36542 29426
rect 36542 29374 36594 29426
rect 36594 29374 36596 29426
rect 36540 29372 36596 29374
rect 37660 30044 37716 30100
rect 37772 29596 37828 29652
rect 37324 29314 37380 29316
rect 37324 29262 37326 29314
rect 37326 29262 37378 29314
rect 37378 29262 37380 29314
rect 37324 29260 37380 29262
rect 36979 29034 37035 29036
rect 36979 28982 36981 29034
rect 36981 28982 37033 29034
rect 37033 28982 37035 29034
rect 36979 28980 37035 28982
rect 37083 29034 37139 29036
rect 37083 28982 37085 29034
rect 37085 28982 37137 29034
rect 37137 28982 37139 29034
rect 37083 28980 37139 28982
rect 37187 29034 37243 29036
rect 37187 28982 37189 29034
rect 37189 28982 37241 29034
rect 37241 28982 37243 29034
rect 37187 28980 37243 28982
rect 37100 28812 37156 28868
rect 36204 28418 36260 28420
rect 36204 28366 36206 28418
rect 36206 28366 36258 28418
rect 36258 28366 36260 28418
rect 36204 28364 36260 28366
rect 37212 28364 37268 28420
rect 36316 28028 36372 28084
rect 36204 26514 36260 26516
rect 36204 26462 36206 26514
rect 36206 26462 36258 26514
rect 36258 26462 36260 26514
rect 36204 26460 36260 26462
rect 37212 27916 37268 27972
rect 37660 28812 37716 28868
rect 36979 27466 37035 27468
rect 36979 27414 36981 27466
rect 36981 27414 37033 27466
rect 37033 27414 37035 27466
rect 36979 27412 37035 27414
rect 37083 27466 37139 27468
rect 37083 27414 37085 27466
rect 37085 27414 37137 27466
rect 37137 27414 37139 27466
rect 37083 27412 37139 27414
rect 37187 27466 37243 27468
rect 37187 27414 37189 27466
rect 37189 27414 37241 27466
rect 37241 27414 37243 27466
rect 37187 27412 37243 27414
rect 37324 26460 37380 26516
rect 36092 25676 36148 25732
rect 35308 23884 35364 23940
rect 35196 22764 35252 22820
rect 35308 22876 35364 22932
rect 35308 22428 35364 22484
rect 35308 22146 35364 22148
rect 35308 22094 35310 22146
rect 35310 22094 35362 22146
rect 35362 22094 35364 22146
rect 35308 22092 35364 22094
rect 35868 25452 35924 25508
rect 35644 25116 35700 25172
rect 35980 25228 36036 25284
rect 36204 24610 36260 24612
rect 36204 24558 36206 24610
rect 36206 24558 36258 24610
rect 36258 24558 36260 24610
rect 36204 24556 36260 24558
rect 36979 25898 37035 25900
rect 36979 25846 36981 25898
rect 36981 25846 37033 25898
rect 37033 25846 37035 25898
rect 36979 25844 37035 25846
rect 37083 25898 37139 25900
rect 37083 25846 37085 25898
rect 37085 25846 37137 25898
rect 37137 25846 37139 25898
rect 37083 25844 37139 25846
rect 37187 25898 37243 25900
rect 37187 25846 37189 25898
rect 37189 25846 37241 25898
rect 37241 25846 37243 25898
rect 37187 25844 37243 25846
rect 36988 25730 37044 25732
rect 36988 25678 36990 25730
rect 36990 25678 37042 25730
rect 37042 25678 37044 25730
rect 36988 25676 37044 25678
rect 37324 25676 37380 25732
rect 37324 25394 37380 25396
rect 37324 25342 37326 25394
rect 37326 25342 37378 25394
rect 37378 25342 37380 25394
rect 37324 25340 37380 25342
rect 37100 25282 37156 25284
rect 37100 25230 37102 25282
rect 37102 25230 37154 25282
rect 37154 25230 37156 25282
rect 37100 25228 37156 25230
rect 36428 25116 36484 25172
rect 36764 24892 36820 24948
rect 37100 24722 37156 24724
rect 37100 24670 37102 24722
rect 37102 24670 37154 24722
rect 37154 24670 37156 24722
rect 37100 24668 37156 24670
rect 35644 24108 35700 24164
rect 36092 23996 36148 24052
rect 35868 23772 35924 23828
rect 35868 23436 35924 23492
rect 36979 24330 37035 24332
rect 36979 24278 36981 24330
rect 36981 24278 37033 24330
rect 37033 24278 37035 24330
rect 36979 24276 37035 24278
rect 37083 24330 37139 24332
rect 37083 24278 37085 24330
rect 37085 24278 37137 24330
rect 37137 24278 37139 24330
rect 37083 24276 37139 24278
rect 37187 24330 37243 24332
rect 37187 24278 37189 24330
rect 37189 24278 37241 24330
rect 37241 24278 37243 24330
rect 37187 24276 37243 24278
rect 37100 23772 37156 23828
rect 37548 25282 37604 25284
rect 37548 25230 37550 25282
rect 37550 25230 37602 25282
rect 37602 25230 37604 25282
rect 37548 25228 37604 25230
rect 37548 24892 37604 24948
rect 37548 24050 37604 24052
rect 37548 23998 37550 24050
rect 37550 23998 37602 24050
rect 37602 23998 37604 24050
rect 37548 23996 37604 23998
rect 36428 22988 36484 23044
rect 35644 22482 35700 22484
rect 35644 22430 35646 22482
rect 35646 22430 35698 22482
rect 35698 22430 35700 22482
rect 35644 22428 35700 22430
rect 36204 22428 36260 22484
rect 36316 22204 36372 22260
rect 35756 22092 35812 22148
rect 34524 21644 34580 21700
rect 34636 20972 34692 21028
rect 34972 20914 35028 20916
rect 34972 20862 34974 20914
rect 34974 20862 35026 20914
rect 35026 20862 35028 20914
rect 34972 20860 35028 20862
rect 34636 20188 34692 20244
rect 35420 21698 35476 21700
rect 35420 21646 35422 21698
rect 35422 21646 35474 21698
rect 35474 21646 35476 21698
rect 35420 21644 35476 21646
rect 35420 21308 35476 21364
rect 35420 20690 35476 20692
rect 35420 20638 35422 20690
rect 35422 20638 35474 20690
rect 35474 20638 35476 20690
rect 35420 20636 35476 20638
rect 34412 19458 34468 19460
rect 34412 19406 34414 19458
rect 34414 19406 34466 19458
rect 34466 19406 34468 19458
rect 34412 19404 34468 19406
rect 35196 20076 35252 20132
rect 34524 19180 34580 19236
rect 34300 17836 34356 17892
rect 35308 20018 35364 20020
rect 35308 19966 35310 20018
rect 35310 19966 35362 20018
rect 35362 19966 35364 20018
rect 35308 19964 35364 19966
rect 34636 19628 34692 19684
rect 35308 19292 35364 19348
rect 34748 19180 34804 19236
rect 35308 18620 35364 18676
rect 35644 21196 35700 21252
rect 34636 18450 34692 18452
rect 34636 18398 34638 18450
rect 34638 18398 34690 18450
rect 34690 18398 34692 18450
rect 34636 18396 34692 18398
rect 34860 18060 34916 18116
rect 35532 18844 35588 18900
rect 36092 21196 36148 21252
rect 37548 23660 37604 23716
rect 37212 22876 37268 22932
rect 36979 22762 37035 22764
rect 36979 22710 36981 22762
rect 36981 22710 37033 22762
rect 37033 22710 37035 22762
rect 36979 22708 37035 22710
rect 37083 22762 37139 22764
rect 37083 22710 37085 22762
rect 37085 22710 37137 22762
rect 37137 22710 37139 22762
rect 37083 22708 37139 22710
rect 37187 22762 37243 22764
rect 37187 22710 37189 22762
rect 37189 22710 37241 22762
rect 37241 22710 37243 22762
rect 37187 22708 37243 22710
rect 37324 22764 37380 22820
rect 36764 22428 36820 22484
rect 36988 22540 37044 22596
rect 36428 21980 36484 22036
rect 38780 32060 38836 32116
rect 39116 32732 39172 32788
rect 40012 32844 40068 32900
rect 39116 32562 39172 32564
rect 39116 32510 39118 32562
rect 39118 32510 39170 32562
rect 39170 32510 39172 32562
rect 39116 32508 39172 32510
rect 39340 32060 39396 32116
rect 39452 31836 39508 31892
rect 38780 31724 38836 31780
rect 39676 31778 39732 31780
rect 39676 31726 39678 31778
rect 39678 31726 39730 31778
rect 39730 31726 39732 31778
rect 39676 31724 39732 31726
rect 38892 31666 38948 31668
rect 38892 31614 38894 31666
rect 38894 31614 38946 31666
rect 38946 31614 38948 31666
rect 38892 31612 38948 31614
rect 39228 31164 39284 31220
rect 40348 32562 40404 32564
rect 40348 32510 40350 32562
rect 40350 32510 40402 32562
rect 40402 32510 40404 32562
rect 40348 32508 40404 32510
rect 40796 33122 40852 33124
rect 40796 33070 40798 33122
rect 40798 33070 40850 33122
rect 40850 33070 40852 33122
rect 40796 33068 40852 33070
rect 40124 31164 40180 31220
rect 40572 31778 40628 31780
rect 40572 31726 40574 31778
rect 40574 31726 40626 31778
rect 40626 31726 40628 31778
rect 40572 31724 40628 31726
rect 41244 33292 41300 33348
rect 41468 32562 41524 32564
rect 41468 32510 41470 32562
rect 41470 32510 41522 32562
rect 41522 32510 41524 32562
rect 41468 32508 41524 32510
rect 41132 32396 41188 32452
rect 41244 32338 41300 32340
rect 41244 32286 41246 32338
rect 41246 32286 41298 32338
rect 41298 32286 41300 32338
rect 41244 32284 41300 32286
rect 41692 33068 41748 33124
rect 41916 32674 41972 32676
rect 41916 32622 41918 32674
rect 41918 32622 41970 32674
rect 41970 32622 41972 32674
rect 41916 32620 41972 32622
rect 41804 32396 41860 32452
rect 42028 32284 42084 32340
rect 42028 32060 42084 32116
rect 41804 31836 41860 31892
rect 41804 31612 41860 31668
rect 40908 31218 40964 31220
rect 40908 31166 40910 31218
rect 40910 31166 40962 31218
rect 40962 31166 40964 31218
rect 40908 31164 40964 31166
rect 40348 30828 40404 30884
rect 39340 30604 39396 30660
rect 38780 29596 38836 29652
rect 38220 28418 38276 28420
rect 38220 28366 38222 28418
rect 38222 28366 38274 28418
rect 38274 28366 38276 28418
rect 38220 28364 38276 28366
rect 38220 27858 38276 27860
rect 38220 27806 38222 27858
rect 38222 27806 38274 27858
rect 38274 27806 38276 27858
rect 38220 27804 38276 27806
rect 38668 28418 38724 28420
rect 38668 28366 38670 28418
rect 38670 28366 38722 28418
rect 38722 28366 38724 28418
rect 38668 28364 38724 28366
rect 40012 30210 40068 30212
rect 40012 30158 40014 30210
rect 40014 30158 40066 30210
rect 40066 30158 40068 30210
rect 40012 30156 40068 30158
rect 39340 28588 39396 28644
rect 39564 28642 39620 28644
rect 39564 28590 39566 28642
rect 39566 28590 39618 28642
rect 39618 28590 39620 28642
rect 39564 28588 39620 28590
rect 39900 28700 39956 28756
rect 38780 28028 38836 28084
rect 38332 27020 38388 27076
rect 37996 25900 38052 25956
rect 37884 25788 37940 25844
rect 37772 25452 37828 25508
rect 38332 26236 38388 26292
rect 38556 26290 38612 26292
rect 38556 26238 38558 26290
rect 38558 26238 38610 26290
rect 38610 26238 38612 26290
rect 38556 26236 38612 26238
rect 38220 25900 38276 25956
rect 39116 25900 39172 25956
rect 38332 25452 38388 25508
rect 38556 25506 38612 25508
rect 38556 25454 38558 25506
rect 38558 25454 38610 25506
rect 38610 25454 38612 25506
rect 38556 25452 38612 25454
rect 38108 24834 38164 24836
rect 38108 24782 38110 24834
rect 38110 24782 38162 24834
rect 38162 24782 38164 24834
rect 38108 24780 38164 24782
rect 38444 24722 38500 24724
rect 38444 24670 38446 24722
rect 38446 24670 38498 24722
rect 38498 24670 38500 24722
rect 38444 24668 38500 24670
rect 37884 24220 37940 24276
rect 37996 23996 38052 24052
rect 38108 24556 38164 24612
rect 37884 23266 37940 23268
rect 37884 23214 37886 23266
rect 37886 23214 37938 23266
rect 37938 23214 37940 23266
rect 37884 23212 37940 23214
rect 37996 23660 38052 23716
rect 37772 22764 37828 22820
rect 37996 22652 38052 22708
rect 37772 22594 37828 22596
rect 37772 22542 37774 22594
rect 37774 22542 37826 22594
rect 37826 22542 37828 22594
rect 37772 22540 37828 22542
rect 37436 21644 37492 21700
rect 36204 20412 36260 20468
rect 36092 20300 36148 20356
rect 36428 20802 36484 20804
rect 36428 20750 36430 20802
rect 36430 20750 36482 20802
rect 36482 20750 36484 20802
rect 36428 20748 36484 20750
rect 36979 21194 37035 21196
rect 36979 21142 36981 21194
rect 36981 21142 37033 21194
rect 37033 21142 37035 21194
rect 36979 21140 37035 21142
rect 37083 21194 37139 21196
rect 37083 21142 37085 21194
rect 37085 21142 37137 21194
rect 37137 21142 37139 21194
rect 37083 21140 37139 21142
rect 37187 21194 37243 21196
rect 37187 21142 37189 21194
rect 37189 21142 37241 21194
rect 37241 21142 37243 21194
rect 37187 21140 37243 21142
rect 37436 21308 37492 21364
rect 37436 20914 37492 20916
rect 37436 20862 37438 20914
rect 37438 20862 37490 20914
rect 37490 20862 37492 20914
rect 37436 20860 37492 20862
rect 38220 24332 38276 24388
rect 38220 23324 38276 23380
rect 38444 24050 38500 24052
rect 38444 23998 38446 24050
rect 38446 23998 38498 24050
rect 38498 23998 38500 24050
rect 38444 23996 38500 23998
rect 38332 23042 38388 23044
rect 38332 22990 38334 23042
rect 38334 22990 38386 23042
rect 38386 22990 38388 23042
rect 38332 22988 38388 22990
rect 38220 22876 38276 22932
rect 38892 24892 38948 24948
rect 38892 24668 38948 24724
rect 38780 24610 38836 24612
rect 38780 24558 38782 24610
rect 38782 24558 38834 24610
rect 38834 24558 38836 24610
rect 38780 24556 38836 24558
rect 38556 23884 38612 23940
rect 38556 23436 38612 23492
rect 38556 23100 38612 23156
rect 37660 22258 37716 22260
rect 37660 22206 37662 22258
rect 37662 22206 37714 22258
rect 37714 22206 37716 22258
rect 37660 22204 37716 22206
rect 37884 22204 37940 22260
rect 38444 22316 38500 22372
rect 38108 22204 38164 22260
rect 38108 21980 38164 22036
rect 38444 21756 38500 21812
rect 37772 21196 37828 21252
rect 37996 21644 38052 21700
rect 37660 21084 37716 21140
rect 36652 20300 36708 20356
rect 36204 19852 36260 19908
rect 35980 19346 36036 19348
rect 35980 19294 35982 19346
rect 35982 19294 36034 19346
rect 36034 19294 36036 19346
rect 35980 19292 36036 19294
rect 35756 19068 35812 19124
rect 36092 19068 36148 19124
rect 36428 18844 36484 18900
rect 35084 17724 35140 17780
rect 34412 17612 34468 17668
rect 34748 17666 34804 17668
rect 34748 17614 34750 17666
rect 34750 17614 34802 17666
rect 34802 17614 34804 17666
rect 34748 17612 34804 17614
rect 36316 18674 36372 18676
rect 36316 18622 36318 18674
rect 36318 18622 36370 18674
rect 36370 18622 36372 18674
rect 36316 18620 36372 18622
rect 36764 20412 36820 20468
rect 38668 21644 38724 21700
rect 38780 22764 38836 22820
rect 38108 20802 38164 20804
rect 38108 20750 38110 20802
rect 38110 20750 38162 20802
rect 38162 20750 38164 20802
rect 38108 20748 38164 20750
rect 37996 20636 38052 20692
rect 37548 19852 37604 19908
rect 36979 19626 37035 19628
rect 36979 19574 36981 19626
rect 36981 19574 37033 19626
rect 37033 19574 37035 19626
rect 36979 19572 37035 19574
rect 37083 19626 37139 19628
rect 37083 19574 37085 19626
rect 37085 19574 37137 19626
rect 37137 19574 37139 19626
rect 37083 19572 37139 19574
rect 37187 19626 37243 19628
rect 37187 19574 37189 19626
rect 37189 19574 37241 19626
rect 37241 19574 37243 19626
rect 37187 19572 37243 19574
rect 36764 18620 36820 18676
rect 36876 18396 36932 18452
rect 35868 18338 35924 18340
rect 35868 18286 35870 18338
rect 35870 18286 35922 18338
rect 35922 18286 35924 18338
rect 35868 18284 35924 18286
rect 37660 19628 37716 19684
rect 37884 20076 37940 20132
rect 37548 18732 37604 18788
rect 37660 19180 37716 19236
rect 37324 18450 37380 18452
rect 37324 18398 37326 18450
rect 37326 18398 37378 18450
rect 37378 18398 37380 18450
rect 37324 18396 37380 18398
rect 35868 17948 35924 18004
rect 36988 18172 37044 18228
rect 33740 17052 33796 17108
rect 33404 16994 33460 16996
rect 33404 16942 33406 16994
rect 33406 16942 33458 16994
rect 33458 16942 33460 16994
rect 33404 16940 33460 16942
rect 33852 16994 33908 16996
rect 33852 16942 33854 16994
rect 33854 16942 33906 16994
rect 33906 16942 33908 16994
rect 33852 16940 33908 16942
rect 33964 16882 34020 16884
rect 33964 16830 33966 16882
rect 33966 16830 34018 16882
rect 34018 16830 34020 16882
rect 33964 16828 34020 16830
rect 34076 16604 34132 16660
rect 32844 15932 32900 15988
rect 32956 15874 33012 15876
rect 32956 15822 32958 15874
rect 32958 15822 33010 15874
rect 33010 15822 33012 15874
rect 32956 15820 33012 15822
rect 33404 15708 33460 15764
rect 32844 15260 32900 15316
rect 32956 15596 33012 15652
rect 32508 14306 32564 14308
rect 32508 14254 32510 14306
rect 32510 14254 32562 14306
rect 32562 14254 32564 14306
rect 32508 14252 32564 14254
rect 33628 15596 33684 15652
rect 33404 15260 33460 15316
rect 33516 15372 33572 15428
rect 33964 15260 34020 15316
rect 34412 17442 34468 17444
rect 34412 17390 34414 17442
rect 34414 17390 34466 17442
rect 34466 17390 34468 17442
rect 34412 17388 34468 17390
rect 34748 17106 34804 17108
rect 34748 17054 34750 17106
rect 34750 17054 34802 17106
rect 34802 17054 34804 17106
rect 34748 17052 34804 17054
rect 34636 16940 34692 16996
rect 34412 16882 34468 16884
rect 34412 16830 34414 16882
rect 34414 16830 34466 16882
rect 34466 16830 34468 16882
rect 34412 16828 34468 16830
rect 33068 14306 33124 14308
rect 33068 14254 33070 14306
rect 33070 14254 33122 14306
rect 33122 14254 33124 14306
rect 33068 14252 33124 14254
rect 32060 13580 32116 13636
rect 31836 12572 31892 12628
rect 32284 13634 32340 13636
rect 32284 13582 32286 13634
rect 32286 13582 32338 13634
rect 32338 13582 32340 13634
rect 32284 13580 32340 13582
rect 32508 13634 32564 13636
rect 32508 13582 32510 13634
rect 32510 13582 32562 13634
rect 32562 13582 32564 13634
rect 32508 13580 32564 13582
rect 32396 13468 32452 13524
rect 33404 13580 33460 13636
rect 33292 13468 33348 13524
rect 33740 13916 33796 13972
rect 33180 12012 33236 12068
rect 32172 11900 32228 11956
rect 33068 11900 33124 11956
rect 32508 11788 32564 11844
rect 31836 11452 31892 11508
rect 32396 11452 32452 11508
rect 32060 11228 32116 11284
rect 31724 11004 31780 11060
rect 30716 8540 30772 8596
rect 30940 9548 30996 9604
rect 31052 9436 31108 9492
rect 31164 10108 31220 10164
rect 31500 10668 31556 10724
rect 31724 9884 31780 9940
rect 31388 9714 31444 9716
rect 31388 9662 31390 9714
rect 31390 9662 31442 9714
rect 31442 9662 31444 9714
rect 31388 9660 31444 9662
rect 31724 9212 31780 9268
rect 30380 8204 30436 8260
rect 29825 7866 29881 7868
rect 29825 7814 29827 7866
rect 29827 7814 29879 7866
rect 29879 7814 29881 7866
rect 29825 7812 29881 7814
rect 29929 7866 29985 7868
rect 29929 7814 29931 7866
rect 29931 7814 29983 7866
rect 29983 7814 29985 7866
rect 29929 7812 29985 7814
rect 30033 7866 30089 7868
rect 30033 7814 30035 7866
rect 30035 7814 30087 7866
rect 30087 7814 30089 7866
rect 30033 7812 30089 7814
rect 32172 10834 32228 10836
rect 32172 10782 32174 10834
rect 32174 10782 32226 10834
rect 32226 10782 32228 10834
rect 32172 10780 32228 10782
rect 32060 10220 32116 10276
rect 32508 9884 32564 9940
rect 32844 11116 32900 11172
rect 32620 11004 32676 11060
rect 33628 13692 33684 13748
rect 34076 14306 34132 14308
rect 34076 14254 34078 14306
rect 34078 14254 34130 14306
rect 34130 14254 34132 14306
rect 34076 14252 34132 14254
rect 33964 13634 34020 13636
rect 33964 13582 33966 13634
rect 33966 13582 34018 13634
rect 34018 13582 34020 13634
rect 33964 13580 34020 13582
rect 33964 12796 34020 12852
rect 33628 11452 33684 11508
rect 33404 11340 33460 11396
rect 33404 10610 33460 10612
rect 33404 10558 33406 10610
rect 33406 10558 33458 10610
rect 33458 10558 33460 10610
rect 33404 10556 33460 10558
rect 33852 11900 33908 11956
rect 33964 12012 34020 12068
rect 33740 10444 33796 10500
rect 34188 13634 34244 13636
rect 34188 13582 34190 13634
rect 34190 13582 34242 13634
rect 34242 13582 34244 13634
rect 34188 13580 34244 13582
rect 34972 17388 35028 17444
rect 35084 17276 35140 17332
rect 35532 17666 35588 17668
rect 35532 17614 35534 17666
rect 35534 17614 35586 17666
rect 35586 17614 35588 17666
rect 35532 17612 35588 17614
rect 35644 17500 35700 17556
rect 35868 17052 35924 17108
rect 35980 16604 36036 16660
rect 36204 16882 36260 16884
rect 36204 16830 36206 16882
rect 36206 16830 36258 16882
rect 36258 16830 36260 16882
rect 36204 16828 36260 16830
rect 36652 16882 36708 16884
rect 36652 16830 36654 16882
rect 36654 16830 36706 16882
rect 36706 16830 36708 16882
rect 36652 16828 36708 16830
rect 36428 16716 36484 16772
rect 36092 16156 36148 16212
rect 36316 16268 36372 16324
rect 36428 16044 36484 16100
rect 36540 15986 36596 15988
rect 36540 15934 36542 15986
rect 36542 15934 36594 15986
rect 36594 15934 36596 15986
rect 36540 15932 36596 15934
rect 34972 14418 35028 14420
rect 34972 14366 34974 14418
rect 34974 14366 35026 14418
rect 35026 14366 35028 14418
rect 34972 14364 35028 14366
rect 34636 14306 34692 14308
rect 34636 14254 34638 14306
rect 34638 14254 34690 14306
rect 34690 14254 34692 14306
rect 34636 14252 34692 14254
rect 34412 13916 34468 13972
rect 34412 12066 34468 12068
rect 34412 12014 34414 12066
rect 34414 12014 34466 12066
rect 34466 12014 34468 12066
rect 34412 12012 34468 12014
rect 34076 11676 34132 11732
rect 33180 10220 33236 10276
rect 32172 9154 32228 9156
rect 32172 9102 32174 9154
rect 32174 9102 32226 9154
rect 32226 9102 32228 9154
rect 32172 9100 32228 9102
rect 32844 9212 32900 9268
rect 33180 9436 33236 9492
rect 31500 8876 31556 8932
rect 31052 8428 31108 8484
rect 30940 8034 30996 8036
rect 30940 7982 30942 8034
rect 30942 7982 30994 8034
rect 30994 7982 30996 8034
rect 30940 7980 30996 7982
rect 30380 7532 30436 7588
rect 29596 7308 29652 7364
rect 29148 6860 29204 6916
rect 30940 7586 30996 7588
rect 30940 7534 30942 7586
rect 30942 7534 30994 7586
rect 30994 7534 30996 7586
rect 30940 7532 30996 7534
rect 31276 8540 31332 8596
rect 31388 7420 31444 7476
rect 31052 7308 31108 7364
rect 30044 6972 30100 7028
rect 29820 6636 29876 6692
rect 29148 6578 29204 6580
rect 29148 6526 29150 6578
rect 29150 6526 29202 6578
rect 29202 6526 29204 6578
rect 29148 6524 29204 6526
rect 29708 6466 29764 6468
rect 29708 6414 29710 6466
rect 29710 6414 29762 6466
rect 29762 6414 29764 6466
rect 29708 6412 29764 6414
rect 29825 6298 29881 6300
rect 29825 6246 29827 6298
rect 29827 6246 29879 6298
rect 29879 6246 29881 6298
rect 29825 6244 29881 6246
rect 29929 6298 29985 6300
rect 29929 6246 29931 6298
rect 29931 6246 29983 6298
rect 29983 6246 29985 6298
rect 29929 6244 29985 6246
rect 30033 6298 30089 6300
rect 30033 6246 30035 6298
rect 30035 6246 30087 6298
rect 30087 6246 30089 6298
rect 30033 6244 30089 6246
rect 29708 6076 29764 6132
rect 28924 5906 28980 5908
rect 28924 5854 28926 5906
rect 28926 5854 28978 5906
rect 28978 5854 28980 5906
rect 28924 5852 28980 5854
rect 28588 5180 28644 5236
rect 28364 4732 28420 4788
rect 27804 4396 27860 4452
rect 27692 4060 27748 4116
rect 27916 4172 27972 4228
rect 25900 2828 25956 2884
rect 27356 3500 27412 3556
rect 28812 4508 28868 4564
rect 28476 3724 28532 3780
rect 28588 4060 28644 4116
rect 29708 5516 29764 5572
rect 29260 5404 29316 5460
rect 29596 5346 29652 5348
rect 29596 5294 29598 5346
rect 29598 5294 29650 5346
rect 29650 5294 29652 5346
rect 29596 5292 29652 5294
rect 29372 4732 29428 4788
rect 29484 4060 29540 4116
rect 30380 5964 30436 6020
rect 29825 4730 29881 4732
rect 29825 4678 29827 4730
rect 29827 4678 29879 4730
rect 29879 4678 29881 4730
rect 29825 4676 29881 4678
rect 29929 4730 29985 4732
rect 29929 4678 29931 4730
rect 29931 4678 29983 4730
rect 29983 4678 29985 4730
rect 29929 4676 29985 4678
rect 30033 4730 30089 4732
rect 30033 4678 30035 4730
rect 30035 4678 30087 4730
rect 30087 4678 30089 4730
rect 30033 4676 30089 4678
rect 30604 5964 30660 6020
rect 30380 4508 30436 4564
rect 30604 4450 30660 4452
rect 30604 4398 30606 4450
rect 30606 4398 30658 4450
rect 30658 4398 30660 4450
rect 30604 4396 30660 4398
rect 29820 4338 29876 4340
rect 29820 4286 29822 4338
rect 29822 4286 29874 4338
rect 29874 4286 29876 4338
rect 29820 4284 29876 4286
rect 30828 6578 30884 6580
rect 30828 6526 30830 6578
rect 30830 6526 30882 6578
rect 30882 6526 30884 6578
rect 30828 6524 30884 6526
rect 31164 6412 31220 6468
rect 31052 5794 31108 5796
rect 31052 5742 31054 5794
rect 31054 5742 31106 5794
rect 31106 5742 31108 5794
rect 31052 5740 31108 5742
rect 31388 6300 31444 6356
rect 32060 8092 32116 8148
rect 31612 7980 31668 8036
rect 31612 7084 31668 7140
rect 33180 8258 33236 8260
rect 33180 8206 33182 8258
rect 33182 8206 33234 8258
rect 33234 8206 33236 8258
rect 33180 8204 33236 8206
rect 32732 8092 32788 8148
rect 33516 10220 33572 10276
rect 33516 9436 33572 9492
rect 33628 9826 33684 9828
rect 33628 9774 33630 9826
rect 33630 9774 33682 9826
rect 33682 9774 33684 9826
rect 33628 9772 33684 9774
rect 33740 8540 33796 8596
rect 33404 8316 33460 8372
rect 35196 14364 35252 14420
rect 34860 12908 34916 12964
rect 34972 12796 35028 12852
rect 34860 12572 34916 12628
rect 34860 12066 34916 12068
rect 34860 12014 34862 12066
rect 34862 12014 34914 12066
rect 34914 12014 34916 12066
rect 34860 12012 34916 12014
rect 33964 10668 34020 10724
rect 34300 11170 34356 11172
rect 34300 11118 34302 11170
rect 34302 11118 34354 11170
rect 34354 11118 34356 11170
rect 34300 11116 34356 11118
rect 34524 11004 34580 11060
rect 34076 10332 34132 10388
rect 34300 10610 34356 10612
rect 34300 10558 34302 10610
rect 34302 10558 34354 10610
rect 34354 10558 34356 10610
rect 34300 10556 34356 10558
rect 34300 9996 34356 10052
rect 34636 8876 34692 8932
rect 34860 11340 34916 11396
rect 34860 9996 34916 10052
rect 35084 10332 35140 10388
rect 35644 14924 35700 14980
rect 35756 15484 35812 15540
rect 35644 14252 35700 14308
rect 35420 14028 35476 14084
rect 35308 11116 35364 11172
rect 35420 13804 35476 13860
rect 35420 11004 35476 11060
rect 35420 10108 35476 10164
rect 35308 9772 35364 9828
rect 35196 9212 35252 9268
rect 34860 8930 34916 8932
rect 34860 8878 34862 8930
rect 34862 8878 34914 8930
rect 34914 8878 34916 8930
rect 34860 8876 34916 8878
rect 33852 8204 33908 8260
rect 34300 8316 34356 8372
rect 33628 7980 33684 8036
rect 32284 7420 32340 7476
rect 32732 7196 32788 7252
rect 31612 5180 31668 5236
rect 31724 6524 31780 6580
rect 32620 6748 32676 6804
rect 32508 6636 32564 6692
rect 31836 6018 31892 6020
rect 31836 5966 31838 6018
rect 31838 5966 31890 6018
rect 31890 5966 31892 6018
rect 31836 5964 31892 5966
rect 32396 5292 32452 5348
rect 33180 7084 33236 7140
rect 32956 6636 33012 6692
rect 32844 6578 32900 6580
rect 32844 6526 32846 6578
rect 32846 6526 32898 6578
rect 32898 6526 32900 6578
rect 32844 6524 32900 6526
rect 33292 6636 33348 6692
rect 33516 7644 33572 7700
rect 34188 8092 34244 8148
rect 33740 7474 33796 7476
rect 33740 7422 33742 7474
rect 33742 7422 33794 7474
rect 33794 7422 33796 7474
rect 33740 7420 33796 7422
rect 33852 7362 33908 7364
rect 33852 7310 33854 7362
rect 33854 7310 33906 7362
rect 33906 7310 33908 7362
rect 33852 7308 33908 7310
rect 34300 6972 34356 7028
rect 33628 6636 33684 6692
rect 34524 7756 34580 7812
rect 34300 6690 34356 6692
rect 34300 6638 34302 6690
rect 34302 6638 34354 6690
rect 34354 6638 34356 6690
rect 34300 6636 34356 6638
rect 32956 5906 33012 5908
rect 32956 5854 32958 5906
rect 32958 5854 33010 5906
rect 33010 5854 33012 5906
rect 32956 5852 33012 5854
rect 33068 5180 33124 5236
rect 32396 4844 32452 4900
rect 29932 4226 29988 4228
rect 29932 4174 29934 4226
rect 29934 4174 29986 4226
rect 29986 4174 29988 4226
rect 29932 4172 29988 4174
rect 29708 3778 29764 3780
rect 29708 3726 29710 3778
rect 29710 3726 29762 3778
rect 29762 3726 29764 3778
rect 29708 3724 29764 3726
rect 29932 3724 29988 3780
rect 30604 3554 30660 3556
rect 30604 3502 30606 3554
rect 30606 3502 30658 3554
rect 30658 3502 30660 3554
rect 30604 3500 30660 3502
rect 30940 3442 30996 3444
rect 30940 3390 30942 3442
rect 30942 3390 30994 3442
rect 30994 3390 30996 3442
rect 30940 3388 30996 3390
rect 28924 3276 28980 3332
rect 29825 3162 29881 3164
rect 29825 3110 29827 3162
rect 29827 3110 29879 3162
rect 29879 3110 29881 3162
rect 29825 3108 29881 3110
rect 29929 3162 29985 3164
rect 29929 3110 29931 3162
rect 29931 3110 29983 3162
rect 29983 3110 29985 3162
rect 29929 3108 29985 3110
rect 30033 3162 30089 3164
rect 30033 3110 30035 3162
rect 30035 3110 30087 3162
rect 30087 3110 30089 3162
rect 30033 3108 30089 3110
rect 30268 2940 30324 2996
rect 32620 4508 32676 4564
rect 33292 4338 33348 4340
rect 33292 4286 33294 4338
rect 33294 4286 33346 4338
rect 33346 4286 33348 4338
rect 33292 4284 33348 4286
rect 32508 4226 32564 4228
rect 32508 4174 32510 4226
rect 32510 4174 32562 4226
rect 32562 4174 32564 4226
rect 32508 4172 32564 4174
rect 33292 3612 33348 3668
rect 33964 6018 34020 6020
rect 33964 5966 33966 6018
rect 33966 5966 34018 6018
rect 34018 5966 34020 6018
rect 33964 5964 34020 5966
rect 33852 5906 33908 5908
rect 33852 5854 33854 5906
rect 33854 5854 33906 5906
rect 33906 5854 33908 5906
rect 33852 5852 33908 5854
rect 34076 5628 34132 5684
rect 33628 4844 33684 4900
rect 34524 5964 34580 6020
rect 34300 5628 34356 5684
rect 34076 4562 34132 4564
rect 34076 4510 34078 4562
rect 34078 4510 34130 4562
rect 34130 4510 34132 4562
rect 34076 4508 34132 4510
rect 33852 4450 33908 4452
rect 33852 4398 33854 4450
rect 33854 4398 33906 4450
rect 33906 4398 33908 4450
rect 33852 4396 33908 4398
rect 34524 5234 34580 5236
rect 34524 5182 34526 5234
rect 34526 5182 34578 5234
rect 34578 5182 34580 5234
rect 34524 5180 34580 5182
rect 34748 8370 34804 8372
rect 34748 8318 34750 8370
rect 34750 8318 34802 8370
rect 34802 8318 34804 8370
rect 34748 8316 34804 8318
rect 36979 18058 37035 18060
rect 36979 18006 36981 18058
rect 36981 18006 37033 18058
rect 37033 18006 37035 18058
rect 36979 18004 37035 18006
rect 37083 18058 37139 18060
rect 37083 18006 37085 18058
rect 37085 18006 37137 18058
rect 37137 18006 37139 18058
rect 37083 18004 37139 18006
rect 37187 18058 37243 18060
rect 37187 18006 37189 18058
rect 37189 18006 37241 18058
rect 37241 18006 37243 18058
rect 37187 18004 37243 18006
rect 37100 17778 37156 17780
rect 37100 17726 37102 17778
rect 37102 17726 37154 17778
rect 37154 17726 37156 17778
rect 37100 17724 37156 17726
rect 37324 17724 37380 17780
rect 37548 17948 37604 18004
rect 36876 16882 36932 16884
rect 36876 16830 36878 16882
rect 36878 16830 36930 16882
rect 36930 16830 36932 16882
rect 36876 16828 36932 16830
rect 37772 19068 37828 19124
rect 38444 20018 38500 20020
rect 38444 19966 38446 20018
rect 38446 19966 38498 20018
rect 38498 19966 38500 20018
rect 38444 19964 38500 19966
rect 38668 19628 38724 19684
rect 38780 20018 38836 20020
rect 38780 19966 38782 20018
rect 38782 19966 38834 20018
rect 38834 19966 38836 20018
rect 38780 19964 38836 19966
rect 39340 25676 39396 25732
rect 39116 25564 39172 25620
rect 39452 25452 39508 25508
rect 39228 24834 39284 24836
rect 39228 24782 39230 24834
rect 39230 24782 39282 24834
rect 39282 24782 39284 24834
rect 39228 24780 39284 24782
rect 41468 30882 41524 30884
rect 41468 30830 41470 30882
rect 41470 30830 41522 30882
rect 41522 30830 41524 30882
rect 41468 30828 41524 30830
rect 41244 30770 41300 30772
rect 41244 30718 41246 30770
rect 41246 30718 41298 30770
rect 41298 30718 41300 30770
rect 41244 30716 41300 30718
rect 41468 30268 41524 30324
rect 41244 28924 41300 28980
rect 40796 28700 40852 28756
rect 41580 28642 41636 28644
rect 41580 28590 41582 28642
rect 41582 28590 41634 28642
rect 41634 28590 41636 28642
rect 41580 28588 41636 28590
rect 40684 28530 40740 28532
rect 40684 28478 40686 28530
rect 40686 28478 40738 28530
rect 40738 28478 40740 28530
rect 40684 28476 40740 28478
rect 41244 28476 41300 28532
rect 41020 28082 41076 28084
rect 41020 28030 41022 28082
rect 41022 28030 41074 28082
rect 41074 28030 41076 28082
rect 41020 28028 41076 28030
rect 40236 27916 40292 27972
rect 40908 27970 40964 27972
rect 40908 27918 40910 27970
rect 40910 27918 40962 27970
rect 40962 27918 40964 27970
rect 40908 27916 40964 27918
rect 41244 27916 41300 27972
rect 40124 26402 40180 26404
rect 40124 26350 40126 26402
rect 40126 26350 40178 26402
rect 40178 26350 40180 26402
rect 40124 26348 40180 26350
rect 41020 26402 41076 26404
rect 41020 26350 41022 26402
rect 41022 26350 41074 26402
rect 41074 26350 41076 26402
rect 41020 26348 41076 26350
rect 40348 26290 40404 26292
rect 40348 26238 40350 26290
rect 40350 26238 40402 26290
rect 40402 26238 40404 26290
rect 40348 26236 40404 26238
rect 41132 26290 41188 26292
rect 41132 26238 41134 26290
rect 41134 26238 41186 26290
rect 41186 26238 41188 26290
rect 41132 26236 41188 26238
rect 40012 25452 40068 25508
rect 39788 25340 39844 25396
rect 39116 24220 39172 24276
rect 39004 23826 39060 23828
rect 39004 23774 39006 23826
rect 39006 23774 39058 23826
rect 39058 23774 39060 23826
rect 39004 23772 39060 23774
rect 40572 25116 40628 25172
rect 40012 24556 40068 24612
rect 41244 24668 41300 24724
rect 39900 23938 39956 23940
rect 39900 23886 39902 23938
rect 39902 23886 39954 23938
rect 39954 23886 39956 23938
rect 39900 23884 39956 23886
rect 39788 23660 39844 23716
rect 39676 23548 39732 23604
rect 39564 23324 39620 23380
rect 39564 23100 39620 23156
rect 39228 22540 39284 22596
rect 39676 22428 39732 22484
rect 39228 22204 39284 22260
rect 39004 22092 39060 22148
rect 39228 21532 39284 21588
rect 39676 21756 39732 21812
rect 40908 23548 40964 23604
rect 39900 23324 39956 23380
rect 40460 22876 40516 22932
rect 39900 22316 39956 22372
rect 40236 22652 40292 22708
rect 40236 22092 40292 22148
rect 40348 21644 40404 21700
rect 39452 21532 39508 21588
rect 40124 21586 40180 21588
rect 40124 21534 40126 21586
rect 40126 21534 40178 21586
rect 40178 21534 40180 21586
rect 40124 21532 40180 21534
rect 39340 21474 39396 21476
rect 39340 21422 39342 21474
rect 39342 21422 39394 21474
rect 39394 21422 39396 21474
rect 39340 21420 39396 21422
rect 38556 19516 38612 19572
rect 37996 19346 38052 19348
rect 37996 19294 37998 19346
rect 37998 19294 38050 19346
rect 38050 19294 38052 19346
rect 37996 19292 38052 19294
rect 37884 18620 37940 18676
rect 36979 16490 37035 16492
rect 36979 16438 36981 16490
rect 36981 16438 37033 16490
rect 37033 16438 37035 16490
rect 36979 16436 37035 16438
rect 37083 16490 37139 16492
rect 37083 16438 37085 16490
rect 37085 16438 37137 16490
rect 37137 16438 37139 16490
rect 37083 16436 37139 16438
rect 37187 16490 37243 16492
rect 37187 16438 37189 16490
rect 37189 16438 37241 16490
rect 37241 16438 37243 16490
rect 37187 16436 37243 16438
rect 36988 16098 37044 16100
rect 36988 16046 36990 16098
rect 36990 16046 37042 16098
rect 37042 16046 37044 16098
rect 36988 16044 37044 16046
rect 37212 15986 37268 15988
rect 37212 15934 37214 15986
rect 37214 15934 37266 15986
rect 37266 15934 37268 15986
rect 37212 15932 37268 15934
rect 36979 14922 37035 14924
rect 36979 14870 36981 14922
rect 36981 14870 37033 14922
rect 37033 14870 37035 14922
rect 36979 14868 37035 14870
rect 37083 14922 37139 14924
rect 37083 14870 37085 14922
rect 37085 14870 37137 14922
rect 37137 14870 37139 14922
rect 37083 14868 37139 14870
rect 37187 14922 37243 14924
rect 37187 14870 37189 14922
rect 37189 14870 37241 14922
rect 37241 14870 37243 14922
rect 37187 14868 37243 14870
rect 37324 14700 37380 14756
rect 36204 14588 36260 14644
rect 37100 14530 37156 14532
rect 37100 14478 37102 14530
rect 37102 14478 37154 14530
rect 37154 14478 37156 14530
rect 37100 14476 37156 14478
rect 37660 14476 37716 14532
rect 36428 13858 36484 13860
rect 36428 13806 36430 13858
rect 36430 13806 36482 13858
rect 36482 13806 36484 13858
rect 36428 13804 36484 13806
rect 37436 13804 37492 13860
rect 36979 13354 37035 13356
rect 36979 13302 36981 13354
rect 36981 13302 37033 13354
rect 37033 13302 37035 13354
rect 36979 13300 37035 13302
rect 37083 13354 37139 13356
rect 37083 13302 37085 13354
rect 37085 13302 37137 13354
rect 37137 13302 37139 13354
rect 37083 13300 37139 13302
rect 37187 13354 37243 13356
rect 37187 13302 37189 13354
rect 37189 13302 37241 13354
rect 37241 13302 37243 13354
rect 37187 13300 37243 13302
rect 37660 12908 37716 12964
rect 35644 12124 35700 12180
rect 36764 12178 36820 12180
rect 36764 12126 36766 12178
rect 36766 12126 36818 12178
rect 36818 12126 36820 12178
rect 36764 12124 36820 12126
rect 37660 12178 37716 12180
rect 37660 12126 37662 12178
rect 37662 12126 37714 12178
rect 37714 12126 37716 12178
rect 37660 12124 37716 12126
rect 36316 12012 36372 12068
rect 37884 12066 37940 12068
rect 37884 12014 37886 12066
rect 37886 12014 37938 12066
rect 37938 12014 37940 12066
rect 37884 12012 37940 12014
rect 36979 11786 37035 11788
rect 36979 11734 36981 11786
rect 36981 11734 37033 11786
rect 37033 11734 37035 11786
rect 36979 11732 37035 11734
rect 37083 11786 37139 11788
rect 37083 11734 37085 11786
rect 37085 11734 37137 11786
rect 37137 11734 37139 11786
rect 37083 11732 37139 11734
rect 37187 11786 37243 11788
rect 37187 11734 37189 11786
rect 37189 11734 37241 11786
rect 37241 11734 37243 11786
rect 37187 11732 37243 11734
rect 35756 11228 35812 11284
rect 35756 11004 35812 11060
rect 35756 10444 35812 10500
rect 35868 10386 35924 10388
rect 35868 10334 35870 10386
rect 35870 10334 35922 10386
rect 35922 10334 35924 10386
rect 35868 10332 35924 10334
rect 35756 9996 35812 10052
rect 36316 10722 36372 10724
rect 36316 10670 36318 10722
rect 36318 10670 36370 10722
rect 36370 10670 36372 10722
rect 36316 10668 36372 10670
rect 38780 18674 38836 18676
rect 38780 18622 38782 18674
rect 38782 18622 38834 18674
rect 38834 18622 38836 18674
rect 38780 18620 38836 18622
rect 38332 18396 38388 18452
rect 38108 17724 38164 17780
rect 38108 16882 38164 16884
rect 38108 16830 38110 16882
rect 38110 16830 38162 16882
rect 38162 16830 38164 16882
rect 38108 16828 38164 16830
rect 38220 16268 38276 16324
rect 38108 16210 38164 16212
rect 38108 16158 38110 16210
rect 38110 16158 38162 16210
rect 38162 16158 38164 16210
rect 38108 16156 38164 16158
rect 38220 16044 38276 16100
rect 38668 16940 38724 16996
rect 37996 11452 38052 11508
rect 37324 11282 37380 11284
rect 37324 11230 37326 11282
rect 37326 11230 37378 11282
rect 37378 11230 37380 11282
rect 37324 11228 37380 11230
rect 37212 10722 37268 10724
rect 37212 10670 37214 10722
rect 37214 10670 37266 10722
rect 37266 10670 37268 10722
rect 37212 10668 37268 10670
rect 36979 10218 37035 10220
rect 36979 10166 36981 10218
rect 36981 10166 37033 10218
rect 37033 10166 37035 10218
rect 36979 10164 37035 10166
rect 37083 10218 37139 10220
rect 37083 10166 37085 10218
rect 37085 10166 37137 10218
rect 37137 10166 37139 10218
rect 37083 10164 37139 10166
rect 37187 10218 37243 10220
rect 37187 10166 37189 10218
rect 37189 10166 37241 10218
rect 37241 10166 37243 10218
rect 37187 10164 37243 10166
rect 35644 8988 35700 9044
rect 35980 8818 36036 8820
rect 35980 8766 35982 8818
rect 35982 8766 36034 8818
rect 36034 8766 36036 8818
rect 35980 8764 36036 8766
rect 38332 9324 38388 9380
rect 35420 8316 35476 8372
rect 35980 8316 36036 8372
rect 36092 8258 36148 8260
rect 36092 8206 36094 8258
rect 36094 8206 36146 8258
rect 36146 8206 36148 8258
rect 36092 8204 36148 8206
rect 35868 7980 35924 8036
rect 35420 7698 35476 7700
rect 35420 7646 35422 7698
rect 35422 7646 35474 7698
rect 35474 7646 35476 7698
rect 35420 7644 35476 7646
rect 34972 7084 35028 7140
rect 34748 6972 34804 7028
rect 35084 6802 35140 6804
rect 35084 6750 35086 6802
rect 35086 6750 35138 6802
rect 35138 6750 35140 6802
rect 35084 6748 35140 6750
rect 34860 6690 34916 6692
rect 34860 6638 34862 6690
rect 34862 6638 34914 6690
rect 34914 6638 34916 6690
rect 34860 6636 34916 6638
rect 34748 6130 34804 6132
rect 34748 6078 34750 6130
rect 34750 6078 34802 6130
rect 34802 6078 34804 6130
rect 34748 6076 34804 6078
rect 36979 8650 37035 8652
rect 36979 8598 36981 8650
rect 36981 8598 37033 8650
rect 37033 8598 37035 8650
rect 36979 8596 37035 8598
rect 37083 8650 37139 8652
rect 37083 8598 37085 8650
rect 37085 8598 37137 8650
rect 37137 8598 37139 8650
rect 37083 8596 37139 8598
rect 37187 8650 37243 8652
rect 37187 8598 37189 8650
rect 37189 8598 37241 8650
rect 37241 8598 37243 8650
rect 37187 8596 37243 8598
rect 37212 8204 37268 8260
rect 36428 7756 36484 7812
rect 36876 8092 36932 8148
rect 37772 8316 37828 8372
rect 36876 7586 36932 7588
rect 36876 7534 36878 7586
rect 36878 7534 36930 7586
rect 36930 7534 36932 7586
rect 36876 7532 36932 7534
rect 37772 7756 37828 7812
rect 37436 7196 37492 7252
rect 38220 7420 38276 7476
rect 36979 7082 37035 7084
rect 36979 7030 36981 7082
rect 36981 7030 37033 7082
rect 37033 7030 37035 7082
rect 36979 7028 37035 7030
rect 37083 7082 37139 7084
rect 37083 7030 37085 7082
rect 37085 7030 37137 7082
rect 37137 7030 37139 7082
rect 37083 7028 37139 7030
rect 37187 7082 37243 7084
rect 37187 7030 37189 7082
rect 37189 7030 37241 7082
rect 37241 7030 37243 7082
rect 37187 7028 37243 7030
rect 35980 6802 36036 6804
rect 35980 6750 35982 6802
rect 35982 6750 36034 6802
rect 36034 6750 36036 6802
rect 35980 6748 36036 6750
rect 36540 6748 36596 6804
rect 35756 6690 35812 6692
rect 35756 6638 35758 6690
rect 35758 6638 35810 6690
rect 35810 6638 35812 6690
rect 35756 6636 35812 6638
rect 35644 6076 35700 6132
rect 35196 5628 35252 5684
rect 37324 6018 37380 6020
rect 37324 5966 37326 6018
rect 37326 5966 37378 6018
rect 37378 5966 37380 6018
rect 37324 5964 37380 5966
rect 36979 5514 37035 5516
rect 36979 5462 36981 5514
rect 36981 5462 37033 5514
rect 37033 5462 37035 5514
rect 36979 5460 37035 5462
rect 37083 5514 37139 5516
rect 37083 5462 37085 5514
rect 37085 5462 37137 5514
rect 37137 5462 37139 5514
rect 37083 5460 37139 5462
rect 37187 5514 37243 5516
rect 37187 5462 37189 5514
rect 37189 5462 37241 5514
rect 37241 5462 37243 5514
rect 37187 5460 37243 5462
rect 37100 5292 37156 5348
rect 35756 5234 35812 5236
rect 35756 5182 35758 5234
rect 35758 5182 35810 5234
rect 35810 5182 35812 5234
rect 35756 5180 35812 5182
rect 34524 4898 34580 4900
rect 34524 4846 34526 4898
rect 34526 4846 34578 4898
rect 34578 4846 34580 4898
rect 34524 4844 34580 4846
rect 34972 5068 35028 5124
rect 34188 4338 34244 4340
rect 34188 4286 34190 4338
rect 34190 4286 34242 4338
rect 34242 4286 34244 4338
rect 34188 4284 34244 4286
rect 34636 4508 34692 4564
rect 36092 4956 36148 5012
rect 37548 5010 37604 5012
rect 37548 4958 37550 5010
rect 37550 4958 37602 5010
rect 37602 4958 37604 5010
rect 37548 4956 37604 4958
rect 37100 4620 37156 4676
rect 38108 6412 38164 6468
rect 38332 5682 38388 5684
rect 38332 5630 38334 5682
rect 38334 5630 38386 5682
rect 38386 5630 38388 5682
rect 38332 5628 38388 5630
rect 37772 4396 37828 4452
rect 38332 4620 38388 4676
rect 34636 3948 34692 4004
rect 37324 4060 37380 4116
rect 36979 3946 37035 3948
rect 36979 3894 36981 3946
rect 36981 3894 37033 3946
rect 37033 3894 37035 3946
rect 36979 3892 37035 3894
rect 37083 3946 37139 3948
rect 37083 3894 37085 3946
rect 37085 3894 37137 3946
rect 37137 3894 37139 3946
rect 37083 3892 37139 3894
rect 37187 3946 37243 3948
rect 37187 3894 37189 3946
rect 37189 3894 37241 3946
rect 37241 3894 37243 3946
rect 37187 3892 37243 3894
rect 34636 3724 34692 3780
rect 35084 3554 35140 3556
rect 35084 3502 35086 3554
rect 35086 3502 35138 3554
rect 35138 3502 35140 3554
rect 35084 3500 35140 3502
rect 32844 3442 32900 3444
rect 32844 3390 32846 3442
rect 32846 3390 32898 3442
rect 32898 3390 32900 3442
rect 32844 3388 32900 3390
rect 31276 2380 31332 2436
rect 28924 2268 28980 2324
rect 34188 3442 34244 3444
rect 34188 3390 34190 3442
rect 34190 3390 34242 3442
rect 34242 3390 34244 3442
rect 34188 3388 34244 3390
rect 33740 3330 33796 3332
rect 33740 3278 33742 3330
rect 33742 3278 33794 3330
rect 33794 3278 33796 3330
rect 33740 3276 33796 3278
rect 38556 14700 38612 14756
rect 38668 15820 38724 15876
rect 38892 16044 38948 16100
rect 38668 14530 38724 14532
rect 38668 14478 38670 14530
rect 38670 14478 38722 14530
rect 38722 14478 38724 14530
rect 38668 14476 38724 14478
rect 38892 14700 38948 14756
rect 39228 19852 39284 19908
rect 39452 20636 39508 20692
rect 39676 20018 39732 20020
rect 39676 19966 39678 20018
rect 39678 19966 39730 20018
rect 39730 19966 39732 20018
rect 39676 19964 39732 19966
rect 39340 19628 39396 19684
rect 39340 17724 39396 17780
rect 39564 16828 39620 16884
rect 39900 16098 39956 16100
rect 39900 16046 39902 16098
rect 39902 16046 39954 16098
rect 39954 16046 39956 16098
rect 39900 16044 39956 16046
rect 40684 22092 40740 22148
rect 40348 19740 40404 19796
rect 40460 20524 40516 20580
rect 40124 19516 40180 19572
rect 40908 21532 40964 21588
rect 41356 22258 41412 22260
rect 41356 22206 41358 22258
rect 41358 22206 41410 22258
rect 41410 22206 41412 22258
rect 41356 22204 41412 22206
rect 42028 26796 42084 26852
rect 42252 34860 42308 34916
rect 42700 35810 42756 35812
rect 42700 35758 42702 35810
rect 42702 35758 42754 35810
rect 42754 35758 42756 35810
rect 42700 35756 42756 35758
rect 43932 36594 43988 36596
rect 43932 36542 43934 36594
rect 43934 36542 43986 36594
rect 43986 36542 43988 36594
rect 43932 36540 43988 36542
rect 44132 36090 44188 36092
rect 44132 36038 44134 36090
rect 44134 36038 44186 36090
rect 44186 36038 44188 36090
rect 44132 36036 44188 36038
rect 44236 36090 44292 36092
rect 44236 36038 44238 36090
rect 44238 36038 44290 36090
rect 44290 36038 44292 36090
rect 44236 36036 44292 36038
rect 44340 36090 44396 36092
rect 44340 36038 44342 36090
rect 44342 36038 44394 36090
rect 44394 36038 44396 36090
rect 44340 36036 44396 36038
rect 42812 35196 42868 35252
rect 42924 34914 42980 34916
rect 42924 34862 42926 34914
rect 42926 34862 42978 34914
rect 42978 34862 42980 34914
rect 42924 34860 42980 34862
rect 44828 35532 44884 35588
rect 43820 34748 43876 34804
rect 45836 37324 45892 37380
rect 45612 35586 45668 35588
rect 45612 35534 45614 35586
rect 45614 35534 45666 35586
rect 45666 35534 45668 35586
rect 45612 35532 45668 35534
rect 45500 34860 45556 34916
rect 46732 36482 46788 36484
rect 46732 36430 46734 36482
rect 46734 36430 46786 36482
rect 46786 36430 46788 36482
rect 46732 36428 46788 36430
rect 46060 36370 46116 36372
rect 46060 36318 46062 36370
rect 46062 36318 46114 36370
rect 46114 36318 46116 36370
rect 46060 36316 46116 36318
rect 47740 36428 47796 36484
rect 48860 36482 48916 36484
rect 48860 36430 48862 36482
rect 48862 36430 48914 36482
rect 48914 36430 48916 36482
rect 48860 36428 48916 36430
rect 46732 35868 46788 35924
rect 46844 35980 46900 36036
rect 44132 34522 44188 34524
rect 44132 34470 44134 34522
rect 44134 34470 44186 34522
rect 44186 34470 44188 34522
rect 44132 34468 44188 34470
rect 44236 34522 44292 34524
rect 44236 34470 44238 34522
rect 44238 34470 44290 34522
rect 44290 34470 44292 34522
rect 44236 34468 44292 34470
rect 44340 34522 44396 34524
rect 44340 34470 44342 34522
rect 44342 34470 44394 34522
rect 44394 34470 44396 34522
rect 44340 34468 44396 34470
rect 46060 35644 46116 35700
rect 46284 35532 46340 35588
rect 45836 34636 45892 34692
rect 43820 33740 43876 33796
rect 43932 33346 43988 33348
rect 43932 33294 43934 33346
rect 43934 33294 43986 33346
rect 43986 33294 43988 33346
rect 43932 33292 43988 33294
rect 43708 33234 43764 33236
rect 43708 33182 43710 33234
rect 43710 33182 43762 33234
rect 43762 33182 43764 33234
rect 43708 33180 43764 33182
rect 44132 32954 44188 32956
rect 43372 32844 43428 32900
rect 44132 32902 44134 32954
rect 44134 32902 44186 32954
rect 44186 32902 44188 32954
rect 44132 32900 44188 32902
rect 44236 32954 44292 32956
rect 44236 32902 44238 32954
rect 44238 32902 44290 32954
rect 44290 32902 44292 32954
rect 44236 32900 44292 32902
rect 44340 32954 44396 32956
rect 44340 32902 44342 32954
rect 44342 32902 44394 32954
rect 44394 32902 44396 32954
rect 44340 32900 44396 32902
rect 43932 32786 43988 32788
rect 43932 32734 43934 32786
rect 43934 32734 43986 32786
rect 43986 32734 43988 32786
rect 43932 32732 43988 32734
rect 43932 32508 43988 32564
rect 42700 32284 42756 32340
rect 42588 31612 42644 31668
rect 42588 29932 42644 29988
rect 42700 30940 42756 30996
rect 42364 27746 42420 27748
rect 42364 27694 42366 27746
rect 42366 27694 42418 27746
rect 42418 27694 42420 27746
rect 42364 27692 42420 27694
rect 44044 32060 44100 32116
rect 43708 31890 43764 31892
rect 43708 31838 43710 31890
rect 43710 31838 43762 31890
rect 43762 31838 43764 31890
rect 43708 31836 43764 31838
rect 45164 32732 45220 32788
rect 44828 32562 44884 32564
rect 44828 32510 44830 32562
rect 44830 32510 44882 32562
rect 44882 32510 44884 32562
rect 44828 32508 44884 32510
rect 43148 31612 43204 31668
rect 43036 30604 43092 30660
rect 42812 30098 42868 30100
rect 42812 30046 42814 30098
rect 42814 30046 42866 30098
rect 42866 30046 42868 30098
rect 42812 30044 42868 30046
rect 44132 31386 44188 31388
rect 44132 31334 44134 31386
rect 44134 31334 44186 31386
rect 44186 31334 44188 31386
rect 44132 31332 44188 31334
rect 44236 31386 44292 31388
rect 44236 31334 44238 31386
rect 44238 31334 44290 31386
rect 44290 31334 44292 31386
rect 44236 31332 44292 31334
rect 44340 31386 44396 31388
rect 44340 31334 44342 31386
rect 44342 31334 44394 31386
rect 44394 31334 44396 31386
rect 44340 31332 44396 31334
rect 46284 33346 46340 33348
rect 46284 33294 46286 33346
rect 46286 33294 46338 33346
rect 46338 33294 46340 33346
rect 46284 33292 46340 33294
rect 47628 35308 47684 35364
rect 47292 35196 47348 35252
rect 47516 35084 47572 35140
rect 46844 34802 46900 34804
rect 46844 34750 46846 34802
rect 46846 34750 46898 34802
rect 46898 34750 46900 34802
rect 46844 34748 46900 34750
rect 46732 33292 46788 33348
rect 47292 33234 47348 33236
rect 47292 33182 47294 33234
rect 47294 33182 47346 33234
rect 47346 33182 47348 33234
rect 47292 33180 47348 33182
rect 45388 32450 45444 32452
rect 45388 32398 45390 32450
rect 45390 32398 45442 32450
rect 45442 32398 45444 32450
rect 45388 32396 45444 32398
rect 45724 32172 45780 32228
rect 45612 31948 45668 32004
rect 45500 31836 45556 31892
rect 45052 31778 45108 31780
rect 45052 31726 45054 31778
rect 45054 31726 45106 31778
rect 45106 31726 45108 31778
rect 45052 31724 45108 31726
rect 45388 31724 45444 31780
rect 43932 30994 43988 30996
rect 43932 30942 43934 30994
rect 43934 30942 43986 30994
rect 43986 30942 43988 30994
rect 43932 30940 43988 30942
rect 43484 29932 43540 29988
rect 42812 29538 42868 29540
rect 42812 29486 42814 29538
rect 42814 29486 42866 29538
rect 42866 29486 42868 29538
rect 42812 29484 42868 29486
rect 44492 30770 44548 30772
rect 44492 30718 44494 30770
rect 44494 30718 44546 30770
rect 44546 30718 44548 30770
rect 44492 30716 44548 30718
rect 44828 30380 44884 30436
rect 44604 30268 44660 30324
rect 43596 28924 43652 28980
rect 43372 28812 43428 28868
rect 43372 27858 43428 27860
rect 43372 27806 43374 27858
rect 43374 27806 43426 27858
rect 43426 27806 43428 27858
rect 43372 27804 43428 27806
rect 43372 27580 43428 27636
rect 41916 25004 41972 25060
rect 42252 26908 42308 26964
rect 41916 24834 41972 24836
rect 41916 24782 41918 24834
rect 41918 24782 41970 24834
rect 41970 24782 41972 24834
rect 41916 24780 41972 24782
rect 43260 26908 43316 26964
rect 42476 25116 42532 25172
rect 43484 26796 43540 26852
rect 44132 29818 44188 29820
rect 44132 29766 44134 29818
rect 44134 29766 44186 29818
rect 44186 29766 44188 29818
rect 44132 29764 44188 29766
rect 44236 29818 44292 29820
rect 44236 29766 44238 29818
rect 44238 29766 44290 29818
rect 44290 29766 44292 29818
rect 44236 29764 44292 29766
rect 44340 29818 44396 29820
rect 44340 29766 44342 29818
rect 44342 29766 44394 29818
rect 44394 29766 44396 29818
rect 44340 29764 44396 29766
rect 44156 29426 44212 29428
rect 44156 29374 44158 29426
rect 44158 29374 44210 29426
rect 44210 29374 44212 29426
rect 44156 29372 44212 29374
rect 44044 28924 44100 28980
rect 43932 28700 43988 28756
rect 43596 25676 43652 25732
rect 43596 25452 43652 25508
rect 42812 24834 42868 24836
rect 42812 24782 42814 24834
rect 42814 24782 42866 24834
rect 42866 24782 42868 24834
rect 42812 24780 42868 24782
rect 42924 24722 42980 24724
rect 42924 24670 42926 24722
rect 42926 24670 42978 24722
rect 42978 24670 42980 24722
rect 42924 24668 42980 24670
rect 41692 23548 41748 23604
rect 41468 22092 41524 22148
rect 41692 22930 41748 22932
rect 41692 22878 41694 22930
rect 41694 22878 41746 22930
rect 41746 22878 41748 22930
rect 41692 22876 41748 22878
rect 41692 22092 41748 22148
rect 41468 20972 41524 21028
rect 41244 20860 41300 20916
rect 40796 20578 40852 20580
rect 40796 20526 40798 20578
rect 40798 20526 40850 20578
rect 40850 20526 40852 20578
rect 40796 20524 40852 20526
rect 40460 19292 40516 19348
rect 40684 19740 40740 19796
rect 40124 18172 40180 18228
rect 40348 17778 40404 17780
rect 40348 17726 40350 17778
rect 40350 17726 40402 17778
rect 40402 17726 40404 17778
rect 40348 17724 40404 17726
rect 40236 16940 40292 16996
rect 40460 16098 40516 16100
rect 40460 16046 40462 16098
rect 40462 16046 40514 16098
rect 40514 16046 40516 16098
rect 40460 16044 40516 16046
rect 39564 15484 39620 15540
rect 39340 14924 39396 14980
rect 40012 15372 40068 15428
rect 39340 14476 39396 14532
rect 39228 14418 39284 14420
rect 39228 14366 39230 14418
rect 39230 14366 39282 14418
rect 39282 14366 39284 14418
rect 39228 14364 39284 14366
rect 38780 14252 38836 14308
rect 38556 12962 38612 12964
rect 38556 12910 38558 12962
rect 38558 12910 38610 12962
rect 38610 12910 38612 12962
rect 38556 12908 38612 12910
rect 38556 10668 38612 10724
rect 39340 13468 39396 13524
rect 39340 12012 39396 12068
rect 39228 11788 39284 11844
rect 38780 11340 38836 11396
rect 39340 10668 39396 10724
rect 38892 10610 38948 10612
rect 38892 10558 38894 10610
rect 38894 10558 38946 10610
rect 38946 10558 38948 10610
rect 38892 10556 38948 10558
rect 38668 10108 38724 10164
rect 39676 14476 39732 14532
rect 41020 19628 41076 19684
rect 41916 20972 41972 21028
rect 41580 20524 41636 20580
rect 42028 20690 42084 20692
rect 42028 20638 42030 20690
rect 42030 20638 42082 20690
rect 42082 20638 42084 20690
rect 42028 20636 42084 20638
rect 41356 19010 41412 19012
rect 41356 18958 41358 19010
rect 41358 18958 41410 19010
rect 41410 18958 41412 19010
rect 41356 18956 41412 18958
rect 40908 16828 40964 16884
rect 41132 17836 41188 17892
rect 40684 15260 40740 15316
rect 40796 16716 40852 16772
rect 40236 14700 40292 14756
rect 40348 14530 40404 14532
rect 40348 14478 40350 14530
rect 40350 14478 40402 14530
rect 40402 14478 40404 14530
rect 40348 14476 40404 14478
rect 40908 16492 40964 16548
rect 41468 17836 41524 17892
rect 41244 16994 41300 16996
rect 41244 16942 41246 16994
rect 41246 16942 41298 16994
rect 41298 16942 41300 16994
rect 41244 16940 41300 16942
rect 41132 16882 41188 16884
rect 41132 16830 41134 16882
rect 41134 16830 41186 16882
rect 41186 16830 41188 16882
rect 41132 16828 41188 16830
rect 41468 16716 41524 16772
rect 40908 16156 40964 16212
rect 40908 15596 40964 15652
rect 41020 15538 41076 15540
rect 41020 15486 41022 15538
rect 41022 15486 41074 15538
rect 41074 15486 41076 15538
rect 41020 15484 41076 15486
rect 41244 15314 41300 15316
rect 41244 15262 41246 15314
rect 41246 15262 41298 15314
rect 41298 15262 41300 15314
rect 41244 15260 41300 15262
rect 41132 14530 41188 14532
rect 41132 14478 41134 14530
rect 41134 14478 41186 14530
rect 41186 14478 41188 14530
rect 41132 14476 41188 14478
rect 39788 13634 39844 13636
rect 39788 13582 39790 13634
rect 39790 13582 39842 13634
rect 39842 13582 39844 13634
rect 39788 13580 39844 13582
rect 40012 13522 40068 13524
rect 40012 13470 40014 13522
rect 40014 13470 40066 13522
rect 40066 13470 40068 13522
rect 40012 13468 40068 13470
rect 41132 13634 41188 13636
rect 41132 13582 41134 13634
rect 41134 13582 41186 13634
rect 41186 13582 41188 13634
rect 41132 13580 41188 13582
rect 40012 12796 40068 12852
rect 40124 12290 40180 12292
rect 40124 12238 40126 12290
rect 40126 12238 40178 12290
rect 40178 12238 40180 12290
rect 40124 12236 40180 12238
rect 41132 12796 41188 12852
rect 41132 12236 41188 12292
rect 39564 11506 39620 11508
rect 39564 11454 39566 11506
rect 39566 11454 39618 11506
rect 39618 11454 39620 11506
rect 39564 11452 39620 11454
rect 39564 10780 39620 10836
rect 41020 12066 41076 12068
rect 41020 12014 41022 12066
rect 41022 12014 41074 12066
rect 41074 12014 41076 12066
rect 41020 12012 41076 12014
rect 39452 9996 39508 10052
rect 39004 9324 39060 9380
rect 39452 9100 39508 9156
rect 38668 8818 38724 8820
rect 38668 8766 38670 8818
rect 38670 8766 38722 8818
rect 38722 8766 38724 8818
rect 38668 8764 38724 8766
rect 38780 8428 38836 8484
rect 38556 8092 38612 8148
rect 38668 7868 38724 7924
rect 38892 8316 38948 8372
rect 41356 13356 41412 13412
rect 39900 9660 39956 9716
rect 39676 9548 39732 9604
rect 39452 7644 39508 7700
rect 40348 9324 40404 9380
rect 40012 9154 40068 9156
rect 40012 9102 40014 9154
rect 40014 9102 40066 9154
rect 40066 9102 40068 9154
rect 40012 9100 40068 9102
rect 40908 10610 40964 10612
rect 40908 10558 40910 10610
rect 40910 10558 40962 10610
rect 40962 10558 40964 10610
rect 40908 10556 40964 10558
rect 41244 11676 41300 11732
rect 41132 10498 41188 10500
rect 41132 10446 41134 10498
rect 41134 10446 41186 10498
rect 41186 10446 41188 10498
rect 41132 10444 41188 10446
rect 41468 10498 41524 10500
rect 41468 10446 41470 10498
rect 41470 10446 41522 10498
rect 41522 10446 41524 10498
rect 41468 10444 41524 10446
rect 41804 19180 41860 19236
rect 42028 18956 42084 19012
rect 42028 18450 42084 18452
rect 42028 18398 42030 18450
rect 42030 18398 42082 18450
rect 42082 18398 42084 18450
rect 42028 18396 42084 18398
rect 42028 16828 42084 16884
rect 42700 23660 42756 23716
rect 43820 27804 43876 27860
rect 44268 28642 44324 28644
rect 44268 28590 44270 28642
rect 44270 28590 44322 28642
rect 44322 28590 44324 28642
rect 44268 28588 44324 28590
rect 44132 28250 44188 28252
rect 44132 28198 44134 28250
rect 44134 28198 44186 28250
rect 44186 28198 44188 28250
rect 44132 28196 44188 28198
rect 44236 28250 44292 28252
rect 44236 28198 44238 28250
rect 44238 28198 44290 28250
rect 44290 28198 44292 28250
rect 44236 28196 44292 28198
rect 44340 28250 44396 28252
rect 44340 28198 44342 28250
rect 44342 28198 44394 28250
rect 44394 28198 44396 28250
rect 44340 28196 44396 28198
rect 44268 27858 44324 27860
rect 44268 27806 44270 27858
rect 44270 27806 44322 27858
rect 44322 27806 44324 27858
rect 44268 27804 44324 27806
rect 43932 27692 43988 27748
rect 44716 28812 44772 28868
rect 45948 31106 46004 31108
rect 45948 31054 45950 31106
rect 45950 31054 46002 31106
rect 46002 31054 46004 31106
rect 45948 31052 46004 31054
rect 45500 30716 45556 30772
rect 44940 29596 44996 29652
rect 45724 30156 45780 30212
rect 44940 28924 44996 28980
rect 44828 28364 44884 28420
rect 45052 27746 45108 27748
rect 45052 27694 45054 27746
rect 45054 27694 45106 27746
rect 45106 27694 45108 27746
rect 45052 27692 45108 27694
rect 44940 27020 44996 27076
rect 44132 26682 44188 26684
rect 44132 26630 44134 26682
rect 44134 26630 44186 26682
rect 44186 26630 44188 26682
rect 44132 26628 44188 26630
rect 44236 26682 44292 26684
rect 44236 26630 44238 26682
rect 44238 26630 44290 26682
rect 44290 26630 44292 26682
rect 44236 26628 44292 26630
rect 44340 26682 44396 26684
rect 44340 26630 44342 26682
rect 44342 26630 44394 26682
rect 44394 26630 44396 26682
rect 44340 26628 44396 26630
rect 44492 26402 44548 26404
rect 44492 26350 44494 26402
rect 44494 26350 44546 26402
rect 44546 26350 44548 26402
rect 44492 26348 44548 26350
rect 44604 26290 44660 26292
rect 44604 26238 44606 26290
rect 44606 26238 44658 26290
rect 44658 26238 44660 26290
rect 44604 26236 44660 26238
rect 43932 25676 43988 25732
rect 44132 25114 44188 25116
rect 44132 25062 44134 25114
rect 44134 25062 44186 25114
rect 44186 25062 44188 25114
rect 44132 25060 44188 25062
rect 44236 25114 44292 25116
rect 44236 25062 44238 25114
rect 44238 25062 44290 25114
rect 44290 25062 44292 25114
rect 44236 25060 44292 25062
rect 44340 25114 44396 25116
rect 44340 25062 44342 25114
rect 44342 25062 44394 25114
rect 44394 25062 44396 25114
rect 44340 25060 44396 25062
rect 43932 24892 43988 24948
rect 44044 24668 44100 24724
rect 43932 24332 43988 24388
rect 43596 23996 43652 24052
rect 43932 23996 43988 24052
rect 43708 23884 43764 23940
rect 42812 23378 42868 23380
rect 42812 23326 42814 23378
rect 42814 23326 42866 23378
rect 42866 23326 42868 23378
rect 42812 23324 42868 23326
rect 43260 23324 43316 23380
rect 42924 23100 42980 23156
rect 42588 22876 42644 22932
rect 42364 19964 42420 20020
rect 42924 21586 42980 21588
rect 42924 21534 42926 21586
rect 42926 21534 42978 21586
rect 42978 21534 42980 21586
rect 42924 21532 42980 21534
rect 43484 23436 43540 23492
rect 43820 23436 43876 23492
rect 43148 21308 43204 21364
rect 42924 20524 42980 20580
rect 42700 18674 42756 18676
rect 42700 18622 42702 18674
rect 42702 18622 42754 18674
rect 42754 18622 42756 18674
rect 42700 18620 42756 18622
rect 44132 23546 44188 23548
rect 44132 23494 44134 23546
rect 44134 23494 44186 23546
rect 44186 23494 44188 23546
rect 44132 23492 44188 23494
rect 44236 23546 44292 23548
rect 44236 23494 44238 23546
rect 44238 23494 44290 23546
rect 44290 23494 44292 23546
rect 44236 23492 44292 23494
rect 44340 23546 44396 23548
rect 44340 23494 44342 23546
rect 44342 23494 44394 23546
rect 44394 23494 44396 23546
rect 44340 23492 44396 23494
rect 44380 22930 44436 22932
rect 44380 22878 44382 22930
rect 44382 22878 44434 22930
rect 44434 22878 44436 22930
rect 44380 22876 44436 22878
rect 44044 22428 44100 22484
rect 45500 29596 45556 29652
rect 45276 28642 45332 28644
rect 45276 28590 45278 28642
rect 45278 28590 45330 28642
rect 45330 28590 45332 28642
rect 45276 28588 45332 28590
rect 45724 29538 45780 29540
rect 45724 29486 45726 29538
rect 45726 29486 45778 29538
rect 45778 29486 45780 29538
rect 45724 29484 45780 29486
rect 46620 31836 46676 31892
rect 46284 31724 46340 31780
rect 47180 32060 47236 32116
rect 46956 32002 47012 32004
rect 46956 31950 46958 32002
rect 46958 31950 47010 32002
rect 47010 31950 47012 32002
rect 46956 31948 47012 31950
rect 46844 31612 46900 31668
rect 47516 33292 47572 33348
rect 48300 36204 48356 36260
rect 48748 35810 48804 35812
rect 48748 35758 48750 35810
rect 48750 35758 48802 35810
rect 48802 35758 48804 35810
rect 48748 35756 48804 35758
rect 49196 36370 49252 36372
rect 49196 36318 49198 36370
rect 49198 36318 49250 36370
rect 49250 36318 49252 36370
rect 49196 36316 49252 36318
rect 52108 36988 52164 37044
rect 51286 36874 51342 36876
rect 51286 36822 51288 36874
rect 51288 36822 51340 36874
rect 51340 36822 51342 36874
rect 51286 36820 51342 36822
rect 51390 36874 51446 36876
rect 51390 36822 51392 36874
rect 51392 36822 51444 36874
rect 51444 36822 51446 36874
rect 51390 36820 51446 36822
rect 51494 36874 51550 36876
rect 51494 36822 51496 36874
rect 51496 36822 51548 36874
rect 51548 36822 51550 36874
rect 51494 36820 51550 36822
rect 49980 36316 50036 36372
rect 50540 36370 50596 36372
rect 50540 36318 50542 36370
rect 50542 36318 50594 36370
rect 50594 36318 50596 36370
rect 50540 36316 50596 36318
rect 49308 36092 49364 36148
rect 48860 35532 48916 35588
rect 49084 35810 49140 35812
rect 49084 35758 49086 35810
rect 49086 35758 49138 35810
rect 49138 35758 49140 35810
rect 49084 35756 49140 35758
rect 47964 34860 48020 34916
rect 47740 34130 47796 34132
rect 47740 34078 47742 34130
rect 47742 34078 47794 34130
rect 47794 34078 47796 34130
rect 47740 34076 47796 34078
rect 48972 34972 49028 35028
rect 48188 34636 48244 34692
rect 48748 34130 48804 34132
rect 48748 34078 48750 34130
rect 48750 34078 48802 34130
rect 48802 34078 48804 34130
rect 48748 34076 48804 34078
rect 51436 35922 51492 35924
rect 51436 35870 51438 35922
rect 51438 35870 51490 35922
rect 51490 35870 51492 35922
rect 51436 35868 51492 35870
rect 50204 35644 50260 35700
rect 49196 35420 49252 35476
rect 49420 35420 49476 35476
rect 49868 34802 49924 34804
rect 49868 34750 49870 34802
rect 49870 34750 49922 34802
rect 49922 34750 49924 34802
rect 49868 34748 49924 34750
rect 49980 34412 50036 34468
rect 47964 33852 48020 33908
rect 47628 33516 47684 33572
rect 48188 33346 48244 33348
rect 48188 33294 48190 33346
rect 48190 33294 48242 33346
rect 48242 33294 48244 33346
rect 48188 33292 48244 33294
rect 48860 33628 48916 33684
rect 48748 33180 48804 33236
rect 47628 33068 47684 33124
rect 48524 33068 48580 33124
rect 46396 29596 46452 29652
rect 46284 29372 46340 29428
rect 46060 29260 46116 29316
rect 45724 28700 45780 28756
rect 45276 28364 45332 28420
rect 45276 27468 45332 27524
rect 45500 28252 45556 28308
rect 45500 27858 45556 27860
rect 45500 27806 45502 27858
rect 45502 27806 45554 27858
rect 45554 27806 45556 27858
rect 45500 27804 45556 27806
rect 46396 28754 46452 28756
rect 46396 28702 46398 28754
rect 46398 28702 46450 28754
rect 46450 28702 46452 28754
rect 46396 28700 46452 28702
rect 46284 28252 46340 28308
rect 45948 27858 46004 27860
rect 45948 27806 45950 27858
rect 45950 27806 46002 27858
rect 46002 27806 46004 27858
rect 45948 27804 46004 27806
rect 46620 27468 46676 27524
rect 46956 27298 47012 27300
rect 46956 27246 46958 27298
rect 46958 27246 47010 27298
rect 47010 27246 47012 27298
rect 46956 27244 47012 27246
rect 46844 27132 46900 27188
rect 45500 27020 45556 27076
rect 46284 27074 46340 27076
rect 46284 27022 46286 27074
rect 46286 27022 46338 27074
rect 46338 27022 46340 27074
rect 46284 27020 46340 27022
rect 46620 26402 46676 26404
rect 46620 26350 46622 26402
rect 46622 26350 46674 26402
rect 46674 26350 46676 26402
rect 46620 26348 46676 26350
rect 45948 26236 46004 26292
rect 45052 24722 45108 24724
rect 45052 24670 45054 24722
rect 45054 24670 45106 24722
rect 45106 24670 45108 24722
rect 45052 24668 45108 24670
rect 44492 22428 44548 22484
rect 45052 24444 45108 24500
rect 45164 23996 45220 24052
rect 45276 24892 45332 24948
rect 45948 25340 46004 25396
rect 45836 24892 45892 24948
rect 46956 26178 47012 26180
rect 46956 26126 46958 26178
rect 46958 26126 47010 26178
rect 47010 26126 47012 26178
rect 46956 26124 47012 26126
rect 48188 31778 48244 31780
rect 48188 31726 48190 31778
rect 48190 31726 48242 31778
rect 48242 31726 48244 31778
rect 48188 31724 48244 31726
rect 48076 30828 48132 30884
rect 47180 30210 47236 30212
rect 47180 30158 47182 30210
rect 47182 30158 47234 30210
rect 47234 30158 47236 30210
rect 47180 30156 47236 30158
rect 47964 29820 48020 29876
rect 48188 30716 48244 30772
rect 48748 32674 48804 32676
rect 48748 32622 48750 32674
rect 48750 32622 48802 32674
rect 48802 32622 48804 32674
rect 48748 32620 48804 32622
rect 49308 31948 49364 32004
rect 49084 31836 49140 31892
rect 48860 31724 48916 31780
rect 50092 33516 50148 33572
rect 51772 35810 51828 35812
rect 51772 35758 51774 35810
rect 51774 35758 51826 35810
rect 51826 35758 51828 35810
rect 51772 35756 51828 35758
rect 50876 35586 50932 35588
rect 50876 35534 50878 35586
rect 50878 35534 50930 35586
rect 50930 35534 50932 35586
rect 50876 35532 50932 35534
rect 52220 36428 52276 36484
rect 52780 35868 52836 35924
rect 51286 35306 51342 35308
rect 51286 35254 51288 35306
rect 51288 35254 51340 35306
rect 51340 35254 51342 35306
rect 51286 35252 51342 35254
rect 51390 35306 51446 35308
rect 51390 35254 51392 35306
rect 51392 35254 51444 35306
rect 51444 35254 51446 35306
rect 51390 35252 51446 35254
rect 51494 35306 51550 35308
rect 51494 35254 51496 35306
rect 51496 35254 51548 35306
rect 51548 35254 51550 35306
rect 51494 35252 51550 35254
rect 51212 35026 51268 35028
rect 51212 34974 51214 35026
rect 51214 34974 51266 35026
rect 51266 34974 51268 35026
rect 51212 34972 51268 34974
rect 52780 35532 52836 35588
rect 53788 36482 53844 36484
rect 53788 36430 53790 36482
rect 53790 36430 53842 36482
rect 53842 36430 53844 36482
rect 53788 36428 53844 36430
rect 56252 37212 56308 37268
rect 55020 36652 55076 36708
rect 54460 36428 54516 36484
rect 55468 36482 55524 36484
rect 55468 36430 55470 36482
rect 55470 36430 55522 36482
rect 55522 36430 55524 36482
rect 55468 36428 55524 36430
rect 53564 35980 53620 36036
rect 52892 34972 52948 35028
rect 54684 35922 54740 35924
rect 54684 35870 54686 35922
rect 54686 35870 54738 35922
rect 54738 35870 54740 35922
rect 54684 35868 54740 35870
rect 51548 34802 51604 34804
rect 51548 34750 51550 34802
rect 51550 34750 51602 34802
rect 51602 34750 51604 34802
rect 51548 34748 51604 34750
rect 50652 34636 50708 34692
rect 50988 34636 51044 34692
rect 50540 34412 50596 34468
rect 50540 34076 50596 34132
rect 50204 33628 50260 33684
rect 50540 33740 50596 33796
rect 50428 33234 50484 33236
rect 50428 33182 50430 33234
rect 50430 33182 50482 33234
rect 50482 33182 50484 33234
rect 50428 33180 50484 33182
rect 51660 34690 51716 34692
rect 51660 34638 51662 34690
rect 51662 34638 51714 34690
rect 51714 34638 51716 34690
rect 51660 34636 51716 34638
rect 51884 34300 51940 34356
rect 51548 34130 51604 34132
rect 51548 34078 51550 34130
rect 51550 34078 51602 34130
rect 51602 34078 51604 34130
rect 51548 34076 51604 34078
rect 50988 33740 51044 33796
rect 51286 33738 51342 33740
rect 51286 33686 51288 33738
rect 51288 33686 51340 33738
rect 51340 33686 51342 33738
rect 51286 33684 51342 33686
rect 51390 33738 51446 33740
rect 51390 33686 51392 33738
rect 51392 33686 51444 33738
rect 51444 33686 51446 33738
rect 51390 33684 51446 33686
rect 51494 33738 51550 33740
rect 51494 33686 51496 33738
rect 51496 33686 51548 33738
rect 51548 33686 51550 33738
rect 51494 33684 51550 33686
rect 51212 33570 51268 33572
rect 51212 33518 51214 33570
rect 51214 33518 51266 33570
rect 51266 33518 51268 33570
rect 51212 33516 51268 33518
rect 51548 33516 51604 33572
rect 49532 31948 49588 32004
rect 50204 31948 50260 32004
rect 48972 29820 49028 29876
rect 48188 29202 48244 29204
rect 48188 29150 48190 29202
rect 48190 29150 48242 29202
rect 48242 29150 48244 29202
rect 48188 29148 48244 29150
rect 48972 29650 49028 29652
rect 48972 29598 48974 29650
rect 48974 29598 49026 29650
rect 49026 29598 49028 29650
rect 48972 29596 49028 29598
rect 47852 27858 47908 27860
rect 47852 27806 47854 27858
rect 47854 27806 47906 27858
rect 47906 27806 47908 27858
rect 47852 27804 47908 27806
rect 48076 27858 48132 27860
rect 48076 27806 48078 27858
rect 48078 27806 48130 27858
rect 48130 27806 48132 27858
rect 48076 27804 48132 27806
rect 47516 27356 47572 27412
rect 47180 27132 47236 27188
rect 47292 27020 47348 27076
rect 47068 26012 47124 26068
rect 47740 27298 47796 27300
rect 47740 27246 47742 27298
rect 47742 27246 47794 27298
rect 47794 27246 47796 27298
rect 47740 27244 47796 27246
rect 47852 27074 47908 27076
rect 47852 27022 47854 27074
rect 47854 27022 47906 27074
rect 47906 27022 47908 27074
rect 47852 27020 47908 27022
rect 47516 26572 47572 26628
rect 46172 25618 46228 25620
rect 46172 25566 46174 25618
rect 46174 25566 46226 25618
rect 46226 25566 46228 25618
rect 46172 25564 46228 25566
rect 46060 24668 46116 24724
rect 45052 23884 45108 23940
rect 44380 22370 44436 22372
rect 44380 22318 44382 22370
rect 44382 22318 44434 22370
rect 44434 22318 44436 22370
rect 44380 22316 44436 22318
rect 44132 21978 44188 21980
rect 44132 21926 44134 21978
rect 44134 21926 44186 21978
rect 44186 21926 44188 21978
rect 44132 21924 44188 21926
rect 44236 21978 44292 21980
rect 44236 21926 44238 21978
rect 44238 21926 44290 21978
rect 44290 21926 44292 21978
rect 44236 21924 44292 21926
rect 44340 21978 44396 21980
rect 44340 21926 44342 21978
rect 44342 21926 44394 21978
rect 44394 21926 44396 21978
rect 44340 21924 44396 21926
rect 44492 21586 44548 21588
rect 44492 21534 44494 21586
rect 44494 21534 44546 21586
rect 44546 21534 44548 21586
rect 44492 21532 44548 21534
rect 44380 20860 44436 20916
rect 44132 20410 44188 20412
rect 44132 20358 44134 20410
rect 44134 20358 44186 20410
rect 44186 20358 44188 20410
rect 44132 20356 44188 20358
rect 44236 20410 44292 20412
rect 44236 20358 44238 20410
rect 44238 20358 44290 20410
rect 44290 20358 44292 20410
rect 44236 20356 44292 20358
rect 44340 20410 44396 20412
rect 44340 20358 44342 20410
rect 44342 20358 44394 20410
rect 44394 20358 44396 20410
rect 44340 20356 44396 20358
rect 43932 20076 43988 20132
rect 43260 19964 43316 20020
rect 42924 18284 42980 18340
rect 43260 19234 43316 19236
rect 43260 19182 43262 19234
rect 43262 19182 43314 19234
rect 43314 19182 43316 19234
rect 43260 19180 43316 19182
rect 44044 19964 44100 20020
rect 43932 19740 43988 19796
rect 43260 18284 43316 18340
rect 42924 17836 42980 17892
rect 42252 16716 42308 16772
rect 42364 16322 42420 16324
rect 42364 16270 42366 16322
rect 42366 16270 42418 16322
rect 42418 16270 42420 16322
rect 42364 16268 42420 16270
rect 41804 15426 41860 15428
rect 41804 15374 41806 15426
rect 41806 15374 41858 15426
rect 41858 15374 41860 15426
rect 41804 15372 41860 15374
rect 41916 13020 41972 13076
rect 42140 15314 42196 15316
rect 42140 15262 42142 15314
rect 42142 15262 42194 15314
rect 42194 15262 42196 15314
rect 42140 15260 42196 15262
rect 43148 17724 43204 17780
rect 43036 17164 43092 17220
rect 44132 18842 44188 18844
rect 44132 18790 44134 18842
rect 44134 18790 44186 18842
rect 44186 18790 44188 18842
rect 44132 18788 44188 18790
rect 44236 18842 44292 18844
rect 44236 18790 44238 18842
rect 44238 18790 44290 18842
rect 44290 18790 44292 18842
rect 44236 18788 44292 18790
rect 44340 18842 44396 18844
rect 44340 18790 44342 18842
rect 44342 18790 44394 18842
rect 44394 18790 44396 18842
rect 44340 18788 44396 18790
rect 44492 18620 44548 18676
rect 44716 23660 44772 23716
rect 44828 23436 44884 23492
rect 44828 21474 44884 21476
rect 44828 21422 44830 21474
rect 44830 21422 44882 21474
rect 44882 21422 44884 21474
rect 44828 21420 44884 21422
rect 45836 23884 45892 23940
rect 47068 25618 47124 25620
rect 47068 25566 47070 25618
rect 47070 25566 47122 25618
rect 47122 25566 47124 25618
rect 47068 25564 47124 25566
rect 46508 25394 46564 25396
rect 46508 25342 46510 25394
rect 46510 25342 46562 25394
rect 46562 25342 46564 25394
rect 46508 25340 46564 25342
rect 46620 24892 46676 24948
rect 46396 24668 46452 24724
rect 46508 24108 46564 24164
rect 45948 23660 46004 23716
rect 45724 23548 45780 23604
rect 45276 23436 45332 23492
rect 45276 23266 45332 23268
rect 45276 23214 45278 23266
rect 45278 23214 45330 23266
rect 45330 23214 45332 23266
rect 45276 23212 45332 23214
rect 45164 22204 45220 22260
rect 44716 20076 44772 20132
rect 44828 19068 44884 19124
rect 44380 18450 44436 18452
rect 44380 18398 44382 18450
rect 44382 18398 44434 18450
rect 44434 18398 44436 18450
rect 44380 18396 44436 18398
rect 44156 18338 44212 18340
rect 44156 18286 44158 18338
rect 44158 18286 44210 18338
rect 44210 18286 44212 18338
rect 44156 18284 44212 18286
rect 43820 17612 43876 17668
rect 42700 16882 42756 16884
rect 42700 16830 42702 16882
rect 42702 16830 42754 16882
rect 42754 16830 42756 16882
rect 42700 16828 42756 16830
rect 42924 16268 42980 16324
rect 44132 17274 44188 17276
rect 44132 17222 44134 17274
rect 44134 17222 44186 17274
rect 44186 17222 44188 17274
rect 44132 17220 44188 17222
rect 44236 17274 44292 17276
rect 44236 17222 44238 17274
rect 44238 17222 44290 17274
rect 44290 17222 44292 17274
rect 44236 17220 44292 17222
rect 44340 17274 44396 17276
rect 44340 17222 44342 17274
rect 44342 17222 44394 17274
rect 44394 17222 44396 17274
rect 44340 17220 44396 17222
rect 43932 16716 43988 16772
rect 44156 16268 44212 16324
rect 44132 15706 44188 15708
rect 44132 15654 44134 15706
rect 44134 15654 44186 15706
rect 44186 15654 44188 15706
rect 44132 15652 44188 15654
rect 44236 15706 44292 15708
rect 44236 15654 44238 15706
rect 44238 15654 44290 15706
rect 44290 15654 44292 15706
rect 44236 15652 44292 15654
rect 44340 15706 44396 15708
rect 44340 15654 44342 15706
rect 44342 15654 44394 15706
rect 44394 15654 44396 15706
rect 44340 15652 44396 15654
rect 44268 15484 44324 15540
rect 43820 15148 43876 15204
rect 42476 15090 42532 15092
rect 42476 15038 42478 15090
rect 42478 15038 42530 15090
rect 42530 15038 42532 15090
rect 42476 15036 42532 15038
rect 42476 13468 42532 13524
rect 43932 14588 43988 14644
rect 44268 14530 44324 14532
rect 44268 14478 44270 14530
rect 44270 14478 44322 14530
rect 44322 14478 44324 14530
rect 44268 14476 44324 14478
rect 42812 14140 42868 14196
rect 42476 11788 42532 11844
rect 42028 11676 42084 11732
rect 41692 10668 41748 10724
rect 41804 10780 41860 10836
rect 42252 10332 42308 10388
rect 40684 9714 40740 9716
rect 40684 9662 40686 9714
rect 40686 9662 40738 9714
rect 40738 9662 40740 9714
rect 40684 9660 40740 9662
rect 39900 8428 39956 8484
rect 38780 6860 38836 6916
rect 38668 6018 38724 6020
rect 38668 5966 38670 6018
rect 38670 5966 38722 6018
rect 38722 5966 38724 6018
rect 38668 5964 38724 5966
rect 40236 8652 40292 8708
rect 40908 9266 40964 9268
rect 40908 9214 40910 9266
rect 40910 9214 40962 9266
rect 40962 9214 40964 9266
rect 40908 9212 40964 9214
rect 40796 8652 40852 8708
rect 41244 8988 41300 9044
rect 40236 7868 40292 7924
rect 41804 9772 41860 9828
rect 41692 9714 41748 9716
rect 41692 9662 41694 9714
rect 41694 9662 41746 9714
rect 41746 9662 41748 9714
rect 41692 9660 41748 9662
rect 41468 9602 41524 9604
rect 41468 9550 41470 9602
rect 41470 9550 41522 9602
rect 41522 9550 41524 9602
rect 41468 9548 41524 9550
rect 41804 8764 41860 8820
rect 41580 7980 41636 8036
rect 40908 7474 40964 7476
rect 40908 7422 40910 7474
rect 40910 7422 40962 7474
rect 40962 7422 40964 7474
rect 40908 7420 40964 7422
rect 40796 6466 40852 6468
rect 40796 6414 40798 6466
rect 40798 6414 40850 6466
rect 40850 6414 40852 6466
rect 40796 6412 40852 6414
rect 38556 5740 38612 5796
rect 39116 5740 39172 5796
rect 38780 5122 38836 5124
rect 38780 5070 38782 5122
rect 38782 5070 38834 5122
rect 38834 5070 38836 5122
rect 38780 5068 38836 5070
rect 38556 4844 38612 4900
rect 38892 4450 38948 4452
rect 38892 4398 38894 4450
rect 38894 4398 38946 4450
rect 38946 4398 38948 4450
rect 38892 4396 38948 4398
rect 39676 5628 39732 5684
rect 40236 5906 40292 5908
rect 40236 5854 40238 5906
rect 40238 5854 40290 5906
rect 40290 5854 40292 5906
rect 40236 5852 40292 5854
rect 41020 5794 41076 5796
rect 41020 5742 41022 5794
rect 41022 5742 41074 5794
rect 41074 5742 41076 5794
rect 41020 5740 41076 5742
rect 42140 9884 42196 9940
rect 42028 9212 42084 9268
rect 43484 13858 43540 13860
rect 43484 13806 43486 13858
rect 43486 13806 43538 13858
rect 43538 13806 43540 13858
rect 43484 13804 43540 13806
rect 43484 13580 43540 13636
rect 42924 12012 42980 12068
rect 44132 14138 44188 14140
rect 44132 14086 44134 14138
rect 44134 14086 44186 14138
rect 44186 14086 44188 14138
rect 44132 14084 44188 14086
rect 44236 14138 44292 14140
rect 44236 14086 44238 14138
rect 44238 14086 44290 14138
rect 44290 14086 44292 14138
rect 44236 14084 44292 14086
rect 44340 14138 44396 14140
rect 44340 14086 44342 14138
rect 44342 14086 44394 14138
rect 44394 14086 44396 14138
rect 44340 14084 44396 14086
rect 43932 13468 43988 13524
rect 43596 13244 43652 13300
rect 44716 17836 44772 17892
rect 44940 20188 44996 20244
rect 45164 19346 45220 19348
rect 45164 19294 45166 19346
rect 45166 19294 45218 19346
rect 45218 19294 45220 19346
rect 45164 19292 45220 19294
rect 45164 18338 45220 18340
rect 45164 18286 45166 18338
rect 45166 18286 45218 18338
rect 45218 18286 45220 18338
rect 45164 18284 45220 18286
rect 44604 15538 44660 15540
rect 44604 15486 44606 15538
rect 44606 15486 44658 15538
rect 44658 15486 44660 15538
rect 44604 15484 44660 15486
rect 45612 23212 45668 23268
rect 46508 23212 46564 23268
rect 45388 23154 45444 23156
rect 45388 23102 45390 23154
rect 45390 23102 45442 23154
rect 45442 23102 45444 23154
rect 45388 23100 45444 23102
rect 45500 22370 45556 22372
rect 45500 22318 45502 22370
rect 45502 22318 45554 22370
rect 45554 22318 45556 22370
rect 45500 22316 45556 22318
rect 45724 22316 45780 22372
rect 45388 20076 45444 20132
rect 45276 17164 45332 17220
rect 45164 16716 45220 16772
rect 44940 16604 44996 16660
rect 45276 16098 45332 16100
rect 45276 16046 45278 16098
rect 45278 16046 45330 16098
rect 45330 16046 45332 16098
rect 45276 16044 45332 16046
rect 45836 22258 45892 22260
rect 45836 22206 45838 22258
rect 45838 22206 45890 22258
rect 45890 22206 45892 22258
rect 45836 22204 45892 22206
rect 46396 22428 46452 22484
rect 46956 24668 47012 24724
rect 48188 26962 48244 26964
rect 48188 26910 48190 26962
rect 48190 26910 48242 26962
rect 48242 26910 48244 26962
rect 48188 26908 48244 26910
rect 48412 27132 48468 27188
rect 49308 30882 49364 30884
rect 49308 30830 49310 30882
rect 49310 30830 49362 30882
rect 49362 30830 49364 30882
rect 49308 30828 49364 30830
rect 49196 30156 49252 30212
rect 49196 29148 49252 29204
rect 49308 28140 49364 28196
rect 51324 33234 51380 33236
rect 51324 33182 51326 33234
rect 51326 33182 51378 33234
rect 51378 33182 51380 33234
rect 51324 33180 51380 33182
rect 50876 31948 50932 32004
rect 50764 30770 50820 30772
rect 50764 30718 50766 30770
rect 50766 30718 50818 30770
rect 50818 30718 50820 30770
rect 50764 30716 50820 30718
rect 50652 30380 50708 30436
rect 50428 30210 50484 30212
rect 50428 30158 50430 30210
rect 50430 30158 50482 30210
rect 50482 30158 50484 30210
rect 50428 30156 50484 30158
rect 50316 29260 50372 29316
rect 49532 29148 49588 29204
rect 47964 26178 48020 26180
rect 47964 26126 47966 26178
rect 47966 26126 48018 26178
rect 48018 26126 48020 26178
rect 47964 26124 48020 26126
rect 49308 27020 49364 27076
rect 49980 28812 50036 28868
rect 50540 27916 50596 27972
rect 50316 27858 50372 27860
rect 50316 27806 50318 27858
rect 50318 27806 50370 27858
rect 50370 27806 50372 27858
rect 50316 27804 50372 27806
rect 50764 27804 50820 27860
rect 50204 27580 50260 27636
rect 50876 27580 50932 27636
rect 49644 27020 49700 27076
rect 47852 25452 47908 25508
rect 46844 23714 46900 23716
rect 46844 23662 46846 23714
rect 46846 23662 46898 23714
rect 46898 23662 46900 23714
rect 46844 23660 46900 23662
rect 46956 23042 47012 23044
rect 46956 22990 46958 23042
rect 46958 22990 47010 23042
rect 47010 22990 47012 23042
rect 46956 22988 47012 22990
rect 46620 22204 46676 22260
rect 46732 22764 46788 22820
rect 47628 24610 47684 24612
rect 47628 24558 47630 24610
rect 47630 24558 47682 24610
rect 47682 24558 47684 24610
rect 47628 24556 47684 24558
rect 47404 23772 47460 23828
rect 47628 24108 47684 24164
rect 48188 25676 48244 25732
rect 48636 25506 48692 25508
rect 48636 25454 48638 25506
rect 48638 25454 48690 25506
rect 48690 25454 48692 25506
rect 48636 25452 48692 25454
rect 48188 24892 48244 24948
rect 49532 26908 49588 26964
rect 49308 26572 49364 26628
rect 48636 24108 48692 24164
rect 47180 23212 47236 23268
rect 46172 21810 46228 21812
rect 46172 21758 46174 21810
rect 46174 21758 46226 21810
rect 46226 21758 46228 21810
rect 46172 21756 46228 21758
rect 46060 21644 46116 21700
rect 45948 21308 46004 21364
rect 45948 21084 46004 21140
rect 46060 20636 46116 20692
rect 46172 20524 46228 20580
rect 46396 21644 46452 21700
rect 46844 21362 46900 21364
rect 46844 21310 46846 21362
rect 46846 21310 46898 21362
rect 46898 21310 46900 21362
rect 46844 21308 46900 21310
rect 46732 21196 46788 21252
rect 47180 22092 47236 22148
rect 47404 22988 47460 23044
rect 47404 22428 47460 22484
rect 47404 22258 47460 22260
rect 47404 22206 47406 22258
rect 47406 22206 47458 22258
rect 47458 22206 47460 22258
rect 47404 22204 47460 22206
rect 47964 23660 48020 23716
rect 48188 23212 48244 23268
rect 48300 23660 48356 23716
rect 48076 23154 48132 23156
rect 48076 23102 48078 23154
rect 48078 23102 48130 23154
rect 48130 23102 48132 23154
rect 48076 23100 48132 23102
rect 48188 23042 48244 23044
rect 48188 22990 48190 23042
rect 48190 22990 48242 23042
rect 48242 22990 48244 23042
rect 48188 22988 48244 22990
rect 48524 22988 48580 23044
rect 48076 22652 48132 22708
rect 47852 22092 47908 22148
rect 47964 22204 48020 22260
rect 47068 21532 47124 21588
rect 47516 21698 47572 21700
rect 47516 21646 47518 21698
rect 47518 21646 47570 21698
rect 47570 21646 47572 21698
rect 47516 21644 47572 21646
rect 48076 21698 48132 21700
rect 48076 21646 48078 21698
rect 48078 21646 48130 21698
rect 48130 21646 48132 21698
rect 48076 21644 48132 21646
rect 47852 21420 47908 21476
rect 46620 20690 46676 20692
rect 46620 20638 46622 20690
rect 46622 20638 46674 20690
rect 46674 20638 46676 20690
rect 46620 20636 46676 20638
rect 46508 19964 46564 20020
rect 45724 19010 45780 19012
rect 45724 18958 45726 19010
rect 45726 18958 45778 19010
rect 45778 18958 45780 19010
rect 45724 18956 45780 18958
rect 45724 18060 45780 18116
rect 45724 16940 45780 16996
rect 45612 16604 45668 16660
rect 45500 15820 45556 15876
rect 45724 15932 45780 15988
rect 45164 15596 45220 15652
rect 44268 13244 44324 13300
rect 44940 13804 44996 13860
rect 44716 13020 44772 13076
rect 43820 12012 43876 12068
rect 43260 11228 43316 11284
rect 42812 10220 42868 10276
rect 42812 9996 42868 10052
rect 43036 9996 43092 10052
rect 42252 9436 42308 9492
rect 42476 9602 42532 9604
rect 42476 9550 42478 9602
rect 42478 9550 42530 9602
rect 42530 9550 42532 9602
rect 42476 9548 42532 9550
rect 42700 9602 42756 9604
rect 42700 9550 42702 9602
rect 42702 9550 42754 9602
rect 42754 9550 42756 9602
rect 42700 9548 42756 9550
rect 43148 9602 43204 9604
rect 43148 9550 43150 9602
rect 43150 9550 43202 9602
rect 43202 9550 43204 9602
rect 43148 9548 43204 9550
rect 42588 9100 42644 9156
rect 43036 9042 43092 9044
rect 43036 8990 43038 9042
rect 43038 8990 43090 9042
rect 43090 8990 43092 9042
rect 43036 8988 43092 8990
rect 42028 6860 42084 6916
rect 42364 7980 42420 8036
rect 42588 7644 42644 7700
rect 43036 8764 43092 8820
rect 42476 6748 42532 6804
rect 42140 6636 42196 6692
rect 41244 6018 41300 6020
rect 41244 5966 41246 6018
rect 41246 5966 41298 6018
rect 41298 5966 41300 6018
rect 41244 5964 41300 5966
rect 41692 6578 41748 6580
rect 41692 6526 41694 6578
rect 41694 6526 41746 6578
rect 41746 6526 41748 6578
rect 41692 6524 41748 6526
rect 42364 6524 42420 6580
rect 41692 5740 41748 5796
rect 41804 5180 41860 5236
rect 39900 4956 39956 5012
rect 40348 5068 40404 5124
rect 40684 5122 40740 5124
rect 40684 5070 40686 5122
rect 40686 5070 40738 5122
rect 40738 5070 40740 5122
rect 40684 5068 40740 5070
rect 41020 5010 41076 5012
rect 41020 4958 41022 5010
rect 41022 4958 41074 5010
rect 41074 4958 41076 5010
rect 41020 4956 41076 4958
rect 39228 4732 39284 4788
rect 40236 4844 40292 4900
rect 40124 4620 40180 4676
rect 41468 4620 41524 4676
rect 39340 4338 39396 4340
rect 39340 4286 39342 4338
rect 39342 4286 39394 4338
rect 39394 4286 39396 4338
rect 39340 4284 39396 4286
rect 40460 4338 40516 4340
rect 40460 4286 40462 4338
rect 40462 4286 40514 4338
rect 40514 4286 40516 4338
rect 40460 4284 40516 4286
rect 41132 4338 41188 4340
rect 41132 4286 41134 4338
rect 41134 4286 41186 4338
rect 41186 4286 41188 4338
rect 41132 4284 41188 4286
rect 40796 4172 40852 4228
rect 42476 5906 42532 5908
rect 42476 5854 42478 5906
rect 42478 5854 42530 5906
rect 42530 5854 42532 5906
rect 42476 5852 42532 5854
rect 42364 5068 42420 5124
rect 42700 4898 42756 4900
rect 42700 4846 42702 4898
rect 42702 4846 42754 4898
rect 42754 4846 42756 4898
rect 42700 4844 42756 4846
rect 43596 11676 43652 11732
rect 44132 12570 44188 12572
rect 44132 12518 44134 12570
rect 44134 12518 44186 12570
rect 44186 12518 44188 12570
rect 44132 12516 44188 12518
rect 44236 12570 44292 12572
rect 44236 12518 44238 12570
rect 44238 12518 44290 12570
rect 44290 12518 44292 12570
rect 44236 12516 44292 12518
rect 44340 12570 44396 12572
rect 44340 12518 44342 12570
rect 44342 12518 44394 12570
rect 44394 12518 44396 12570
rect 44340 12516 44396 12518
rect 44044 12402 44100 12404
rect 44044 12350 44046 12402
rect 44046 12350 44098 12402
rect 44098 12350 44100 12402
rect 44044 12348 44100 12350
rect 45724 15484 45780 15540
rect 46060 19906 46116 19908
rect 46060 19854 46062 19906
rect 46062 19854 46114 19906
rect 46114 19854 46116 19906
rect 46060 19852 46116 19854
rect 46060 18956 46116 19012
rect 45948 17666 46004 17668
rect 45948 17614 45950 17666
rect 45950 17614 46002 17666
rect 46002 17614 46004 17666
rect 45948 17612 46004 17614
rect 45948 17164 46004 17220
rect 46732 19068 46788 19124
rect 46956 19180 47012 19236
rect 46172 16940 46228 16996
rect 46172 16098 46228 16100
rect 46172 16046 46174 16098
rect 46174 16046 46226 16098
rect 46226 16046 46228 16098
rect 46172 16044 46228 16046
rect 46284 15986 46340 15988
rect 46284 15934 46286 15986
rect 46286 15934 46338 15986
rect 46338 15934 46340 15986
rect 46284 15932 46340 15934
rect 46060 15820 46116 15876
rect 46060 15314 46116 15316
rect 46060 15262 46062 15314
rect 46062 15262 46114 15314
rect 46114 15262 46116 15314
rect 46060 15260 46116 15262
rect 45500 14588 45556 14644
rect 45276 13804 45332 13860
rect 45612 13468 45668 13524
rect 45164 13020 45220 13076
rect 45052 12348 45108 12404
rect 44716 12290 44772 12292
rect 44716 12238 44718 12290
rect 44718 12238 44770 12290
rect 44770 12238 44772 12290
rect 44716 12236 44772 12238
rect 45164 12460 45220 12516
rect 44380 12012 44436 12068
rect 43932 11228 43988 11284
rect 45276 12124 45332 12180
rect 45388 12236 45444 12292
rect 45388 11900 45444 11956
rect 45164 11282 45220 11284
rect 45164 11230 45166 11282
rect 45166 11230 45218 11282
rect 45218 11230 45220 11282
rect 45164 11228 45220 11230
rect 44132 11002 44188 11004
rect 44132 10950 44134 11002
rect 44134 10950 44186 11002
rect 44186 10950 44188 11002
rect 44132 10948 44188 10950
rect 44236 11002 44292 11004
rect 44236 10950 44238 11002
rect 44238 10950 44290 11002
rect 44290 10950 44292 11002
rect 44236 10948 44292 10950
rect 44340 11002 44396 11004
rect 44340 10950 44342 11002
rect 44342 10950 44394 11002
rect 44394 10950 44396 11002
rect 44340 10948 44396 10950
rect 43596 10556 43652 10612
rect 43596 9884 43652 9940
rect 43484 9772 43540 9828
rect 43932 9772 43988 9828
rect 43708 9714 43764 9716
rect 43708 9662 43710 9714
rect 43710 9662 43762 9714
rect 43762 9662 43764 9714
rect 43708 9660 43764 9662
rect 43260 8652 43316 8708
rect 44268 9996 44324 10052
rect 43932 9436 43988 9492
rect 44132 9434 44188 9436
rect 44132 9382 44134 9434
rect 44134 9382 44186 9434
rect 44186 9382 44188 9434
rect 44132 9380 44188 9382
rect 44236 9434 44292 9436
rect 44236 9382 44238 9434
rect 44238 9382 44290 9434
rect 44290 9382 44292 9434
rect 44236 9380 44292 9382
rect 44340 9434 44396 9436
rect 44340 9382 44342 9434
rect 44342 9382 44394 9434
rect 44394 9382 44396 9434
rect 44340 9380 44396 9382
rect 43932 8988 43988 9044
rect 44044 8428 44100 8484
rect 44716 10610 44772 10612
rect 44716 10558 44718 10610
rect 44718 10558 44770 10610
rect 44770 10558 44772 10610
rect 44716 10556 44772 10558
rect 44716 10108 44772 10164
rect 45052 9996 45108 10052
rect 45276 9772 45332 9828
rect 45388 9660 45444 9716
rect 46844 18172 46900 18228
rect 46508 17052 46564 17108
rect 46508 16604 46564 16660
rect 46396 15484 46452 15540
rect 47628 21196 47684 21252
rect 47180 21084 47236 21140
rect 47852 20972 47908 21028
rect 48076 21420 48132 21476
rect 47628 20690 47684 20692
rect 47628 20638 47630 20690
rect 47630 20638 47682 20690
rect 47682 20638 47684 20690
rect 47628 20636 47684 20638
rect 47852 20130 47908 20132
rect 47852 20078 47854 20130
rect 47854 20078 47906 20130
rect 47906 20078 47908 20130
rect 47852 20076 47908 20078
rect 47404 19852 47460 19908
rect 47180 19516 47236 19572
rect 47404 19292 47460 19348
rect 47292 19122 47348 19124
rect 47292 19070 47294 19122
rect 47294 19070 47346 19122
rect 47346 19070 47348 19122
rect 47292 19068 47348 19070
rect 47852 19234 47908 19236
rect 47852 19182 47854 19234
rect 47854 19182 47906 19234
rect 47906 19182 47908 19234
rect 47852 19180 47908 19182
rect 48860 23042 48916 23044
rect 48860 22990 48862 23042
rect 48862 22990 48914 23042
rect 48914 22990 48916 23042
rect 48860 22988 48916 22990
rect 49308 26236 49364 26292
rect 49084 25676 49140 25732
rect 50540 26962 50596 26964
rect 50540 26910 50542 26962
rect 50542 26910 50594 26962
rect 50594 26910 50596 26962
rect 50540 26908 50596 26910
rect 50764 26796 50820 26852
rect 50428 26290 50484 26292
rect 50428 26238 50430 26290
rect 50430 26238 50482 26290
rect 50482 26238 50484 26290
rect 50428 26236 50484 26238
rect 50204 25900 50260 25956
rect 49196 25228 49252 25284
rect 49420 24780 49476 24836
rect 49084 24556 49140 24612
rect 49308 24108 49364 24164
rect 53340 34130 53396 34132
rect 53340 34078 53342 34130
rect 53342 34078 53394 34130
rect 53394 34078 53396 34130
rect 53340 34076 53396 34078
rect 53228 33516 53284 33572
rect 53116 33458 53172 33460
rect 53116 33406 53118 33458
rect 53118 33406 53170 33458
rect 53170 33406 53172 33458
rect 53116 33404 53172 33406
rect 52892 33180 52948 33236
rect 51772 33122 51828 33124
rect 51772 33070 51774 33122
rect 51774 33070 51826 33122
rect 51826 33070 51828 33122
rect 51772 33068 51828 33070
rect 51286 32170 51342 32172
rect 51286 32118 51288 32170
rect 51288 32118 51340 32170
rect 51340 32118 51342 32170
rect 51286 32116 51342 32118
rect 51390 32170 51446 32172
rect 51390 32118 51392 32170
rect 51392 32118 51444 32170
rect 51444 32118 51446 32170
rect 51390 32116 51446 32118
rect 51494 32170 51550 32172
rect 51494 32118 51496 32170
rect 51496 32118 51548 32170
rect 51548 32118 51550 32170
rect 51494 32116 51550 32118
rect 53116 32508 53172 32564
rect 51286 30602 51342 30604
rect 51286 30550 51288 30602
rect 51288 30550 51340 30602
rect 51340 30550 51342 30602
rect 51286 30548 51342 30550
rect 51390 30602 51446 30604
rect 51390 30550 51392 30602
rect 51392 30550 51444 30602
rect 51444 30550 51446 30602
rect 51390 30548 51446 30550
rect 51494 30602 51550 30604
rect 51494 30550 51496 30602
rect 51496 30550 51548 30602
rect 51548 30550 51550 30602
rect 51494 30548 51550 30550
rect 51212 29314 51268 29316
rect 51212 29262 51214 29314
rect 51214 29262 51266 29314
rect 51266 29262 51268 29314
rect 51212 29260 51268 29262
rect 51660 29484 51716 29540
rect 51772 29372 51828 29428
rect 51286 29034 51342 29036
rect 51286 28982 51288 29034
rect 51288 28982 51340 29034
rect 51340 28982 51342 29034
rect 51286 28980 51342 28982
rect 51390 29034 51446 29036
rect 51390 28982 51392 29034
rect 51392 28982 51444 29034
rect 51444 28982 51446 29034
rect 51390 28980 51446 28982
rect 51494 29034 51550 29036
rect 51494 28982 51496 29034
rect 51496 28982 51548 29034
rect 51548 28982 51550 29034
rect 51494 28980 51550 28982
rect 51548 28812 51604 28868
rect 51436 28642 51492 28644
rect 51436 28590 51438 28642
rect 51438 28590 51490 28642
rect 51490 28590 51492 28642
rect 51436 28588 51492 28590
rect 51436 27858 51492 27860
rect 51436 27806 51438 27858
rect 51438 27806 51490 27858
rect 51490 27806 51492 27858
rect 51436 27804 51492 27806
rect 51884 28700 51940 28756
rect 52780 29986 52836 29988
rect 52780 29934 52782 29986
rect 52782 29934 52834 29986
rect 52834 29934 52836 29986
rect 52780 29932 52836 29934
rect 53004 29932 53060 29988
rect 53004 29426 53060 29428
rect 53004 29374 53006 29426
rect 53006 29374 53058 29426
rect 53058 29374 53060 29426
rect 53004 29372 53060 29374
rect 52668 28812 52724 28868
rect 52780 28754 52836 28756
rect 52780 28702 52782 28754
rect 52782 28702 52834 28754
rect 52834 28702 52836 28754
rect 52780 28700 52836 28702
rect 52108 28530 52164 28532
rect 52108 28478 52110 28530
rect 52110 28478 52162 28530
rect 52162 28478 52164 28530
rect 52108 28476 52164 28478
rect 51772 28028 51828 28084
rect 51884 27970 51940 27972
rect 51884 27918 51886 27970
rect 51886 27918 51938 27970
rect 51938 27918 51940 27970
rect 51884 27916 51940 27918
rect 51286 27466 51342 27468
rect 51286 27414 51288 27466
rect 51288 27414 51340 27466
rect 51340 27414 51342 27466
rect 51286 27412 51342 27414
rect 51390 27466 51446 27468
rect 51390 27414 51392 27466
rect 51392 27414 51444 27466
rect 51444 27414 51446 27466
rect 51390 27412 51446 27414
rect 51494 27466 51550 27468
rect 51494 27414 51496 27466
rect 51496 27414 51548 27466
rect 51548 27414 51550 27466
rect 51494 27412 51550 27414
rect 51884 27244 51940 27300
rect 51884 26908 51940 26964
rect 51548 26796 51604 26852
rect 51660 26572 51716 26628
rect 52556 28140 52612 28196
rect 52108 27692 52164 27748
rect 52444 27580 52500 27636
rect 51884 26572 51940 26628
rect 53004 27858 53060 27860
rect 53004 27806 53006 27858
rect 53006 27806 53058 27858
rect 53058 27806 53060 27858
rect 53004 27804 53060 27806
rect 52892 27746 52948 27748
rect 52892 27694 52894 27746
rect 52894 27694 52946 27746
rect 52946 27694 52948 27746
rect 52892 27692 52948 27694
rect 52780 27298 52836 27300
rect 52780 27246 52782 27298
rect 52782 27246 52834 27298
rect 52834 27246 52836 27298
rect 52780 27244 52836 27246
rect 52556 27020 52612 27076
rect 51286 25898 51342 25900
rect 51286 25846 51288 25898
rect 51288 25846 51340 25898
rect 51340 25846 51342 25898
rect 51286 25844 51342 25846
rect 51390 25898 51446 25900
rect 51390 25846 51392 25898
rect 51392 25846 51444 25898
rect 51444 25846 51446 25898
rect 51390 25844 51446 25846
rect 51494 25898 51550 25900
rect 51494 25846 51496 25898
rect 51496 25846 51548 25898
rect 51548 25846 51550 25898
rect 51494 25844 51550 25846
rect 51212 25676 51268 25732
rect 51548 25564 51604 25620
rect 52220 26124 52276 26180
rect 51772 25676 51828 25732
rect 50428 24892 50484 24948
rect 50540 24834 50596 24836
rect 50540 24782 50542 24834
rect 50542 24782 50594 24834
rect 50594 24782 50596 24834
rect 50540 24780 50596 24782
rect 50428 24722 50484 24724
rect 50428 24670 50430 24722
rect 50430 24670 50482 24722
rect 50482 24670 50484 24722
rect 50428 24668 50484 24670
rect 49756 24220 49812 24276
rect 49308 23324 49364 23380
rect 49084 23212 49140 23268
rect 48972 22764 49028 22820
rect 48412 22428 48468 22484
rect 48972 22316 49028 22372
rect 48300 21586 48356 21588
rect 48300 21534 48302 21586
rect 48302 21534 48354 21586
rect 48354 21534 48356 21586
rect 48300 21532 48356 21534
rect 48412 21308 48468 21364
rect 48076 20018 48132 20020
rect 48076 19966 48078 20018
rect 48078 19966 48130 20018
rect 48130 19966 48132 20018
rect 48076 19964 48132 19966
rect 47180 18396 47236 18452
rect 47516 17948 47572 18004
rect 46732 16940 46788 16996
rect 46956 17052 47012 17108
rect 47292 16994 47348 16996
rect 47292 16942 47294 16994
rect 47294 16942 47346 16994
rect 47346 16942 47348 16994
rect 47292 16940 47348 16942
rect 46844 16828 46900 16884
rect 46956 16716 47012 16772
rect 46620 15372 46676 15428
rect 46956 16380 47012 16436
rect 47068 16156 47124 16212
rect 47852 18844 47908 18900
rect 47964 18732 48020 18788
rect 48188 19234 48244 19236
rect 48188 19182 48190 19234
rect 48190 19182 48242 19234
rect 48242 19182 48244 19234
rect 48188 19180 48244 19182
rect 48188 18732 48244 18788
rect 48188 18508 48244 18564
rect 47964 18396 48020 18452
rect 47852 17554 47908 17556
rect 47852 17502 47854 17554
rect 47854 17502 47906 17554
rect 47906 17502 47908 17554
rect 47852 17500 47908 17502
rect 49308 22258 49364 22260
rect 49308 22206 49310 22258
rect 49310 22206 49362 22258
rect 49362 22206 49364 22258
rect 49308 22204 49364 22206
rect 50428 23996 50484 24052
rect 49868 23714 49924 23716
rect 49868 23662 49870 23714
rect 49870 23662 49922 23714
rect 49922 23662 49924 23714
rect 49868 23660 49924 23662
rect 50092 23714 50148 23716
rect 50092 23662 50094 23714
rect 50094 23662 50146 23714
rect 50146 23662 50148 23714
rect 50092 23660 50148 23662
rect 49756 23548 49812 23604
rect 49644 23212 49700 23268
rect 49756 23042 49812 23044
rect 49756 22990 49758 23042
rect 49758 22990 49810 23042
rect 49810 22990 49812 23042
rect 49756 22988 49812 22990
rect 50204 23378 50260 23380
rect 50204 23326 50206 23378
rect 50206 23326 50258 23378
rect 50258 23326 50260 23378
rect 50204 23324 50260 23326
rect 51548 24892 51604 24948
rect 51286 24330 51342 24332
rect 51286 24278 51288 24330
rect 51288 24278 51340 24330
rect 51340 24278 51342 24330
rect 51286 24276 51342 24278
rect 51390 24330 51446 24332
rect 51390 24278 51392 24330
rect 51392 24278 51444 24330
rect 51444 24278 51446 24330
rect 51390 24276 51446 24278
rect 51494 24330 51550 24332
rect 51494 24278 51496 24330
rect 51496 24278 51548 24330
rect 51548 24278 51550 24330
rect 51494 24276 51550 24278
rect 50540 23714 50596 23716
rect 50540 23662 50542 23714
rect 50542 23662 50594 23714
rect 50594 23662 50596 23714
rect 50540 23660 50596 23662
rect 50764 23714 50820 23716
rect 50764 23662 50766 23714
rect 50766 23662 50818 23714
rect 50818 23662 50820 23714
rect 50764 23660 50820 23662
rect 50652 23266 50708 23268
rect 50652 23214 50654 23266
rect 50654 23214 50706 23266
rect 50706 23214 50708 23266
rect 50652 23212 50708 23214
rect 50428 22652 50484 22708
rect 49756 21644 49812 21700
rect 48972 20860 49028 20916
rect 49196 20412 49252 20468
rect 48748 19628 48804 19684
rect 48860 20300 48916 20356
rect 49420 20188 49476 20244
rect 48636 19068 48692 19124
rect 48972 20018 49028 20020
rect 48972 19966 48974 20018
rect 48974 19966 49026 20018
rect 49026 19966 49028 20018
rect 48972 19964 49028 19966
rect 48972 19404 49028 19460
rect 49644 20076 49700 20132
rect 49756 20018 49812 20020
rect 49756 19966 49758 20018
rect 49758 19966 49810 20018
rect 49810 19966 49812 20018
rect 49756 19964 49812 19966
rect 50428 22204 50484 22260
rect 50204 22146 50260 22148
rect 50204 22094 50206 22146
rect 50206 22094 50258 22146
rect 50258 22094 50260 22146
rect 50204 22092 50260 22094
rect 50092 21196 50148 21252
rect 50316 21980 50372 22036
rect 49532 19516 49588 19572
rect 50204 20412 50260 20468
rect 51324 23772 51380 23828
rect 51324 23548 51380 23604
rect 51548 23660 51604 23716
rect 51286 22762 51342 22764
rect 51286 22710 51288 22762
rect 51288 22710 51340 22762
rect 51340 22710 51342 22762
rect 51286 22708 51342 22710
rect 51390 22762 51446 22764
rect 51390 22710 51392 22762
rect 51392 22710 51444 22762
rect 51444 22710 51446 22762
rect 51390 22708 51446 22710
rect 51494 22762 51550 22764
rect 51494 22710 51496 22762
rect 51496 22710 51548 22762
rect 51548 22710 51550 22762
rect 51494 22708 51550 22710
rect 52108 25282 52164 25284
rect 52108 25230 52110 25282
rect 52110 25230 52162 25282
rect 52162 25230 52164 25282
rect 52108 25228 52164 25230
rect 52780 25676 52836 25732
rect 52892 25564 52948 25620
rect 53340 32002 53396 32004
rect 53340 31950 53342 32002
rect 53342 31950 53394 32002
rect 53394 31950 53396 32002
rect 53340 31948 53396 31950
rect 56028 36258 56084 36260
rect 56028 36206 56030 36258
rect 56030 36206 56082 36258
rect 56082 36206 56084 36258
rect 56028 36204 56084 36206
rect 55580 35810 55636 35812
rect 55580 35758 55582 35810
rect 55582 35758 55634 35810
rect 55634 35758 55636 35810
rect 55580 35756 55636 35758
rect 55244 35698 55300 35700
rect 55244 35646 55246 35698
rect 55246 35646 55298 35698
rect 55298 35646 55300 35698
rect 55244 35644 55300 35646
rect 55692 35532 55748 35588
rect 55356 35420 55412 35476
rect 55356 34860 55412 34916
rect 55132 34636 55188 34692
rect 54572 34130 54628 34132
rect 54572 34078 54574 34130
rect 54574 34078 54626 34130
rect 54626 34078 54628 34130
rect 54572 34076 54628 34078
rect 55468 34076 55524 34132
rect 55692 34860 55748 34916
rect 54460 33570 54516 33572
rect 54460 33518 54462 33570
rect 54462 33518 54514 33570
rect 54514 33518 54516 33570
rect 54460 33516 54516 33518
rect 56140 35196 56196 35252
rect 56364 37100 56420 37156
rect 56476 36370 56532 36372
rect 56476 36318 56478 36370
rect 56478 36318 56530 36370
rect 56530 36318 56532 36370
rect 56476 36316 56532 36318
rect 56924 36594 56980 36596
rect 56924 36542 56926 36594
rect 56926 36542 56978 36594
rect 56978 36542 56980 36594
rect 56924 36540 56980 36542
rect 58439 36090 58495 36092
rect 58439 36038 58441 36090
rect 58441 36038 58493 36090
rect 58493 36038 58495 36090
rect 58439 36036 58495 36038
rect 58543 36090 58599 36092
rect 58543 36038 58545 36090
rect 58545 36038 58597 36090
rect 58597 36038 58599 36090
rect 58543 36036 58599 36038
rect 58647 36090 58703 36092
rect 58647 36038 58649 36090
rect 58649 36038 58701 36090
rect 58701 36038 58703 36090
rect 58647 36036 58703 36038
rect 56476 35698 56532 35700
rect 56476 35646 56478 35698
rect 56478 35646 56530 35698
rect 56530 35646 56532 35698
rect 56476 35644 56532 35646
rect 56252 34972 56308 35028
rect 55916 34076 55972 34132
rect 54236 32562 54292 32564
rect 54236 32510 54238 32562
rect 54238 32510 54290 32562
rect 54290 32510 54292 32562
rect 54236 32508 54292 32510
rect 54012 32284 54068 32340
rect 55132 32396 55188 32452
rect 53564 31778 53620 31780
rect 53564 31726 53566 31778
rect 53566 31726 53618 31778
rect 53618 31726 53620 31778
rect 53564 31724 53620 31726
rect 53676 30380 53732 30436
rect 53788 30156 53844 30212
rect 53228 29372 53284 29428
rect 53340 29260 53396 29316
rect 54908 31836 54964 31892
rect 54460 30828 54516 30884
rect 54460 30322 54516 30324
rect 54460 30270 54462 30322
rect 54462 30270 54514 30322
rect 54514 30270 54516 30322
rect 54460 30268 54516 30270
rect 54012 29148 54068 29204
rect 54124 30098 54180 30100
rect 54124 30046 54126 30098
rect 54126 30046 54178 30098
rect 54178 30046 54180 30098
rect 54124 30044 54180 30046
rect 53788 29036 53844 29092
rect 53228 28642 53284 28644
rect 53228 28590 53230 28642
rect 53230 28590 53282 28642
rect 53282 28590 53284 28642
rect 53228 28588 53284 28590
rect 54236 29932 54292 29988
rect 54348 29538 54404 29540
rect 54348 29486 54350 29538
rect 54350 29486 54402 29538
rect 54402 29486 54404 29538
rect 54348 29484 54404 29486
rect 54572 29426 54628 29428
rect 54572 29374 54574 29426
rect 54574 29374 54626 29426
rect 54626 29374 54628 29426
rect 54572 29372 54628 29374
rect 54236 29036 54292 29092
rect 55916 32674 55972 32676
rect 55916 32622 55918 32674
rect 55918 32622 55970 32674
rect 55970 32622 55972 32674
rect 55916 32620 55972 32622
rect 56588 35084 56644 35140
rect 56700 35196 56756 35252
rect 56588 34748 56644 34804
rect 56700 34130 56756 34132
rect 56700 34078 56702 34130
rect 56702 34078 56754 34130
rect 56754 34078 56756 34130
rect 56700 34076 56756 34078
rect 55468 31836 55524 31892
rect 57148 32450 57204 32452
rect 57148 32398 57150 32450
rect 57150 32398 57202 32450
rect 57202 32398 57204 32450
rect 57148 32396 57204 32398
rect 56588 31724 56644 31780
rect 55244 30828 55300 30884
rect 56924 31778 56980 31780
rect 56924 31726 56926 31778
rect 56926 31726 56978 31778
rect 56978 31726 56980 31778
rect 56924 31724 56980 31726
rect 55692 30210 55748 30212
rect 55692 30158 55694 30210
rect 55694 30158 55746 30210
rect 55746 30158 55748 30210
rect 55692 30156 55748 30158
rect 55468 30044 55524 30100
rect 55804 30044 55860 30100
rect 56700 30268 56756 30324
rect 57148 30322 57204 30324
rect 57148 30270 57150 30322
rect 57150 30270 57202 30322
rect 57202 30270 57204 30322
rect 57148 30268 57204 30270
rect 56140 29596 56196 29652
rect 56924 29596 56980 29652
rect 54796 29260 54852 29316
rect 54684 28812 54740 28868
rect 55692 28866 55748 28868
rect 55692 28814 55694 28866
rect 55694 28814 55746 28866
rect 55746 28814 55748 28866
rect 55692 28812 55748 28814
rect 54012 28700 54068 28756
rect 53788 28588 53844 28644
rect 54348 28476 54404 28532
rect 54236 28082 54292 28084
rect 54236 28030 54238 28082
rect 54238 28030 54290 28082
rect 54290 28030 54292 28082
rect 54236 28028 54292 28030
rect 55020 28642 55076 28644
rect 55020 28590 55022 28642
rect 55022 28590 55074 28642
rect 55074 28590 55076 28642
rect 55020 28588 55076 28590
rect 55916 29538 55972 29540
rect 55916 29486 55918 29538
rect 55918 29486 55970 29538
rect 55970 29486 55972 29538
rect 55916 29484 55972 29486
rect 55804 28588 55860 28644
rect 55916 29148 55972 29204
rect 53788 27692 53844 27748
rect 54572 27692 54628 27748
rect 53340 26348 53396 26404
rect 53452 26572 53508 26628
rect 53228 26124 53284 26180
rect 53340 25452 53396 25508
rect 53900 26796 53956 26852
rect 53452 25340 53508 25396
rect 51996 24162 52052 24164
rect 51996 24110 51998 24162
rect 51998 24110 52050 24162
rect 52050 24110 52052 24162
rect 51996 24108 52052 24110
rect 51996 22204 52052 22260
rect 50876 21868 50932 21924
rect 50988 21756 51044 21812
rect 50652 21698 50708 21700
rect 50652 21646 50654 21698
rect 50654 21646 50706 21698
rect 50706 21646 50708 21698
rect 50652 21644 50708 21646
rect 51100 21532 51156 21588
rect 50428 20748 50484 20804
rect 50428 20412 50484 20468
rect 50652 21196 50708 21252
rect 50316 20300 50372 20356
rect 50652 20802 50708 20804
rect 50652 20750 50654 20802
rect 50654 20750 50706 20802
rect 50706 20750 50708 20802
rect 50652 20748 50708 20750
rect 50876 20860 50932 20916
rect 51324 22146 51380 22148
rect 51324 22094 51326 22146
rect 51326 22094 51378 22146
rect 51378 22094 51380 22146
rect 51324 22092 51380 22094
rect 51324 21868 51380 21924
rect 50876 20412 50932 20468
rect 50316 20130 50372 20132
rect 50316 20078 50318 20130
rect 50318 20078 50370 20130
rect 50370 20078 50372 20130
rect 50316 20076 50372 20078
rect 49420 19068 49476 19124
rect 48860 18956 48916 19012
rect 49084 18844 49140 18900
rect 47964 17276 48020 17332
rect 47740 17164 47796 17220
rect 47852 16940 47908 16996
rect 47628 16882 47684 16884
rect 47628 16830 47630 16882
rect 47630 16830 47682 16882
rect 47682 16830 47684 16882
rect 47628 16828 47684 16830
rect 47516 16716 47572 16772
rect 46956 15484 47012 15540
rect 47516 15820 47572 15876
rect 46732 15260 46788 15316
rect 47292 15260 47348 15316
rect 46172 14530 46228 14532
rect 46172 14478 46174 14530
rect 46174 14478 46226 14530
rect 46226 14478 46228 14530
rect 46172 14476 46228 14478
rect 46620 14588 46676 14644
rect 46060 12908 46116 12964
rect 46284 13356 46340 13412
rect 46396 12908 46452 12964
rect 46172 12796 46228 12852
rect 45612 12236 45668 12292
rect 45836 12178 45892 12180
rect 45836 12126 45838 12178
rect 45838 12126 45890 12178
rect 45890 12126 45892 12178
rect 45836 12124 45892 12126
rect 45612 11900 45668 11956
rect 45836 11900 45892 11956
rect 46396 12178 46452 12180
rect 46396 12126 46398 12178
rect 46398 12126 46450 12178
rect 46450 12126 46452 12178
rect 46396 12124 46452 12126
rect 46956 15090 47012 15092
rect 46956 15038 46958 15090
rect 46958 15038 47010 15090
rect 47010 15038 47012 15090
rect 46956 15036 47012 15038
rect 46956 14588 47012 14644
rect 47292 13858 47348 13860
rect 47292 13806 47294 13858
rect 47294 13806 47346 13858
rect 47346 13806 47348 13858
rect 47292 13804 47348 13806
rect 46844 12962 46900 12964
rect 46844 12910 46846 12962
rect 46846 12910 46898 12962
rect 46898 12910 46900 12962
rect 46844 12908 46900 12910
rect 46844 12236 46900 12292
rect 46172 12012 46228 12068
rect 45724 11676 45780 11732
rect 46060 11788 46116 11844
rect 45724 11228 45780 11284
rect 45612 9714 45668 9716
rect 45612 9662 45614 9714
rect 45614 9662 45666 9714
rect 45666 9662 45668 9714
rect 45612 9660 45668 9662
rect 45948 11340 46004 11396
rect 45948 9996 46004 10052
rect 45948 9826 46004 9828
rect 45948 9774 45950 9826
rect 45950 9774 46002 9826
rect 46002 9774 46004 9826
rect 45948 9772 46004 9774
rect 46508 11900 46564 11956
rect 46284 11676 46340 11732
rect 46620 11788 46676 11844
rect 46396 11228 46452 11284
rect 47180 12402 47236 12404
rect 47180 12350 47182 12402
rect 47182 12350 47234 12402
rect 47234 12350 47236 12402
rect 47180 12348 47236 12350
rect 47068 12012 47124 12068
rect 48412 16210 48468 16212
rect 48412 16158 48414 16210
rect 48414 16158 48466 16210
rect 48466 16158 48468 16210
rect 48412 16156 48468 16158
rect 48188 16098 48244 16100
rect 48188 16046 48190 16098
rect 48190 16046 48242 16098
rect 48242 16046 48244 16098
rect 48188 16044 48244 16046
rect 47964 15986 48020 15988
rect 47964 15934 47966 15986
rect 47966 15934 48018 15986
rect 48018 15934 48020 15986
rect 47964 15932 48020 15934
rect 48188 15426 48244 15428
rect 48188 15374 48190 15426
rect 48190 15374 48242 15426
rect 48242 15374 48244 15426
rect 48188 15372 48244 15374
rect 48748 17500 48804 17556
rect 49308 18172 49364 18228
rect 48748 16716 48804 16772
rect 48636 16098 48692 16100
rect 48636 16046 48638 16098
rect 48638 16046 48690 16098
rect 48690 16046 48692 16098
rect 48636 16044 48692 16046
rect 48076 14476 48132 14532
rect 47516 13580 47572 13636
rect 47852 13244 47908 13300
rect 48300 14418 48356 14420
rect 48300 14366 48302 14418
rect 48302 14366 48354 14418
rect 48354 14366 48356 14418
rect 48300 14364 48356 14366
rect 48188 14306 48244 14308
rect 48188 14254 48190 14306
rect 48190 14254 48242 14306
rect 48242 14254 48244 14306
rect 48188 14252 48244 14254
rect 48300 13580 48356 13636
rect 48188 13356 48244 13412
rect 48300 13020 48356 13076
rect 47404 12012 47460 12068
rect 47180 11954 47236 11956
rect 47180 11902 47182 11954
rect 47182 11902 47234 11954
rect 47234 11902 47236 11954
rect 47180 11900 47236 11902
rect 46956 11452 47012 11508
rect 47964 11506 48020 11508
rect 47964 11454 47966 11506
rect 47966 11454 48018 11506
rect 48018 11454 48020 11506
rect 47964 11452 48020 11454
rect 48188 11394 48244 11396
rect 48188 11342 48190 11394
rect 48190 11342 48242 11394
rect 48242 11342 48244 11394
rect 48188 11340 48244 11342
rect 45500 9042 45556 9044
rect 45500 8990 45502 9042
rect 45502 8990 45554 9042
rect 45554 8990 45556 9042
rect 45500 8988 45556 8990
rect 45388 8930 45444 8932
rect 45388 8878 45390 8930
rect 45390 8878 45442 8930
rect 45442 8878 45444 8930
rect 45388 8876 45444 8878
rect 44604 8428 44660 8484
rect 45388 8652 45444 8708
rect 46060 9212 46116 9268
rect 46284 8764 46340 8820
rect 46620 9996 46676 10052
rect 46620 9826 46676 9828
rect 46620 9774 46622 9826
rect 46622 9774 46674 9826
rect 46674 9774 46676 9826
rect 46620 9772 46676 9774
rect 46956 9996 47012 10052
rect 46956 9548 47012 9604
rect 47068 8764 47124 8820
rect 45612 8316 45668 8372
rect 46396 8316 46452 8372
rect 43932 8146 43988 8148
rect 43932 8094 43934 8146
rect 43934 8094 43986 8146
rect 43986 8094 43988 8146
rect 43932 8092 43988 8094
rect 43708 7980 43764 8036
rect 44716 7980 44772 8036
rect 44132 7866 44188 7868
rect 44132 7814 44134 7866
rect 44134 7814 44186 7866
rect 44186 7814 44188 7866
rect 44132 7812 44188 7814
rect 44236 7866 44292 7868
rect 44236 7814 44238 7866
rect 44238 7814 44290 7866
rect 44290 7814 44292 7866
rect 44236 7812 44292 7814
rect 44340 7866 44396 7868
rect 44340 7814 44342 7866
rect 44342 7814 44394 7866
rect 44394 7814 44396 7866
rect 44340 7812 44396 7814
rect 43484 7474 43540 7476
rect 43484 7422 43486 7474
rect 43486 7422 43538 7474
rect 43538 7422 43540 7474
rect 43484 7420 43540 7422
rect 43372 7308 43428 7364
rect 43260 6636 43316 6692
rect 44604 7474 44660 7476
rect 44604 7422 44606 7474
rect 44606 7422 44658 7474
rect 44658 7422 44660 7474
rect 44604 7420 44660 7422
rect 44940 8034 44996 8036
rect 44940 7982 44942 8034
rect 44942 7982 44994 8034
rect 44994 7982 44996 8034
rect 44940 7980 44996 7982
rect 44828 7868 44884 7924
rect 44828 7698 44884 7700
rect 44828 7646 44830 7698
rect 44830 7646 44882 7698
rect 44882 7646 44884 7698
rect 44828 7644 44884 7646
rect 46060 8258 46116 8260
rect 46060 8206 46062 8258
rect 46062 8206 46114 8258
rect 46114 8206 46116 8258
rect 46060 8204 46116 8206
rect 45724 7420 45780 7476
rect 46172 8092 46228 8148
rect 46620 8034 46676 8036
rect 46620 7982 46622 8034
rect 46622 7982 46674 8034
rect 46674 7982 46676 8034
rect 46620 7980 46676 7982
rect 46396 7474 46452 7476
rect 46396 7422 46398 7474
rect 46398 7422 46450 7474
rect 46450 7422 46452 7474
rect 46396 7420 46452 7422
rect 44380 6972 44436 7028
rect 45724 6972 45780 7028
rect 44156 6748 44212 6804
rect 44044 6690 44100 6692
rect 44044 6638 44046 6690
rect 44046 6638 44098 6690
rect 44098 6638 44100 6690
rect 44044 6636 44100 6638
rect 43484 5234 43540 5236
rect 43484 5182 43486 5234
rect 43486 5182 43538 5234
rect 43538 5182 43540 5234
rect 43484 5180 43540 5182
rect 45948 6802 46004 6804
rect 45948 6750 45950 6802
rect 45950 6750 46002 6802
rect 46002 6750 46004 6802
rect 45948 6748 46004 6750
rect 44132 6298 44188 6300
rect 44132 6246 44134 6298
rect 44134 6246 44186 6298
rect 44186 6246 44188 6298
rect 44132 6244 44188 6246
rect 44236 6298 44292 6300
rect 44236 6246 44238 6298
rect 44238 6246 44290 6298
rect 44290 6246 44292 6298
rect 44236 6244 44292 6246
rect 44340 6298 44396 6300
rect 44340 6246 44342 6298
rect 44342 6246 44394 6298
rect 44394 6246 44396 6298
rect 44340 6244 44396 6246
rect 44268 5292 44324 5348
rect 43708 5234 43764 5236
rect 43708 5182 43710 5234
rect 43710 5182 43762 5234
rect 43762 5182 43764 5234
rect 43708 5180 43764 5182
rect 46284 6636 46340 6692
rect 46508 7308 46564 7364
rect 46732 7308 46788 7364
rect 45388 5292 45444 5348
rect 44828 5180 44884 5236
rect 44716 4844 44772 4900
rect 43708 4732 43764 4788
rect 42812 4620 42868 4676
rect 43596 4620 43652 4676
rect 43260 4450 43316 4452
rect 43260 4398 43262 4450
rect 43262 4398 43314 4450
rect 43314 4398 43316 4450
rect 43260 4396 43316 4398
rect 42140 4284 42196 4340
rect 42476 4172 42532 4228
rect 43820 4172 43876 4228
rect 44132 4730 44188 4732
rect 44132 4678 44134 4730
rect 44134 4678 44186 4730
rect 44186 4678 44188 4730
rect 44132 4676 44188 4678
rect 44236 4730 44292 4732
rect 44236 4678 44238 4730
rect 44238 4678 44290 4730
rect 44290 4678 44292 4730
rect 44236 4676 44292 4678
rect 44340 4730 44396 4732
rect 44340 4678 44342 4730
rect 44342 4678 44394 4730
rect 44394 4678 44396 4730
rect 44340 4676 44396 4678
rect 44604 3724 44660 3780
rect 45724 4172 45780 4228
rect 45052 3330 45108 3332
rect 45052 3278 45054 3330
rect 45054 3278 45106 3330
rect 45106 3278 45108 3330
rect 45052 3276 45108 3278
rect 44132 3162 44188 3164
rect 44132 3110 44134 3162
rect 44134 3110 44186 3162
rect 44186 3110 44188 3162
rect 44132 3108 44188 3110
rect 44236 3162 44292 3164
rect 44236 3110 44238 3162
rect 44238 3110 44290 3162
rect 44290 3110 44292 3162
rect 44236 3108 44292 3110
rect 44340 3162 44396 3164
rect 44340 3110 44342 3162
rect 44342 3110 44394 3162
rect 44394 3110 44396 3162
rect 44340 3108 44396 3110
rect 47404 9660 47460 9716
rect 47404 8988 47460 9044
rect 47292 8370 47348 8372
rect 47292 8318 47294 8370
rect 47294 8318 47346 8370
rect 47346 8318 47348 8370
rect 47292 8316 47348 8318
rect 47068 8258 47124 8260
rect 47068 8206 47070 8258
rect 47070 8206 47122 8258
rect 47122 8206 47124 8258
rect 47068 8204 47124 8206
rect 47516 8146 47572 8148
rect 47516 8094 47518 8146
rect 47518 8094 47570 8146
rect 47570 8094 47572 8146
rect 47516 8092 47572 8094
rect 46956 7586 47012 7588
rect 46956 7534 46958 7586
rect 46958 7534 47010 7586
rect 47010 7534 47012 7586
rect 46956 7532 47012 7534
rect 47628 7532 47684 7588
rect 48188 9548 48244 9604
rect 48636 15036 48692 15092
rect 49084 17554 49140 17556
rect 49084 17502 49086 17554
rect 49086 17502 49138 17554
rect 49138 17502 49140 17554
rect 49084 17500 49140 17502
rect 48972 17388 49028 17444
rect 48860 16380 48916 16436
rect 48860 16156 48916 16212
rect 49308 16210 49364 16212
rect 49308 16158 49310 16210
rect 49310 16158 49362 16210
rect 49362 16158 49364 16210
rect 49308 16156 49364 16158
rect 49196 15932 49252 15988
rect 49084 15260 49140 15316
rect 48748 14530 48804 14532
rect 48748 14478 48750 14530
rect 48750 14478 48802 14530
rect 48802 14478 48804 14530
rect 48748 14476 48804 14478
rect 48860 14364 48916 14420
rect 48860 13244 48916 13300
rect 48748 11564 48804 11620
rect 48524 9826 48580 9828
rect 48524 9774 48526 9826
rect 48526 9774 48578 9826
rect 48578 9774 48580 9826
rect 48524 9772 48580 9774
rect 48524 8876 48580 8932
rect 48076 8092 48132 8148
rect 48076 7474 48132 7476
rect 48076 7422 48078 7474
rect 48078 7422 48130 7474
rect 48130 7422 48132 7474
rect 48076 7420 48132 7422
rect 46844 6972 46900 7028
rect 46620 4396 46676 4452
rect 45948 3724 46004 3780
rect 47740 6690 47796 6692
rect 47740 6638 47742 6690
rect 47742 6638 47794 6690
rect 47794 6638 47796 6690
rect 47740 6636 47796 6638
rect 48188 7196 48244 7252
rect 47180 5906 47236 5908
rect 47180 5854 47182 5906
rect 47182 5854 47234 5906
rect 47234 5854 47236 5906
rect 47180 5852 47236 5854
rect 47628 5906 47684 5908
rect 47628 5854 47630 5906
rect 47630 5854 47682 5906
rect 47682 5854 47684 5906
rect 47628 5852 47684 5854
rect 47852 5794 47908 5796
rect 47852 5742 47854 5794
rect 47854 5742 47906 5794
rect 47906 5742 47908 5794
rect 47852 5740 47908 5742
rect 47964 5404 48020 5460
rect 48188 5682 48244 5684
rect 48188 5630 48190 5682
rect 48190 5630 48242 5682
rect 48242 5630 48244 5682
rect 48188 5628 48244 5630
rect 47180 5068 47236 5124
rect 48076 5068 48132 5124
rect 47516 4396 47572 4452
rect 46956 3724 47012 3780
rect 45724 2716 45780 2772
rect 38444 2156 38500 2212
rect 47404 3724 47460 3780
rect 47852 4226 47908 4228
rect 47852 4174 47854 4226
rect 47854 4174 47906 4226
rect 47906 4174 47908 4226
rect 47852 4172 47908 4174
rect 48972 9660 49028 9716
rect 48748 8146 48804 8148
rect 48748 8094 48750 8146
rect 48750 8094 48802 8146
rect 48802 8094 48804 8146
rect 48748 8092 48804 8094
rect 48748 7868 48804 7924
rect 49532 18956 49588 19012
rect 49532 18508 49588 18564
rect 51286 21194 51342 21196
rect 51286 21142 51288 21194
rect 51288 21142 51340 21194
rect 51340 21142 51342 21194
rect 51286 21140 51342 21142
rect 51390 21194 51446 21196
rect 51390 21142 51392 21194
rect 51392 21142 51444 21194
rect 51444 21142 51446 21194
rect 51390 21140 51446 21142
rect 51494 21194 51550 21196
rect 51494 21142 51496 21194
rect 51496 21142 51548 21194
rect 51548 21142 51550 21194
rect 51494 21140 51550 21142
rect 51548 20972 51604 21028
rect 51212 20860 51268 20916
rect 51996 20412 52052 20468
rect 51212 20076 51268 20132
rect 51996 20076 52052 20132
rect 49980 19516 50036 19572
rect 49756 19122 49812 19124
rect 49756 19070 49758 19122
rect 49758 19070 49810 19122
rect 49810 19070 49812 19122
rect 49756 19068 49812 19070
rect 50204 19404 50260 19460
rect 50316 19068 50372 19124
rect 50428 19628 50484 19684
rect 50540 19292 50596 19348
rect 49532 17388 49588 17444
rect 49868 17052 49924 17108
rect 50204 18450 50260 18452
rect 50204 18398 50206 18450
rect 50206 18398 50258 18450
rect 50258 18398 50260 18450
rect 50204 18396 50260 18398
rect 50092 18172 50148 18228
rect 49980 16940 50036 16996
rect 50092 17388 50148 17444
rect 49532 16098 49588 16100
rect 49532 16046 49534 16098
rect 49534 16046 49586 16098
rect 49586 16046 49588 16098
rect 49532 16044 49588 16046
rect 49980 15932 50036 15988
rect 50428 18562 50484 18564
rect 50428 18510 50430 18562
rect 50430 18510 50482 18562
rect 50482 18510 50484 18562
rect 50428 18508 50484 18510
rect 51286 19626 51342 19628
rect 51286 19574 51288 19626
rect 51288 19574 51340 19626
rect 51340 19574 51342 19626
rect 51286 19572 51342 19574
rect 51390 19626 51446 19628
rect 51390 19574 51392 19626
rect 51392 19574 51444 19626
rect 51444 19574 51446 19626
rect 51390 19572 51446 19574
rect 51494 19626 51550 19628
rect 51494 19574 51496 19626
rect 51496 19574 51548 19626
rect 51548 19574 51550 19626
rect 51494 19572 51550 19574
rect 51548 19346 51604 19348
rect 51548 19294 51550 19346
rect 51550 19294 51602 19346
rect 51602 19294 51604 19346
rect 51548 19292 51604 19294
rect 50764 18450 50820 18452
rect 50764 18398 50766 18450
rect 50766 18398 50818 18450
rect 50818 18398 50820 18450
rect 50764 18396 50820 18398
rect 50428 17164 50484 17220
rect 50316 16380 50372 16436
rect 50652 16716 50708 16772
rect 51772 19234 51828 19236
rect 51772 19182 51774 19234
rect 51774 19182 51826 19234
rect 51826 19182 51828 19234
rect 51772 19180 51828 19182
rect 51286 18058 51342 18060
rect 51286 18006 51288 18058
rect 51288 18006 51340 18058
rect 51340 18006 51342 18058
rect 51286 18004 51342 18006
rect 51390 18058 51446 18060
rect 51390 18006 51392 18058
rect 51392 18006 51444 18058
rect 51444 18006 51446 18058
rect 51390 18004 51446 18006
rect 51494 18058 51550 18060
rect 51494 18006 51496 18058
rect 51496 18006 51548 18058
rect 51548 18006 51550 18058
rect 51494 18004 51550 18006
rect 52220 24780 52276 24836
rect 52556 24668 52612 24724
rect 53340 25282 53396 25284
rect 53340 25230 53342 25282
rect 53342 25230 53394 25282
rect 53394 25230 53396 25282
rect 53340 25228 53396 25230
rect 53116 24668 53172 24724
rect 53116 24108 53172 24164
rect 53340 24050 53396 24052
rect 53340 23998 53342 24050
rect 53342 23998 53394 24050
rect 53394 23998 53396 24050
rect 53340 23996 53396 23998
rect 52892 23826 52948 23828
rect 52892 23774 52894 23826
rect 52894 23774 52946 23826
rect 52946 23774 52948 23826
rect 52892 23772 52948 23774
rect 52780 23714 52836 23716
rect 52780 23662 52782 23714
rect 52782 23662 52834 23714
rect 52834 23662 52836 23714
rect 52780 23660 52836 23662
rect 52892 22370 52948 22372
rect 52892 22318 52894 22370
rect 52894 22318 52946 22370
rect 52946 22318 52948 22370
rect 52892 22316 52948 22318
rect 52444 22204 52500 22260
rect 52220 21868 52276 21924
rect 53116 22092 53172 22148
rect 52892 20690 52948 20692
rect 52892 20638 52894 20690
rect 52894 20638 52946 20690
rect 52946 20638 52948 20690
rect 52892 20636 52948 20638
rect 52108 19740 52164 19796
rect 53116 20188 53172 20244
rect 52780 20076 52836 20132
rect 52556 19964 52612 20020
rect 53004 20130 53060 20132
rect 53004 20078 53006 20130
rect 53006 20078 53058 20130
rect 53058 20078 53060 20130
rect 53004 20076 53060 20078
rect 52668 19346 52724 19348
rect 52668 19294 52670 19346
rect 52670 19294 52722 19346
rect 52722 19294 52724 19346
rect 52668 19292 52724 19294
rect 52892 19234 52948 19236
rect 52892 19182 52894 19234
rect 52894 19182 52946 19234
rect 52946 19182 52948 19234
rect 52892 19180 52948 19182
rect 53676 21644 53732 21700
rect 54012 26572 54068 26628
rect 54124 26962 54180 26964
rect 54124 26910 54126 26962
rect 54126 26910 54178 26962
rect 54178 26910 54180 26962
rect 54124 26908 54180 26910
rect 54012 26348 54068 26404
rect 54124 26124 54180 26180
rect 54236 25394 54292 25396
rect 54236 25342 54238 25394
rect 54238 25342 54290 25394
rect 54290 25342 54292 25394
rect 54236 25340 54292 25342
rect 54124 25282 54180 25284
rect 54124 25230 54126 25282
rect 54126 25230 54178 25282
rect 54178 25230 54180 25282
rect 54124 25228 54180 25230
rect 55132 27858 55188 27860
rect 55132 27806 55134 27858
rect 55134 27806 55186 27858
rect 55186 27806 55188 27858
rect 55132 27804 55188 27806
rect 54796 27580 54852 27636
rect 54796 27132 54852 27188
rect 55132 26572 55188 26628
rect 56364 28642 56420 28644
rect 56364 28590 56366 28642
rect 56366 28590 56418 28642
rect 56418 28590 56420 28642
rect 56364 28588 56420 28590
rect 56924 28476 56980 28532
rect 57372 30156 57428 30212
rect 58439 34522 58495 34524
rect 58439 34470 58441 34522
rect 58441 34470 58493 34522
rect 58493 34470 58495 34522
rect 58439 34468 58495 34470
rect 58543 34522 58599 34524
rect 58543 34470 58545 34522
rect 58545 34470 58597 34522
rect 58597 34470 58599 34522
rect 58543 34468 58599 34470
rect 58647 34522 58703 34524
rect 58647 34470 58649 34522
rect 58649 34470 58701 34522
rect 58701 34470 58703 34522
rect 58647 34468 58703 34470
rect 58439 32954 58495 32956
rect 58439 32902 58441 32954
rect 58441 32902 58493 32954
rect 58493 32902 58495 32954
rect 58439 32900 58495 32902
rect 58543 32954 58599 32956
rect 58543 32902 58545 32954
rect 58545 32902 58597 32954
rect 58597 32902 58599 32954
rect 58543 32900 58599 32902
rect 58647 32954 58703 32956
rect 58647 32902 58649 32954
rect 58649 32902 58701 32954
rect 58701 32902 58703 32954
rect 58647 32900 58703 32902
rect 58268 32620 58324 32676
rect 58044 31106 58100 31108
rect 58044 31054 58046 31106
rect 58046 31054 58098 31106
rect 58098 31054 58100 31106
rect 58044 31052 58100 31054
rect 58156 31836 58212 31892
rect 57596 30098 57652 30100
rect 57596 30046 57598 30098
rect 57598 30046 57650 30098
rect 57650 30046 57652 30098
rect 57596 30044 57652 30046
rect 57372 28530 57428 28532
rect 57372 28478 57374 28530
rect 57374 28478 57426 28530
rect 57426 28478 57428 28530
rect 57372 28476 57428 28478
rect 56028 27074 56084 27076
rect 56028 27022 56030 27074
rect 56030 27022 56082 27074
rect 56082 27022 56084 27074
rect 56028 27020 56084 27022
rect 55132 25506 55188 25508
rect 55132 25454 55134 25506
rect 55134 25454 55186 25506
rect 55186 25454 55188 25506
rect 55132 25452 55188 25454
rect 54684 24722 54740 24724
rect 54684 24670 54686 24722
rect 54686 24670 54738 24722
rect 54738 24670 54740 24722
rect 54684 24668 54740 24670
rect 54684 24444 54740 24500
rect 54348 23154 54404 23156
rect 54348 23102 54350 23154
rect 54350 23102 54402 23154
rect 54402 23102 54404 23154
rect 54348 23100 54404 23102
rect 54460 22988 54516 23044
rect 54236 22876 54292 22932
rect 54348 21810 54404 21812
rect 54348 21758 54350 21810
rect 54350 21758 54402 21810
rect 54402 21758 54404 21810
rect 54348 21756 54404 21758
rect 53564 20524 53620 20580
rect 53788 19852 53844 19908
rect 53900 19458 53956 19460
rect 53900 19406 53902 19458
rect 53902 19406 53954 19458
rect 53954 19406 53956 19458
rect 53900 19404 53956 19406
rect 50988 17388 51044 17444
rect 50764 17276 50820 17332
rect 50876 17164 50932 17220
rect 51212 17052 51268 17108
rect 50428 15372 50484 15428
rect 50652 16044 50708 16100
rect 49868 14924 49924 14980
rect 49644 14252 49700 14308
rect 49420 13356 49476 13412
rect 49532 12962 49588 12964
rect 49532 12910 49534 12962
rect 49534 12910 49586 12962
rect 49586 12910 49588 12962
rect 49532 12908 49588 12910
rect 49420 11676 49476 11732
rect 49756 11394 49812 11396
rect 49756 11342 49758 11394
rect 49758 11342 49810 11394
rect 49810 11342 49812 11394
rect 49756 11340 49812 11342
rect 50204 14588 50260 14644
rect 50428 13804 50484 13860
rect 50316 13634 50372 13636
rect 50316 13582 50318 13634
rect 50318 13582 50370 13634
rect 50370 13582 50372 13634
rect 50316 13580 50372 13582
rect 50540 12908 50596 12964
rect 50652 14924 50708 14980
rect 51286 16490 51342 16492
rect 51286 16438 51288 16490
rect 51288 16438 51340 16490
rect 51340 16438 51342 16490
rect 51286 16436 51342 16438
rect 51390 16490 51446 16492
rect 51390 16438 51392 16490
rect 51392 16438 51444 16490
rect 51444 16438 51446 16490
rect 51390 16436 51446 16438
rect 51494 16490 51550 16492
rect 51494 16438 51496 16490
rect 51496 16438 51548 16490
rect 51548 16438 51550 16490
rect 51494 16436 51550 16438
rect 51548 16268 51604 16324
rect 51548 15314 51604 15316
rect 51548 15262 51550 15314
rect 51550 15262 51602 15314
rect 51602 15262 51604 15314
rect 51548 15260 51604 15262
rect 53116 17666 53172 17668
rect 53116 17614 53118 17666
rect 53118 17614 53170 17666
rect 53170 17614 53172 17666
rect 53116 17612 53172 17614
rect 51884 16770 51940 16772
rect 51884 16718 51886 16770
rect 51886 16718 51938 16770
rect 51938 16718 51940 16770
rect 51884 16716 51940 16718
rect 52780 16604 52836 16660
rect 52892 16716 52948 16772
rect 53564 16828 53620 16884
rect 53340 16604 53396 16660
rect 52444 15426 52500 15428
rect 52444 15374 52446 15426
rect 52446 15374 52498 15426
rect 52498 15374 52500 15426
rect 52444 15372 52500 15374
rect 52892 15260 52948 15316
rect 51660 15202 51716 15204
rect 51660 15150 51662 15202
rect 51662 15150 51714 15202
rect 51714 15150 51716 15202
rect 51660 15148 51716 15150
rect 52556 15148 52612 15204
rect 51286 14922 51342 14924
rect 51286 14870 51288 14922
rect 51288 14870 51340 14922
rect 51340 14870 51342 14922
rect 51286 14868 51342 14870
rect 51390 14922 51446 14924
rect 51390 14870 51392 14922
rect 51392 14870 51444 14922
rect 51444 14870 51446 14922
rect 51390 14868 51446 14870
rect 51494 14922 51550 14924
rect 51494 14870 51496 14922
rect 51496 14870 51548 14922
rect 51548 14870 51550 14922
rect 51494 14868 51550 14870
rect 51100 14700 51156 14756
rect 50764 12908 50820 12964
rect 51286 13354 51342 13356
rect 51286 13302 51288 13354
rect 51288 13302 51340 13354
rect 51340 13302 51342 13354
rect 51286 13300 51342 13302
rect 51390 13354 51446 13356
rect 51390 13302 51392 13354
rect 51392 13302 51444 13354
rect 51444 13302 51446 13354
rect 51390 13300 51446 13302
rect 51494 13354 51550 13356
rect 51494 13302 51496 13354
rect 51496 13302 51548 13354
rect 51548 13302 51550 13354
rect 51494 13300 51550 13302
rect 51100 12796 51156 12852
rect 51212 12236 51268 12292
rect 51996 14530 52052 14532
rect 51996 14478 51998 14530
rect 51998 14478 52050 14530
rect 52050 14478 52052 14530
rect 51996 14476 52052 14478
rect 52780 15148 52836 15204
rect 53228 15372 53284 15428
rect 52444 14140 52500 14196
rect 51772 13580 51828 13636
rect 51100 12012 51156 12068
rect 50764 11900 50820 11956
rect 50092 11676 50148 11732
rect 50652 11676 50708 11732
rect 50540 11394 50596 11396
rect 50540 11342 50542 11394
rect 50542 11342 50594 11394
rect 50594 11342 50596 11394
rect 50540 11340 50596 11342
rect 50652 10050 50708 10052
rect 50652 9998 50654 10050
rect 50654 9998 50706 10050
rect 50706 9998 50708 10050
rect 50652 9996 50708 9998
rect 49756 9772 49812 9828
rect 52108 12236 52164 12292
rect 51436 11900 51492 11956
rect 51286 11786 51342 11788
rect 51286 11734 51288 11786
rect 51288 11734 51340 11786
rect 51340 11734 51342 11786
rect 51286 11732 51342 11734
rect 51390 11786 51446 11788
rect 51390 11734 51392 11786
rect 51392 11734 51444 11786
rect 51444 11734 51446 11786
rect 51390 11732 51446 11734
rect 51494 11786 51550 11788
rect 51494 11734 51496 11786
rect 51496 11734 51548 11786
rect 51548 11734 51550 11786
rect 51494 11732 51550 11734
rect 51772 12012 51828 12068
rect 52332 11900 52388 11956
rect 51286 10218 51342 10220
rect 51286 10166 51288 10218
rect 51288 10166 51340 10218
rect 51340 10166 51342 10218
rect 51286 10164 51342 10166
rect 51390 10218 51446 10220
rect 51390 10166 51392 10218
rect 51392 10166 51444 10218
rect 51444 10166 51446 10218
rect 51390 10164 51446 10166
rect 51494 10218 51550 10220
rect 51494 10166 51496 10218
rect 51496 10166 51548 10218
rect 51548 10166 51550 10218
rect 51494 10164 51550 10166
rect 49756 9100 49812 9156
rect 50204 9324 50260 9380
rect 49980 8818 50036 8820
rect 49980 8766 49982 8818
rect 49982 8766 50034 8818
rect 50034 8766 50036 8818
rect 49980 8764 50036 8766
rect 50316 8764 50372 8820
rect 49196 7420 49252 7476
rect 49532 7532 49588 7588
rect 50316 7586 50372 7588
rect 50316 7534 50318 7586
rect 50318 7534 50370 7586
rect 50370 7534 50372 7586
rect 50316 7532 50372 7534
rect 50540 7474 50596 7476
rect 50540 7422 50542 7474
rect 50542 7422 50594 7474
rect 50594 7422 50596 7474
rect 50540 7420 50596 7422
rect 48860 6524 48916 6580
rect 50428 6636 50484 6692
rect 50316 6578 50372 6580
rect 50316 6526 50318 6578
rect 50318 6526 50370 6578
rect 50370 6526 50372 6578
rect 50316 6524 50372 6526
rect 48972 5628 49028 5684
rect 48972 5346 49028 5348
rect 48972 5294 48974 5346
rect 48974 5294 49026 5346
rect 49026 5294 49028 5346
rect 48972 5292 49028 5294
rect 48748 5122 48804 5124
rect 48748 5070 48750 5122
rect 48750 5070 48802 5122
rect 48802 5070 48804 5122
rect 48748 5068 48804 5070
rect 50428 5906 50484 5908
rect 50428 5854 50430 5906
rect 50430 5854 50482 5906
rect 50482 5854 50484 5906
rect 50428 5852 50484 5854
rect 49756 5794 49812 5796
rect 49756 5742 49758 5794
rect 49758 5742 49810 5794
rect 49810 5742 49812 5794
rect 49756 5740 49812 5742
rect 49756 5404 49812 5460
rect 50204 5068 50260 5124
rect 49308 4956 49364 5012
rect 50988 9324 51044 9380
rect 50988 9154 51044 9156
rect 50988 9102 50990 9154
rect 50990 9102 51042 9154
rect 51042 9102 51044 9154
rect 50988 9100 51044 9102
rect 51660 9772 51716 9828
rect 51884 9660 51940 9716
rect 51286 8650 51342 8652
rect 51286 8598 51288 8650
rect 51288 8598 51340 8650
rect 51340 8598 51342 8650
rect 51286 8596 51342 8598
rect 51390 8650 51446 8652
rect 51390 8598 51392 8650
rect 51392 8598 51444 8650
rect 51444 8598 51446 8650
rect 51390 8596 51446 8598
rect 51494 8650 51550 8652
rect 51494 8598 51496 8650
rect 51496 8598 51548 8650
rect 51548 8598 51550 8650
rect 51494 8596 51550 8598
rect 52332 9324 52388 9380
rect 52108 8540 52164 8596
rect 51436 8204 51492 8260
rect 51772 7532 51828 7588
rect 51548 7308 51604 7364
rect 51286 7082 51342 7084
rect 51286 7030 51288 7082
rect 51288 7030 51340 7082
rect 51340 7030 51342 7082
rect 51286 7028 51342 7030
rect 51390 7082 51446 7084
rect 51390 7030 51392 7082
rect 51392 7030 51444 7082
rect 51444 7030 51446 7082
rect 51390 7028 51446 7030
rect 51494 7082 51550 7084
rect 51494 7030 51496 7082
rect 51496 7030 51548 7082
rect 51548 7030 51550 7082
rect 51494 7028 51550 7030
rect 51772 7084 51828 7140
rect 50876 6578 50932 6580
rect 50876 6526 50878 6578
rect 50878 6526 50930 6578
rect 50930 6526 50932 6578
rect 50876 6524 50932 6526
rect 51324 6578 51380 6580
rect 51324 6526 51326 6578
rect 51326 6526 51378 6578
rect 51378 6526 51380 6578
rect 51324 6524 51380 6526
rect 50764 5180 50820 5236
rect 51884 6972 51940 7028
rect 50988 5404 51044 5460
rect 51286 5514 51342 5516
rect 51286 5462 51288 5514
rect 51288 5462 51340 5514
rect 51340 5462 51342 5514
rect 51286 5460 51342 5462
rect 51390 5514 51446 5516
rect 51390 5462 51392 5514
rect 51392 5462 51444 5514
rect 51444 5462 51446 5514
rect 51390 5460 51446 5462
rect 51494 5514 51550 5516
rect 51494 5462 51496 5514
rect 51496 5462 51548 5514
rect 51548 5462 51550 5514
rect 51494 5460 51550 5462
rect 53004 13858 53060 13860
rect 53004 13806 53006 13858
rect 53006 13806 53058 13858
rect 53058 13806 53060 13858
rect 53004 13804 53060 13806
rect 53340 13634 53396 13636
rect 53340 13582 53342 13634
rect 53342 13582 53394 13634
rect 53394 13582 53396 13634
rect 53340 13580 53396 13582
rect 53116 9826 53172 9828
rect 53116 9774 53118 9826
rect 53118 9774 53170 9826
rect 53170 9774 53172 9826
rect 53116 9772 53172 9774
rect 52556 9660 52612 9716
rect 52892 9100 52948 9156
rect 52892 8540 52948 8596
rect 53116 9042 53172 9044
rect 53116 8990 53118 9042
rect 53118 8990 53170 9042
rect 53170 8990 53172 9042
rect 53116 8988 53172 8990
rect 52444 7644 52500 7700
rect 53004 8316 53060 8372
rect 54124 20802 54180 20804
rect 54124 20750 54126 20802
rect 54126 20750 54178 20802
rect 54178 20750 54180 20802
rect 54124 20748 54180 20750
rect 54460 20636 54516 20692
rect 55916 26236 55972 26292
rect 55692 26178 55748 26180
rect 55692 26126 55694 26178
rect 55694 26126 55746 26178
rect 55746 26126 55748 26178
rect 55692 26124 55748 26126
rect 55804 25452 55860 25508
rect 55916 25564 55972 25620
rect 56476 26460 56532 26516
rect 56700 26178 56756 26180
rect 56700 26126 56702 26178
rect 56702 26126 56754 26178
rect 56754 26126 56756 26178
rect 56700 26124 56756 26126
rect 54908 22988 54964 23044
rect 55020 22876 55076 22932
rect 55020 22594 55076 22596
rect 55020 22542 55022 22594
rect 55022 22542 55074 22594
rect 55074 22542 55076 22594
rect 55020 22540 55076 22542
rect 55468 22652 55524 22708
rect 57260 27074 57316 27076
rect 57260 27022 57262 27074
rect 57262 27022 57314 27074
rect 57314 27022 57316 27074
rect 57260 27020 57316 27022
rect 57932 29484 57988 29540
rect 57820 28812 57876 28868
rect 57484 27244 57540 27300
rect 57372 26796 57428 26852
rect 56028 23100 56084 23156
rect 56252 23826 56308 23828
rect 56252 23774 56254 23826
rect 56254 23774 56306 23826
rect 56306 23774 56308 23826
rect 56252 23772 56308 23774
rect 55244 21532 55300 21588
rect 54796 20412 54852 20468
rect 55692 21810 55748 21812
rect 55692 21758 55694 21810
rect 55694 21758 55746 21810
rect 55746 21758 55748 21810
rect 55692 21756 55748 21758
rect 55916 21698 55972 21700
rect 55916 21646 55918 21698
rect 55918 21646 55970 21698
rect 55970 21646 55972 21698
rect 55916 21644 55972 21646
rect 55692 20578 55748 20580
rect 55692 20526 55694 20578
rect 55694 20526 55746 20578
rect 55746 20526 55748 20578
rect 55692 20524 55748 20526
rect 56140 20412 56196 20468
rect 55804 20076 55860 20132
rect 55020 19180 55076 19236
rect 55132 18450 55188 18452
rect 55132 18398 55134 18450
rect 55134 18398 55186 18450
rect 55186 18398 55188 18450
rect 55132 18396 55188 18398
rect 54796 18284 54852 18340
rect 54460 17724 54516 17780
rect 54684 17554 54740 17556
rect 54684 17502 54686 17554
rect 54686 17502 54738 17554
rect 54738 17502 54740 17554
rect 54684 17500 54740 17502
rect 54348 16828 54404 16884
rect 55244 17778 55300 17780
rect 55244 17726 55246 17778
rect 55246 17726 55298 17778
rect 55298 17726 55300 17778
rect 55244 17724 55300 17726
rect 54908 16828 54964 16884
rect 55132 16882 55188 16884
rect 55132 16830 55134 16882
rect 55134 16830 55186 16882
rect 55186 16830 55188 16882
rect 55132 16828 55188 16830
rect 54796 15148 54852 15204
rect 55132 15372 55188 15428
rect 54908 14588 54964 14644
rect 56028 19852 56084 19908
rect 55916 19404 55972 19460
rect 57036 23772 57092 23828
rect 57148 26290 57204 26292
rect 57148 26238 57150 26290
rect 57150 26238 57202 26290
rect 57202 26238 57204 26290
rect 57148 26236 57204 26238
rect 56476 23660 56532 23716
rect 55692 19234 55748 19236
rect 55692 19182 55694 19234
rect 55694 19182 55746 19234
rect 55746 19182 55748 19234
rect 55692 19180 55748 19182
rect 55580 18338 55636 18340
rect 55580 18286 55582 18338
rect 55582 18286 55634 18338
rect 55634 18286 55636 18338
rect 55580 18284 55636 18286
rect 56028 18284 56084 18340
rect 55692 17836 55748 17892
rect 55580 17666 55636 17668
rect 55580 17614 55582 17666
rect 55582 17614 55634 17666
rect 55634 17614 55636 17666
rect 55580 17612 55636 17614
rect 55580 17388 55636 17444
rect 56028 17388 56084 17444
rect 55916 17106 55972 17108
rect 55916 17054 55918 17106
rect 55918 17054 55970 17106
rect 55970 17054 55972 17106
rect 55916 17052 55972 17054
rect 55692 16828 55748 16884
rect 55916 15484 55972 15540
rect 55804 15148 55860 15204
rect 56028 15426 56084 15428
rect 56028 15374 56030 15426
rect 56030 15374 56082 15426
rect 56082 15374 56084 15426
rect 56028 15372 56084 15374
rect 56140 15148 56196 15204
rect 55804 14530 55860 14532
rect 55804 14478 55806 14530
rect 55806 14478 55858 14530
rect 55858 14478 55860 14530
rect 55804 14476 55860 14478
rect 54908 13804 54964 13860
rect 56140 14642 56196 14644
rect 56140 14590 56142 14642
rect 56142 14590 56194 14642
rect 56194 14590 56196 14642
rect 56140 14588 56196 14590
rect 56252 14476 56308 14532
rect 55244 12236 55300 12292
rect 55468 13074 55524 13076
rect 55468 13022 55470 13074
rect 55470 13022 55522 13074
rect 55522 13022 55524 13074
rect 55468 13020 55524 13022
rect 54908 11954 54964 11956
rect 54908 11902 54910 11954
rect 54910 11902 54962 11954
rect 54962 11902 54964 11954
rect 54908 11900 54964 11902
rect 56140 12236 56196 12292
rect 55580 12066 55636 12068
rect 55580 12014 55582 12066
rect 55582 12014 55634 12066
rect 55634 12014 55636 12066
rect 55580 12012 55636 12014
rect 56140 11788 56196 11844
rect 53900 10834 53956 10836
rect 53900 10782 53902 10834
rect 53902 10782 53954 10834
rect 53954 10782 53956 10834
rect 53900 10780 53956 10782
rect 53900 10108 53956 10164
rect 53788 9154 53844 9156
rect 53788 9102 53790 9154
rect 53790 9102 53842 9154
rect 53842 9102 53844 9154
rect 53788 9100 53844 9102
rect 54012 8988 54068 9044
rect 54460 9772 54516 9828
rect 54908 10108 54964 10164
rect 55132 9826 55188 9828
rect 55132 9774 55134 9826
rect 55134 9774 55186 9826
rect 55186 9774 55188 9826
rect 55132 9772 55188 9774
rect 54908 8988 54964 9044
rect 54348 8316 54404 8372
rect 54572 8876 54628 8932
rect 54684 8370 54740 8372
rect 54684 8318 54686 8370
rect 54686 8318 54738 8370
rect 54738 8318 54740 8370
rect 54684 8316 54740 8318
rect 54572 8204 54628 8260
rect 55916 9996 55972 10052
rect 55692 8988 55748 9044
rect 55356 8428 55412 8484
rect 55916 8818 55972 8820
rect 55916 8766 55918 8818
rect 55918 8766 55970 8818
rect 55970 8766 55972 8818
rect 55916 8764 55972 8766
rect 53340 8034 53396 8036
rect 53340 7982 53342 8034
rect 53342 7982 53394 8034
rect 53394 7982 53396 8034
rect 53340 7980 53396 7982
rect 54124 7586 54180 7588
rect 54124 7534 54126 7586
rect 54126 7534 54178 7586
rect 54178 7534 54180 7586
rect 54124 7532 54180 7534
rect 54908 7980 54964 8036
rect 53452 6972 53508 7028
rect 53228 6748 53284 6804
rect 53004 6690 53060 6692
rect 53004 6638 53006 6690
rect 53006 6638 53058 6690
rect 53058 6638 53060 6690
rect 53004 6636 53060 6638
rect 53452 6524 53508 6580
rect 51436 5122 51492 5124
rect 51436 5070 51438 5122
rect 51438 5070 51490 5122
rect 51490 5070 51492 5122
rect 51436 5068 51492 5070
rect 51660 5122 51716 5124
rect 51660 5070 51662 5122
rect 51662 5070 51714 5122
rect 51714 5070 51716 5122
rect 51660 5068 51716 5070
rect 52108 5292 52164 5348
rect 53116 5292 53172 5348
rect 51212 5010 51268 5012
rect 51212 4958 51214 5010
rect 51214 4958 51266 5010
rect 51266 4958 51268 5010
rect 51212 4956 51268 4958
rect 53676 6578 53732 6580
rect 53676 6526 53678 6578
rect 53678 6526 53730 6578
rect 53730 6526 53732 6578
rect 53676 6524 53732 6526
rect 54012 6748 54068 6804
rect 54124 6636 54180 6692
rect 55020 7698 55076 7700
rect 55020 7646 55022 7698
rect 55022 7646 55074 7698
rect 55074 7646 55076 7698
rect 55020 7644 55076 7646
rect 55244 7308 55300 7364
rect 54796 6524 54852 6580
rect 54012 5122 54068 5124
rect 54012 5070 54014 5122
rect 54014 5070 54066 5122
rect 54066 5070 54068 5122
rect 54012 5068 54068 5070
rect 51100 4396 51156 4452
rect 52220 4956 52276 5012
rect 51996 4450 52052 4452
rect 51996 4398 51998 4450
rect 51998 4398 52050 4450
rect 52050 4398 52052 4450
rect 51996 4396 52052 4398
rect 54684 5292 54740 5348
rect 55468 8316 55524 8372
rect 57596 25564 57652 25620
rect 57260 24556 57316 24612
rect 58156 28476 58212 28532
rect 58156 24610 58212 24612
rect 58156 24558 58158 24610
rect 58158 24558 58210 24610
rect 58210 24558 58212 24610
rect 58156 24556 58212 24558
rect 57260 23660 57316 23716
rect 56924 23154 56980 23156
rect 56924 23102 56926 23154
rect 56926 23102 56978 23154
rect 56978 23102 56980 23154
rect 56924 23100 56980 23102
rect 56700 22540 56756 22596
rect 57260 22370 57316 22372
rect 57260 22318 57262 22370
rect 57262 22318 57314 22370
rect 57314 22318 57316 22370
rect 57260 22316 57316 22318
rect 57596 22316 57652 22372
rect 56812 20524 56868 20580
rect 56700 20412 56756 20468
rect 57036 20076 57092 20132
rect 56588 19906 56644 19908
rect 56588 19854 56590 19906
rect 56590 19854 56642 19906
rect 56642 19854 56644 19906
rect 56588 19852 56644 19854
rect 56812 19404 56868 19460
rect 56812 18338 56868 18340
rect 56812 18286 56814 18338
rect 56814 18286 56866 18338
rect 56866 18286 56868 18338
rect 56812 18284 56868 18286
rect 56812 16882 56868 16884
rect 56812 16830 56814 16882
rect 56814 16830 56866 16882
rect 56866 16830 56868 16882
rect 56812 16828 56868 16830
rect 57148 17612 57204 17668
rect 57036 17500 57092 17556
rect 57148 17052 57204 17108
rect 57372 21586 57428 21588
rect 57372 21534 57374 21586
rect 57374 21534 57426 21586
rect 57426 21534 57428 21586
rect 57372 21532 57428 21534
rect 58044 21532 58100 21588
rect 57708 17554 57764 17556
rect 57708 17502 57710 17554
rect 57710 17502 57762 17554
rect 57762 17502 57764 17554
rect 57708 17500 57764 17502
rect 57932 17442 57988 17444
rect 57932 17390 57934 17442
rect 57934 17390 57986 17442
rect 57986 17390 57988 17442
rect 57932 17388 57988 17390
rect 57484 15538 57540 15540
rect 57484 15486 57486 15538
rect 57486 15486 57538 15538
rect 57538 15486 57540 15538
rect 57484 15484 57540 15486
rect 57260 14140 57316 14196
rect 56588 12290 56644 12292
rect 56588 12238 56590 12290
rect 56590 12238 56642 12290
rect 56642 12238 56644 12290
rect 56588 12236 56644 12238
rect 57708 15148 57764 15204
rect 57820 14140 57876 14196
rect 57372 13244 57428 13300
rect 57484 13132 57540 13188
rect 57148 12236 57204 12292
rect 56812 12012 56868 12068
rect 57372 12012 57428 12068
rect 56812 11788 56868 11844
rect 57148 11788 57204 11844
rect 58439 31386 58495 31388
rect 58439 31334 58441 31386
rect 58441 31334 58493 31386
rect 58493 31334 58495 31386
rect 58439 31332 58495 31334
rect 58543 31386 58599 31388
rect 58543 31334 58545 31386
rect 58545 31334 58597 31386
rect 58597 31334 58599 31386
rect 58543 31332 58599 31334
rect 58647 31386 58703 31388
rect 58647 31334 58649 31386
rect 58649 31334 58701 31386
rect 58701 31334 58703 31386
rect 58647 31332 58703 31334
rect 58439 29818 58495 29820
rect 58439 29766 58441 29818
rect 58441 29766 58493 29818
rect 58493 29766 58495 29818
rect 58439 29764 58495 29766
rect 58543 29818 58599 29820
rect 58543 29766 58545 29818
rect 58545 29766 58597 29818
rect 58597 29766 58599 29818
rect 58543 29764 58599 29766
rect 58647 29818 58703 29820
rect 58647 29766 58649 29818
rect 58649 29766 58701 29818
rect 58701 29766 58703 29818
rect 58647 29764 58703 29766
rect 58439 28250 58495 28252
rect 58439 28198 58441 28250
rect 58441 28198 58493 28250
rect 58493 28198 58495 28250
rect 58439 28196 58495 28198
rect 58543 28250 58599 28252
rect 58543 28198 58545 28250
rect 58545 28198 58597 28250
rect 58597 28198 58599 28250
rect 58543 28196 58599 28198
rect 58647 28250 58703 28252
rect 58647 28198 58649 28250
rect 58649 28198 58701 28250
rect 58701 28198 58703 28250
rect 58647 28196 58703 28198
rect 58439 26682 58495 26684
rect 58439 26630 58441 26682
rect 58441 26630 58493 26682
rect 58493 26630 58495 26682
rect 58439 26628 58495 26630
rect 58543 26682 58599 26684
rect 58543 26630 58545 26682
rect 58545 26630 58597 26682
rect 58597 26630 58599 26682
rect 58543 26628 58599 26630
rect 58647 26682 58703 26684
rect 58647 26630 58649 26682
rect 58649 26630 58701 26682
rect 58701 26630 58703 26682
rect 58647 26628 58703 26630
rect 58439 25114 58495 25116
rect 58439 25062 58441 25114
rect 58441 25062 58493 25114
rect 58493 25062 58495 25114
rect 58439 25060 58495 25062
rect 58543 25114 58599 25116
rect 58543 25062 58545 25114
rect 58545 25062 58597 25114
rect 58597 25062 58599 25114
rect 58543 25060 58599 25062
rect 58647 25114 58703 25116
rect 58647 25062 58649 25114
rect 58649 25062 58701 25114
rect 58701 25062 58703 25114
rect 58647 25060 58703 25062
rect 58439 23546 58495 23548
rect 58439 23494 58441 23546
rect 58441 23494 58493 23546
rect 58493 23494 58495 23546
rect 58439 23492 58495 23494
rect 58543 23546 58599 23548
rect 58543 23494 58545 23546
rect 58545 23494 58597 23546
rect 58597 23494 58599 23546
rect 58543 23492 58599 23494
rect 58647 23546 58703 23548
rect 58647 23494 58649 23546
rect 58649 23494 58701 23546
rect 58701 23494 58703 23546
rect 58647 23492 58703 23494
rect 58439 21978 58495 21980
rect 58439 21926 58441 21978
rect 58441 21926 58493 21978
rect 58493 21926 58495 21978
rect 58439 21924 58495 21926
rect 58543 21978 58599 21980
rect 58543 21926 58545 21978
rect 58545 21926 58597 21978
rect 58597 21926 58599 21978
rect 58543 21924 58599 21926
rect 58647 21978 58703 21980
rect 58647 21926 58649 21978
rect 58649 21926 58701 21978
rect 58701 21926 58703 21978
rect 58647 21924 58703 21926
rect 58439 20410 58495 20412
rect 58439 20358 58441 20410
rect 58441 20358 58493 20410
rect 58493 20358 58495 20410
rect 58439 20356 58495 20358
rect 58543 20410 58599 20412
rect 58543 20358 58545 20410
rect 58545 20358 58597 20410
rect 58597 20358 58599 20410
rect 58543 20356 58599 20358
rect 58647 20410 58703 20412
rect 58647 20358 58649 20410
rect 58649 20358 58701 20410
rect 58701 20358 58703 20410
rect 58647 20356 58703 20358
rect 58439 18842 58495 18844
rect 58439 18790 58441 18842
rect 58441 18790 58493 18842
rect 58493 18790 58495 18842
rect 58439 18788 58495 18790
rect 58543 18842 58599 18844
rect 58543 18790 58545 18842
rect 58545 18790 58597 18842
rect 58597 18790 58599 18842
rect 58543 18788 58599 18790
rect 58647 18842 58703 18844
rect 58647 18790 58649 18842
rect 58649 18790 58701 18842
rect 58701 18790 58703 18842
rect 58647 18788 58703 18790
rect 58439 17274 58495 17276
rect 58439 17222 58441 17274
rect 58441 17222 58493 17274
rect 58493 17222 58495 17274
rect 58439 17220 58495 17222
rect 58543 17274 58599 17276
rect 58543 17222 58545 17274
rect 58545 17222 58597 17274
rect 58597 17222 58599 17274
rect 58543 17220 58599 17222
rect 58647 17274 58703 17276
rect 58647 17222 58649 17274
rect 58649 17222 58701 17274
rect 58701 17222 58703 17274
rect 58647 17220 58703 17222
rect 58439 15706 58495 15708
rect 58439 15654 58441 15706
rect 58441 15654 58493 15706
rect 58493 15654 58495 15706
rect 58439 15652 58495 15654
rect 58543 15706 58599 15708
rect 58543 15654 58545 15706
rect 58545 15654 58597 15706
rect 58597 15654 58599 15706
rect 58543 15652 58599 15654
rect 58647 15706 58703 15708
rect 58647 15654 58649 15706
rect 58649 15654 58701 15706
rect 58701 15654 58703 15706
rect 58647 15652 58703 15654
rect 58439 14138 58495 14140
rect 58439 14086 58441 14138
rect 58441 14086 58493 14138
rect 58493 14086 58495 14138
rect 58439 14084 58495 14086
rect 58543 14138 58599 14140
rect 58543 14086 58545 14138
rect 58545 14086 58597 14138
rect 58597 14086 58599 14138
rect 58543 14084 58599 14086
rect 58647 14138 58703 14140
rect 58647 14086 58649 14138
rect 58649 14086 58701 14138
rect 58701 14086 58703 14138
rect 58647 14084 58703 14086
rect 58044 13244 58100 13300
rect 57820 13132 57876 13188
rect 57820 11788 57876 11844
rect 56700 9996 56756 10052
rect 56588 9042 56644 9044
rect 56588 8990 56590 9042
rect 56590 8990 56642 9042
rect 56642 8990 56644 9042
rect 56588 8988 56644 8990
rect 56252 8370 56308 8372
rect 56252 8318 56254 8370
rect 56254 8318 56306 8370
rect 56306 8318 56308 8370
rect 56252 8316 56308 8318
rect 56924 8316 56980 8372
rect 55804 8204 55860 8260
rect 56476 8258 56532 8260
rect 56476 8206 56478 8258
rect 56478 8206 56530 8258
rect 56530 8206 56532 8258
rect 56476 8204 56532 8206
rect 58439 12570 58495 12572
rect 58439 12518 58441 12570
rect 58441 12518 58493 12570
rect 58493 12518 58495 12570
rect 58439 12516 58495 12518
rect 58543 12570 58599 12572
rect 58543 12518 58545 12570
rect 58545 12518 58597 12570
rect 58597 12518 58599 12570
rect 58543 12516 58599 12518
rect 58647 12570 58703 12572
rect 58647 12518 58649 12570
rect 58649 12518 58701 12570
rect 58701 12518 58703 12570
rect 58647 12516 58703 12518
rect 58439 11002 58495 11004
rect 58439 10950 58441 11002
rect 58441 10950 58493 11002
rect 58493 10950 58495 11002
rect 58439 10948 58495 10950
rect 58543 11002 58599 11004
rect 58543 10950 58545 11002
rect 58545 10950 58597 11002
rect 58597 10950 58599 11002
rect 58543 10948 58599 10950
rect 58647 11002 58703 11004
rect 58647 10950 58649 11002
rect 58649 10950 58701 11002
rect 58701 10950 58703 11002
rect 58647 10948 58703 10950
rect 58439 9434 58495 9436
rect 58439 9382 58441 9434
rect 58441 9382 58493 9434
rect 58493 9382 58495 9434
rect 58439 9380 58495 9382
rect 58543 9434 58599 9436
rect 58543 9382 58545 9434
rect 58545 9382 58597 9434
rect 58597 9382 58599 9434
rect 58543 9380 58599 9382
rect 58647 9434 58703 9436
rect 58647 9382 58649 9434
rect 58649 9382 58701 9434
rect 58701 9382 58703 9434
rect 58647 9380 58703 9382
rect 57484 8764 57540 8820
rect 57148 7644 57204 7700
rect 56812 6860 56868 6916
rect 57036 7308 57092 7364
rect 56140 6466 56196 6468
rect 56140 6414 56142 6466
rect 56142 6414 56194 6466
rect 56194 6414 56196 6466
rect 56140 6412 56196 6414
rect 57260 8204 57316 8260
rect 58439 7866 58495 7868
rect 58439 7814 58441 7866
rect 58441 7814 58493 7866
rect 58493 7814 58495 7866
rect 58439 7812 58495 7814
rect 58543 7866 58599 7868
rect 58543 7814 58545 7866
rect 58545 7814 58597 7866
rect 58597 7814 58599 7866
rect 58543 7812 58599 7814
rect 58647 7866 58703 7868
rect 58647 7814 58649 7866
rect 58649 7814 58701 7866
rect 58701 7814 58703 7866
rect 58647 7812 58703 7814
rect 57036 6300 57092 6356
rect 55692 5068 55748 5124
rect 56028 5906 56084 5908
rect 56028 5854 56030 5906
rect 56030 5854 56082 5906
rect 56082 5854 56084 5906
rect 56028 5852 56084 5854
rect 56588 5906 56644 5908
rect 56588 5854 56590 5906
rect 56590 5854 56642 5906
rect 56642 5854 56644 5906
rect 56588 5852 56644 5854
rect 57820 6412 57876 6468
rect 58044 6300 58100 6356
rect 58439 6298 58495 6300
rect 58439 6246 58441 6298
rect 58441 6246 58493 6298
rect 58493 6246 58495 6298
rect 58439 6244 58495 6246
rect 58543 6298 58599 6300
rect 58543 6246 58545 6298
rect 58545 6246 58597 6298
rect 58597 6246 58599 6298
rect 58543 6244 58599 6246
rect 58647 6298 58703 6300
rect 58647 6246 58649 6298
rect 58649 6246 58701 6298
rect 58701 6246 58703 6298
rect 58647 6244 58703 6246
rect 56252 5180 56308 5236
rect 56924 5180 56980 5236
rect 56588 5122 56644 5124
rect 56588 5070 56590 5122
rect 56590 5070 56642 5122
rect 56642 5070 56644 5122
rect 56588 5068 56644 5070
rect 58156 5906 58212 5908
rect 58156 5854 58158 5906
rect 58158 5854 58210 5906
rect 58210 5854 58212 5906
rect 58156 5852 58212 5854
rect 58044 5068 58100 5124
rect 58439 4730 58495 4732
rect 58439 4678 58441 4730
rect 58441 4678 58493 4730
rect 58493 4678 58495 4730
rect 58439 4676 58495 4678
rect 58543 4730 58599 4732
rect 58543 4678 58545 4730
rect 58545 4678 58597 4730
rect 58597 4678 58599 4730
rect 58543 4676 58599 4678
rect 58647 4730 58703 4732
rect 58647 4678 58649 4730
rect 58649 4678 58701 4730
rect 58701 4678 58703 4730
rect 58647 4676 58703 4678
rect 56588 4508 56644 4564
rect 51286 3946 51342 3948
rect 51286 3894 51288 3946
rect 51288 3894 51340 3946
rect 51340 3894 51342 3946
rect 51286 3892 51342 3894
rect 51390 3946 51446 3948
rect 51390 3894 51392 3946
rect 51392 3894 51444 3946
rect 51444 3894 51446 3946
rect 51390 3892 51446 3894
rect 51494 3946 51550 3948
rect 51494 3894 51496 3946
rect 51496 3894 51548 3946
rect 51548 3894 51550 3946
rect 51494 3892 51550 3894
rect 50652 3276 50708 3332
rect 52780 2604 52836 2660
rect 58439 3162 58495 3164
rect 58439 3110 58441 3162
rect 58441 3110 58493 3162
rect 58493 3110 58495 3162
rect 58439 3108 58495 3110
rect 58543 3162 58599 3164
rect 58543 3110 58545 3162
rect 58545 3110 58597 3162
rect 58597 3110 58599 3162
rect 58543 3108 58599 3110
rect 58647 3162 58703 3164
rect 58647 3110 58649 3162
rect 58649 3110 58701 3162
rect 58701 3110 58703 3162
rect 58647 3108 58703 3110
<< metal3 >>
rect 13794 37324 13804 37380
rect 13860 37324 45836 37380
rect 45892 37324 45902 37380
rect 0 37268 800 37296
rect 0 37212 3500 37268
rect 3556 37212 3566 37268
rect 27682 37212 27692 37268
rect 27748 37212 56252 37268
rect 56308 37212 56318 37268
rect 0 37184 800 37212
rect 28802 37100 28812 37156
rect 28868 37100 56364 37156
rect 56420 37100 56430 37156
rect 12226 36988 12236 37044
rect 12292 36988 33292 37044
rect 33348 36988 33358 37044
rect 34514 36988 34524 37044
rect 34580 36988 52108 37044
rect 52164 36988 52174 37044
rect 9650 36876 9660 36932
rect 9716 36876 10668 36932
rect 10724 36876 10734 36932
rect 16370 36876 16380 36932
rect 16436 36876 17388 36932
rect 17444 36876 17454 36932
rect 32050 36876 32060 36932
rect 32116 36876 33740 36932
rect 33796 36876 33806 36932
rect 41010 36876 41020 36932
rect 41076 36876 42252 36932
rect 42308 36876 43036 36932
rect 43092 36876 43102 36932
rect 8355 36820 8365 36876
rect 8421 36820 8469 36876
rect 8525 36820 8573 36876
rect 8629 36820 8639 36876
rect 22662 36820 22672 36876
rect 22728 36820 22776 36876
rect 22832 36820 22880 36876
rect 22936 36820 22946 36876
rect 36969 36820 36979 36876
rect 37035 36820 37083 36876
rect 37139 36820 37187 36876
rect 37243 36820 37253 36876
rect 51276 36820 51286 36876
rect 51342 36820 51390 36876
rect 51446 36820 51494 36876
rect 51550 36820 51560 36876
rect 11218 36764 11228 36820
rect 11284 36764 15148 36820
rect 15092 36708 15148 36764
rect 40796 36764 41916 36820
rect 41972 36764 41982 36820
rect 40796 36708 40852 36764
rect 15092 36652 40796 36708
rect 40852 36652 40862 36708
rect 41346 36652 41356 36708
rect 41412 36652 55020 36708
rect 55076 36652 55086 36708
rect 4610 36540 4620 36596
rect 4676 36540 5404 36596
rect 5460 36540 5470 36596
rect 12562 36540 12572 36596
rect 12628 36540 14364 36596
rect 14420 36540 14430 36596
rect 18050 36540 18060 36596
rect 18116 36540 35308 36596
rect 35364 36540 35374 36596
rect 37202 36540 37212 36596
rect 37268 36540 43932 36596
rect 43988 36540 43998 36596
rect 53788 36540 56924 36596
rect 56980 36540 56990 36596
rect 53788 36484 53844 36540
rect 1810 36428 1820 36484
rect 1876 36428 4172 36484
rect 4228 36428 4238 36484
rect 21186 36428 21196 36484
rect 21252 36428 25004 36484
rect 25060 36428 25070 36484
rect 32610 36428 32620 36484
rect 32676 36428 46732 36484
rect 46788 36428 46798 36484
rect 47730 36428 47740 36484
rect 47796 36428 48860 36484
rect 48916 36428 48926 36484
rect 52210 36428 52220 36484
rect 52276 36428 53788 36484
rect 53844 36428 53854 36484
rect 54450 36428 54460 36484
rect 54516 36428 55468 36484
rect 55524 36428 55534 36484
rect 6626 36316 6636 36372
rect 6692 36316 7868 36372
rect 7924 36316 7934 36372
rect 14018 36316 14028 36372
rect 14084 36316 15820 36372
rect 15876 36316 16492 36372
rect 16548 36316 16558 36372
rect 28354 36316 28364 36372
rect 28420 36316 29148 36372
rect 29204 36316 29214 36372
rect 38546 36316 38556 36372
rect 38612 36316 43540 36372
rect 46050 36316 46060 36372
rect 46116 36316 49196 36372
rect 49252 36316 49262 36372
rect 49970 36316 49980 36372
rect 50036 36316 50540 36372
rect 50596 36316 56476 36372
rect 56532 36316 56542 36372
rect 43484 36260 43540 36316
rect 13234 36204 13244 36260
rect 13300 36204 13692 36260
rect 13748 36204 15148 36260
rect 15204 36204 16156 36260
rect 16212 36204 18508 36260
rect 18564 36204 24668 36260
rect 24724 36204 24734 36260
rect 26674 36204 26684 36260
rect 26740 36204 28476 36260
rect 28532 36204 28542 36260
rect 43484 36204 48300 36260
rect 48356 36204 48366 36260
rect 55412 36204 56028 36260
rect 56084 36204 56094 36260
rect 0 36148 800 36176
rect 55412 36148 55468 36204
rect 0 36092 2604 36148
rect 2660 36092 2670 36148
rect 31826 36092 31836 36148
rect 31892 36092 43764 36148
rect 49298 36092 49308 36148
rect 49364 36092 55468 36148
rect 0 36064 800 36092
rect 15508 36036 15518 36092
rect 15574 36036 15622 36092
rect 15678 36036 15726 36092
rect 15782 36036 15792 36092
rect 29815 36036 29825 36092
rect 29881 36036 29929 36092
rect 29985 36036 30033 36092
rect 30089 36036 30099 36092
rect 20290 35980 20300 36036
rect 20356 35980 21308 36036
rect 21364 35980 22764 36036
rect 22820 35980 24332 36036
rect 24388 35980 24398 36036
rect 38612 35980 42756 36036
rect 38612 35924 38668 35980
rect 4946 35868 4956 35924
rect 5012 35868 21644 35924
rect 21700 35868 21710 35924
rect 22866 35868 22876 35924
rect 22932 35868 38668 35924
rect 42700 35812 42756 35980
rect 43708 35812 43764 36092
rect 44122 36036 44132 36092
rect 44188 36036 44236 36092
rect 44292 36036 44340 36092
rect 44396 36036 44406 36092
rect 58429 36036 58439 36092
rect 58495 36036 58543 36092
rect 58599 36036 58647 36092
rect 58703 36036 58713 36092
rect 46834 35980 46844 36036
rect 46900 35980 53564 36036
rect 53620 35980 53630 36036
rect 46722 35868 46732 35924
rect 46788 35868 51436 35924
rect 51492 35868 51502 35924
rect 52770 35868 52780 35924
rect 52836 35868 54684 35924
rect 54740 35868 54750 35924
rect 6962 35756 6972 35812
rect 7028 35756 26908 35812
rect 35522 35756 35532 35812
rect 35588 35756 35868 35812
rect 35924 35756 35934 35812
rect 36418 35756 36428 35812
rect 36484 35756 40908 35812
rect 40964 35756 40974 35812
rect 42690 35756 42700 35812
rect 42756 35756 42766 35812
rect 43708 35756 48748 35812
rect 48804 35756 48814 35812
rect 49074 35756 49084 35812
rect 49140 35756 51772 35812
rect 51828 35756 51838 35812
rect 51996 35756 55580 35812
rect 55636 35756 55646 35812
rect 26852 35700 26908 35756
rect 51996 35700 52052 35756
rect 4162 35644 4172 35700
rect 4228 35644 5068 35700
rect 5124 35644 5852 35700
rect 5908 35644 9044 35700
rect 21634 35644 21644 35700
rect 21700 35644 22652 35700
rect 22708 35644 22718 35700
rect 22866 35644 22876 35700
rect 22932 35644 22942 35700
rect 24658 35644 24668 35700
rect 24724 35644 26012 35700
rect 26068 35644 26684 35700
rect 26740 35644 26750 35700
rect 26852 35644 37772 35700
rect 37828 35644 37838 35700
rect 46050 35644 46060 35700
rect 46116 35644 50204 35700
rect 50260 35644 50270 35700
rect 50428 35644 52052 35700
rect 55234 35644 55244 35700
rect 55300 35644 56476 35700
rect 56532 35644 56542 35700
rect 8988 35588 9044 35644
rect 1698 35532 1708 35588
rect 1764 35532 8428 35588
rect 8978 35532 8988 35588
rect 9044 35532 9772 35588
rect 9828 35532 11116 35588
rect 11172 35532 12796 35588
rect 12852 35532 12862 35588
rect 15922 35532 15932 35588
rect 15988 35532 16940 35588
rect 16996 35532 17006 35588
rect 18162 35532 18172 35588
rect 18228 35532 18844 35588
rect 18900 35532 18910 35588
rect 8372 35476 8428 35532
rect 22876 35476 22932 35644
rect 50428 35588 50484 35644
rect 24210 35532 24220 35588
rect 24276 35532 25676 35588
rect 25732 35532 26908 35588
rect 27794 35532 27804 35588
rect 27860 35532 28924 35588
rect 28980 35532 28990 35588
rect 37426 35532 37436 35588
rect 37492 35532 39788 35588
rect 39844 35532 39854 35588
rect 44818 35532 44828 35588
rect 44884 35532 45612 35588
rect 45668 35532 46284 35588
rect 46340 35532 46350 35588
rect 48850 35532 48860 35588
rect 48916 35532 50484 35588
rect 50866 35532 50876 35588
rect 50932 35532 52780 35588
rect 52836 35532 55692 35588
rect 55748 35532 55758 35588
rect 26852 35476 26908 35532
rect 8372 35420 8876 35476
rect 8932 35420 8942 35476
rect 13122 35420 13132 35476
rect 13188 35420 22932 35476
rect 24546 35420 24556 35476
rect 24612 35420 25900 35476
rect 25956 35420 25966 35476
rect 26852 35420 33964 35476
rect 34020 35420 34524 35476
rect 34580 35420 34590 35476
rect 36418 35420 36428 35476
rect 36484 35420 37996 35476
rect 38052 35420 38062 35476
rect 39218 35420 39228 35476
rect 39284 35420 40236 35476
rect 40292 35420 41020 35476
rect 41076 35420 41086 35476
rect 42130 35420 42140 35476
rect 42196 35420 49196 35476
rect 49252 35420 49262 35476
rect 49410 35420 49420 35476
rect 49476 35420 55356 35476
rect 55412 35420 55422 35476
rect 1474 35308 1484 35364
rect 1540 35308 2156 35364
rect 2212 35308 2222 35364
rect 3826 35308 3836 35364
rect 3892 35308 5628 35364
rect 5684 35308 5694 35364
rect 10434 35308 10444 35364
rect 10500 35308 12124 35364
rect 12180 35308 12190 35364
rect 28466 35308 28476 35364
rect 28532 35308 29596 35364
rect 29652 35308 30156 35364
rect 30212 35308 32172 35364
rect 32228 35308 32238 35364
rect 37650 35308 37660 35364
rect 37716 35308 47628 35364
rect 47684 35308 47694 35364
rect 8355 35252 8365 35308
rect 8421 35252 8469 35308
rect 8525 35252 8573 35308
rect 8629 35252 8639 35308
rect 22662 35252 22672 35308
rect 22728 35252 22776 35308
rect 22832 35252 22880 35308
rect 22936 35252 22946 35308
rect 36969 35252 36979 35308
rect 37035 35252 37083 35308
rect 37139 35252 37187 35308
rect 37243 35252 37253 35308
rect 51276 35252 51286 35308
rect 51342 35252 51390 35308
rect 51446 35252 51494 35308
rect 51550 35252 51560 35308
rect 34290 35196 34300 35252
rect 34356 35196 35084 35252
rect 35140 35196 35150 35252
rect 38770 35196 38780 35252
rect 38836 35196 41132 35252
rect 41188 35196 41198 35252
rect 42802 35196 42812 35252
rect 42868 35196 47292 35252
rect 47348 35196 47358 35252
rect 56130 35196 56140 35252
rect 56196 35196 56700 35252
rect 56756 35196 56766 35252
rect 15922 35084 15932 35140
rect 15988 35084 22428 35140
rect 22484 35084 22494 35140
rect 23986 35084 23996 35140
rect 24052 35084 24444 35140
rect 24500 35084 35308 35140
rect 35364 35084 35374 35140
rect 47506 35084 47516 35140
rect 47572 35084 56588 35140
rect 56644 35084 56654 35140
rect 0 35028 800 35056
rect 0 34972 1708 35028
rect 1764 34972 1774 35028
rect 21410 34972 21420 35028
rect 21476 34972 21486 35028
rect 22306 34972 22316 35028
rect 22372 34972 25228 35028
rect 25284 34972 26348 35028
rect 26404 34972 26414 35028
rect 33730 34972 33740 35028
rect 33796 34972 36988 35028
rect 37044 34972 37054 35028
rect 37202 34972 37212 35028
rect 37268 34972 48972 35028
rect 49028 34972 49038 35028
rect 51202 34972 51212 35028
rect 51268 34972 52892 35028
rect 52948 34972 52958 35028
rect 56242 34972 56252 35028
rect 56308 34972 56318 35028
rect 0 34944 800 34972
rect 21420 34916 21476 34972
rect 1362 34860 1372 34916
rect 1428 34860 2268 34916
rect 2324 34860 2334 34916
rect 3490 34860 3500 34916
rect 3556 34860 3566 34916
rect 4050 34860 4060 34916
rect 4116 34860 5180 34916
rect 5236 34860 5246 34916
rect 21420 34860 21756 34916
rect 21812 34860 26460 34916
rect 26516 34860 26526 34916
rect 31714 34860 31724 34916
rect 31780 34860 42252 34916
rect 42308 34860 42924 34916
rect 42980 34860 42990 34916
rect 45490 34860 45500 34916
rect 45556 34860 47964 34916
rect 48020 34860 48030 34916
rect 55346 34860 55356 34916
rect 55412 34860 55692 34916
rect 55748 34860 55758 34916
rect 3500 34692 3556 34860
rect 56252 34804 56308 34972
rect 13010 34748 13020 34804
rect 13076 34748 14140 34804
rect 14196 34748 17556 34804
rect 17714 34748 17724 34804
rect 17780 34748 18732 34804
rect 18788 34748 18798 34804
rect 20290 34748 20300 34804
rect 20356 34748 21420 34804
rect 21476 34748 21486 34804
rect 22530 34748 22540 34804
rect 22596 34748 23436 34804
rect 23492 34748 23502 34804
rect 26852 34748 31836 34804
rect 31892 34748 31902 34804
rect 37874 34748 37884 34804
rect 37940 34748 38668 34804
rect 38770 34748 38780 34804
rect 38836 34748 39564 34804
rect 39620 34748 39630 34804
rect 43810 34748 43820 34804
rect 43876 34748 46844 34804
rect 46900 34748 46910 34804
rect 49858 34748 49868 34804
rect 49924 34748 51548 34804
rect 51604 34748 51614 34804
rect 56252 34748 56588 34804
rect 56644 34748 56654 34804
rect 2594 34636 2604 34692
rect 2660 34636 3388 34692
rect 3500 34636 9996 34692
rect 10052 34636 10062 34692
rect 3332 34468 3388 34636
rect 17500 34580 17556 34748
rect 17826 34636 17836 34692
rect 17892 34636 20524 34692
rect 20580 34636 21364 34692
rect 22418 34636 22428 34692
rect 22484 34636 24220 34692
rect 24276 34636 26124 34692
rect 26180 34636 26190 34692
rect 21308 34580 21364 34636
rect 26852 34580 26908 34748
rect 38612 34692 38668 34748
rect 32946 34636 32956 34692
rect 33012 34636 33852 34692
rect 33908 34636 33918 34692
rect 34178 34636 34188 34692
rect 34244 34636 36540 34692
rect 36596 34636 36606 34692
rect 38612 34636 39004 34692
rect 39060 34636 39070 34692
rect 45826 34636 45836 34692
rect 45892 34636 48188 34692
rect 48244 34636 48254 34692
rect 50642 34636 50652 34692
rect 50708 34636 50988 34692
rect 51044 34636 51660 34692
rect 51716 34636 55132 34692
rect 55188 34636 55198 34692
rect 17500 34524 18172 34580
rect 18228 34524 18238 34580
rect 19058 34524 19068 34580
rect 19124 34524 20972 34580
rect 21028 34524 21038 34580
rect 21298 34524 21308 34580
rect 21364 34524 26908 34580
rect 29334 34524 29372 34580
rect 29428 34524 29438 34580
rect 31602 34524 31612 34580
rect 31668 34524 38444 34580
rect 38500 34524 38510 34580
rect 15508 34468 15518 34524
rect 15574 34468 15622 34524
rect 15678 34468 15726 34524
rect 15782 34468 15792 34524
rect 29815 34468 29825 34524
rect 29881 34468 29929 34524
rect 29985 34468 30033 34524
rect 30089 34468 30099 34524
rect 44122 34468 44132 34524
rect 44188 34468 44236 34524
rect 44292 34468 44340 34524
rect 44396 34468 44406 34524
rect 58429 34468 58439 34524
rect 58495 34468 58543 34524
rect 58599 34468 58647 34524
rect 58703 34468 58713 34524
rect 3332 34412 11564 34468
rect 11620 34412 11630 34468
rect 49970 34412 49980 34468
rect 50036 34412 50540 34468
rect 50596 34412 50606 34468
rect 1810 34300 1820 34356
rect 1876 34300 6636 34356
rect 6692 34300 6702 34356
rect 8372 34300 11676 34356
rect 11732 34300 11742 34356
rect 11890 34300 11900 34356
rect 11956 34300 12796 34356
rect 12852 34300 12862 34356
rect 27570 34300 27580 34356
rect 27636 34300 29372 34356
rect 29428 34300 29438 34356
rect 29922 34300 29932 34356
rect 29988 34300 30940 34356
rect 30996 34300 31006 34356
rect 33506 34300 33516 34356
rect 33572 34300 34860 34356
rect 34916 34300 34926 34356
rect 35970 34300 35980 34356
rect 36036 34300 36764 34356
rect 36820 34300 36830 34356
rect 38612 34300 51884 34356
rect 51940 34300 51950 34356
rect 8372 34244 8428 34300
rect 3042 34188 3052 34244
rect 3108 34188 8428 34244
rect 9996 34188 19628 34244
rect 19684 34188 19694 34244
rect 22082 34188 22092 34244
rect 22148 34188 22540 34244
rect 22596 34188 22606 34244
rect 9996 34132 10052 34188
rect 38612 34132 38668 34300
rect 40002 34188 40012 34244
rect 40068 34188 41580 34244
rect 41636 34188 41646 34244
rect 2370 34076 2380 34132
rect 2436 34076 4396 34132
rect 4452 34076 4462 34132
rect 8194 34076 8204 34132
rect 8260 34076 10052 34132
rect 10210 34076 10220 34132
rect 10276 34076 18956 34132
rect 19012 34076 19022 34132
rect 25218 34076 25228 34132
rect 25284 34076 26012 34132
rect 26068 34076 31500 34132
rect 31556 34076 31566 34132
rect 32162 34076 32172 34132
rect 32228 34076 32956 34132
rect 33012 34076 33022 34132
rect 34188 34076 38668 34132
rect 39554 34076 39564 34132
rect 39620 34076 40124 34132
rect 40180 34076 41020 34132
rect 41076 34076 41086 34132
rect 47730 34076 47740 34132
rect 47796 34076 48748 34132
rect 48804 34076 48814 34132
rect 50530 34076 50540 34132
rect 50596 34076 51548 34132
rect 51604 34076 51614 34132
rect 53330 34076 53340 34132
rect 53396 34076 54572 34132
rect 54628 34076 55468 34132
rect 55524 34076 55534 34132
rect 55906 34076 55916 34132
rect 55972 34076 56700 34132
rect 56756 34076 56766 34132
rect 4620 33964 11116 34020
rect 11172 33964 12908 34020
rect 12964 33964 12974 34020
rect 23314 33964 23324 34020
rect 23380 33964 29876 34020
rect 32386 33964 32396 34020
rect 32452 33964 32732 34020
rect 32788 33964 33964 34020
rect 34020 33964 34030 34020
rect 0 33908 800 33936
rect 0 33852 1708 33908
rect 1764 33852 1774 33908
rect 2706 33852 2716 33908
rect 2772 33852 4060 33908
rect 4116 33852 4126 33908
rect 0 33824 800 33852
rect 4620 33796 4676 33964
rect 29820 33908 29876 33964
rect 18834 33852 18844 33908
rect 18900 33852 19516 33908
rect 19572 33852 20524 33908
rect 20580 33852 20590 33908
rect 22754 33852 22764 33908
rect 22820 33852 23996 33908
rect 24052 33852 25340 33908
rect 25396 33852 25406 33908
rect 25666 33852 25676 33908
rect 25732 33852 26908 33908
rect 26964 33852 26974 33908
rect 27570 33852 27580 33908
rect 27636 33852 28476 33908
rect 28532 33852 28542 33908
rect 29820 33852 32844 33908
rect 32900 33852 32910 33908
rect 34188 33796 34244 34076
rect 36194 33964 36204 34020
rect 36260 33964 36876 34020
rect 36932 33964 37324 34020
rect 37380 33964 40908 34020
rect 40964 33964 40974 34020
rect 35522 33852 35532 33908
rect 35588 33852 40012 33908
rect 40068 33852 40078 33908
rect 47954 33852 47964 33908
rect 48020 33852 51716 33908
rect 1138 33740 1148 33796
rect 1204 33740 3500 33796
rect 3556 33740 4620 33796
rect 4676 33740 4686 33796
rect 18274 33740 18284 33796
rect 18340 33740 19852 33796
rect 19908 33740 19918 33796
rect 24434 33740 24444 33796
rect 24500 33740 34244 33796
rect 37986 33740 37996 33796
rect 38052 33740 43820 33796
rect 43876 33740 43886 33796
rect 50530 33740 50540 33796
rect 50596 33740 50988 33796
rect 51044 33740 51054 33796
rect 8355 33684 8365 33740
rect 8421 33684 8469 33740
rect 8525 33684 8573 33740
rect 8629 33684 8639 33740
rect 22662 33684 22672 33740
rect 22728 33684 22776 33740
rect 22832 33684 22880 33740
rect 22936 33684 22946 33740
rect 36969 33684 36979 33740
rect 37035 33684 37083 33740
rect 37139 33684 37187 33740
rect 37243 33684 37253 33740
rect 51276 33684 51286 33740
rect 51342 33684 51390 33740
rect 51446 33684 51494 33740
rect 51550 33684 51560 33740
rect 11778 33628 11788 33684
rect 11844 33628 12572 33684
rect 12628 33628 21980 33684
rect 22036 33628 22046 33684
rect 27346 33628 27356 33684
rect 27412 33628 36428 33684
rect 36484 33628 36494 33684
rect 48850 33628 48860 33684
rect 48916 33628 50204 33684
rect 50260 33628 50270 33684
rect 51660 33572 51716 33852
rect 8866 33516 8876 33572
rect 8932 33516 47628 33572
rect 47684 33516 47694 33572
rect 50082 33516 50092 33572
rect 50148 33516 51212 33572
rect 51268 33516 51278 33572
rect 51538 33516 51548 33572
rect 51604 33516 51716 33572
rect 53218 33516 53228 33572
rect 53284 33516 54460 33572
rect 54516 33516 54526 33572
rect 1698 33404 1708 33460
rect 1764 33404 6188 33460
rect 6244 33404 6254 33460
rect 8194 33404 8204 33460
rect 8260 33404 9324 33460
rect 9380 33404 9390 33460
rect 9986 33404 9996 33460
rect 10052 33404 12012 33460
rect 12068 33404 12078 33460
rect 18722 33404 18732 33460
rect 18788 33404 20188 33460
rect 20244 33404 21980 33460
rect 22036 33404 27580 33460
rect 27636 33404 27646 33460
rect 28578 33404 28588 33460
rect 28644 33404 29596 33460
rect 29652 33404 29662 33460
rect 33282 33404 33292 33460
rect 33348 33404 34636 33460
rect 34692 33404 34702 33460
rect 34850 33404 34860 33460
rect 34916 33404 35420 33460
rect 35476 33404 35486 33460
rect 48748 33404 53116 33460
rect 53172 33404 53182 33460
rect 1810 33292 1820 33348
rect 1876 33292 3276 33348
rect 3332 33292 3342 33348
rect 4610 33292 4620 33348
rect 4676 33292 8540 33348
rect 8596 33292 8606 33348
rect 26852 33292 27244 33348
rect 27300 33292 27310 33348
rect 27682 33292 27692 33348
rect 27748 33292 28812 33348
rect 28868 33292 28878 33348
rect 29138 33292 29148 33348
rect 29204 33292 29484 33348
rect 29540 33292 29550 33348
rect 34962 33292 34972 33348
rect 35028 33292 35532 33348
rect 35588 33292 35598 33348
rect 36418 33292 36428 33348
rect 36484 33292 37100 33348
rect 37156 33292 37166 33348
rect 37426 33292 37436 33348
rect 37492 33292 38220 33348
rect 38276 33292 39452 33348
rect 39508 33292 39518 33348
rect 40226 33292 40236 33348
rect 40292 33292 41244 33348
rect 41300 33292 41310 33348
rect 43922 33292 43932 33348
rect 43988 33292 46284 33348
rect 46340 33292 46732 33348
rect 46788 33292 46798 33348
rect 46956 33292 47516 33348
rect 47572 33292 48188 33348
rect 48244 33292 48254 33348
rect 13010 33180 13020 33236
rect 13076 33180 13916 33236
rect 13972 33180 13982 33236
rect 26852 33124 26908 33292
rect 46956 33236 47012 33292
rect 48748 33236 48804 33404
rect 34514 33180 34524 33236
rect 34580 33180 35420 33236
rect 35476 33180 37548 33236
rect 37604 33180 37614 33236
rect 43698 33180 43708 33236
rect 43764 33180 47012 33236
rect 47282 33180 47292 33236
rect 47348 33180 48748 33236
rect 48804 33180 48814 33236
rect 49196 33180 50428 33236
rect 50484 33180 51324 33236
rect 51380 33180 52892 33236
rect 52948 33180 52958 33236
rect 49196 33124 49252 33180
rect 3042 33068 3052 33124
rect 3108 33068 7084 33124
rect 7140 33068 7150 33124
rect 19842 33068 19852 33124
rect 19908 33068 26572 33124
rect 26628 33068 26908 33124
rect 29362 33068 29372 33124
rect 29428 33068 30492 33124
rect 30548 33068 30940 33124
rect 30996 33068 38668 33124
rect 40786 33068 40796 33124
rect 40852 33068 41692 33124
rect 41748 33068 41758 33124
rect 47618 33068 47628 33124
rect 47684 33068 47694 33124
rect 48514 33068 48524 33124
rect 48580 33068 49252 33124
rect 50372 33068 51772 33124
rect 51828 33068 51838 33124
rect 38612 33012 38668 33068
rect 47628 33012 47684 33068
rect 50372 33012 50428 33068
rect 3714 32956 3724 33012
rect 3780 32956 7756 33012
rect 7812 32956 7822 33012
rect 19506 32956 19516 33012
rect 19572 32956 20188 33012
rect 20244 32956 21532 33012
rect 21588 32956 29652 33012
rect 30594 32956 30604 33012
rect 30660 32956 31836 33012
rect 31892 32956 32620 33012
rect 32676 32956 36988 33012
rect 37044 32956 37054 33012
rect 38612 32956 43764 33012
rect 47628 32956 50428 33012
rect 15508 32900 15518 32956
rect 15574 32900 15622 32956
rect 15678 32900 15726 32956
rect 15782 32900 15792 32956
rect 4162 32844 4172 32900
rect 4228 32844 6748 32900
rect 6804 32844 7196 32900
rect 7252 32844 7262 32900
rect 9202 32844 9212 32900
rect 9268 32844 10668 32900
rect 10724 32844 10734 32900
rect 16146 32844 16156 32900
rect 16212 32844 16828 32900
rect 16884 32844 16894 32900
rect 21858 32844 21868 32900
rect 21924 32844 23100 32900
rect 23156 32844 23884 32900
rect 23940 32844 23950 32900
rect 0 32788 800 32816
rect 29596 32788 29652 32956
rect 29815 32900 29825 32956
rect 29881 32900 29929 32956
rect 29985 32900 30033 32956
rect 30089 32900 30099 32956
rect 38770 32844 38780 32900
rect 38836 32844 40012 32900
rect 40068 32844 43372 32900
rect 43428 32844 43438 32900
rect 0 32732 1596 32788
rect 1652 32732 1662 32788
rect 9650 32732 9660 32788
rect 9716 32732 10332 32788
rect 10388 32732 10398 32788
rect 11778 32732 11788 32788
rect 11844 32732 18060 32788
rect 18116 32732 18126 32788
rect 21410 32732 21420 32788
rect 21476 32732 28028 32788
rect 28084 32732 28094 32788
rect 29596 32732 38892 32788
rect 38948 32732 38958 32788
rect 39106 32732 39116 32788
rect 39172 32732 39182 32788
rect 0 32704 800 32732
rect 39116 32676 39172 32732
rect 43708 32676 43764 32956
rect 44122 32900 44132 32956
rect 44188 32900 44236 32956
rect 44292 32900 44340 32956
rect 44396 32900 44406 32956
rect 58429 32900 58439 32956
rect 58495 32900 58543 32956
rect 58599 32900 58647 32956
rect 58703 32900 58713 32956
rect 43922 32732 43932 32788
rect 43988 32732 45164 32788
rect 45220 32732 45230 32788
rect 1810 32620 1820 32676
rect 1876 32620 3388 32676
rect 3444 32620 3454 32676
rect 6962 32620 6972 32676
rect 7028 32620 8316 32676
rect 8372 32620 10724 32676
rect 10668 32564 10724 32620
rect 15092 32620 16156 32676
rect 16212 32620 16222 32676
rect 21746 32620 21756 32676
rect 21812 32620 30380 32676
rect 30436 32620 30446 32676
rect 36306 32620 36316 32676
rect 36372 32620 38668 32676
rect 38724 32620 38734 32676
rect 39116 32620 39396 32676
rect 41906 32620 41916 32676
rect 41972 32620 41982 32676
rect 43708 32620 48748 32676
rect 48804 32620 48814 32676
rect 55906 32620 55916 32676
rect 55972 32620 58268 32676
rect 58324 32620 58334 32676
rect 15092 32564 15148 32620
rect 3938 32508 3948 32564
rect 4004 32508 6412 32564
rect 6468 32508 6478 32564
rect 8372 32508 9436 32564
rect 9492 32508 9502 32564
rect 10658 32508 10668 32564
rect 10724 32508 10734 32564
rect 14578 32508 14588 32564
rect 14644 32508 15148 32564
rect 15362 32508 15372 32564
rect 15428 32508 18508 32564
rect 18564 32508 18574 32564
rect 27122 32508 27132 32564
rect 27188 32508 30268 32564
rect 30324 32508 30334 32564
rect 30818 32508 30828 32564
rect 30884 32508 33180 32564
rect 33236 32508 33246 32564
rect 33506 32508 33516 32564
rect 33572 32508 34300 32564
rect 34356 32508 34366 32564
rect 38434 32508 38444 32564
rect 38500 32508 39116 32564
rect 39172 32508 39182 32564
rect 8372 32452 8428 32508
rect 30268 32452 30324 32508
rect 39340 32452 39396 32620
rect 41916 32564 41972 32620
rect 40338 32508 40348 32564
rect 40404 32508 41468 32564
rect 41524 32508 41972 32564
rect 43922 32508 43932 32564
rect 43988 32508 44828 32564
rect 44884 32508 44894 32564
rect 53106 32508 53116 32564
rect 53172 32508 54236 32564
rect 54292 32508 54302 32564
rect 5954 32396 5964 32452
rect 6020 32396 8428 32452
rect 9314 32396 9324 32452
rect 9380 32396 11452 32452
rect 11508 32396 11518 32452
rect 15138 32396 15148 32452
rect 15204 32396 16044 32452
rect 16100 32396 16110 32452
rect 18722 32396 18732 32452
rect 18788 32396 19516 32452
rect 19572 32396 19582 32452
rect 27682 32396 27692 32452
rect 27748 32396 28252 32452
rect 28308 32396 28318 32452
rect 30268 32396 31388 32452
rect 31444 32396 33292 32452
rect 33348 32396 33358 32452
rect 37762 32396 37772 32452
rect 37828 32396 38668 32452
rect 38724 32396 39396 32452
rect 41122 32396 41132 32452
rect 41188 32396 41804 32452
rect 41860 32396 41870 32452
rect 45378 32396 45388 32452
rect 45444 32396 50428 32452
rect 55122 32396 55132 32452
rect 55188 32396 57148 32452
rect 57204 32396 57214 32452
rect 50372 32340 50428 32396
rect 2258 32284 2268 32340
rect 2324 32284 4172 32340
rect 4228 32284 4238 32340
rect 7186 32284 7196 32340
rect 7252 32284 9212 32340
rect 9268 32284 9278 32340
rect 14690 32284 14700 32340
rect 14756 32284 15372 32340
rect 15428 32284 15438 32340
rect 15810 32284 15820 32340
rect 15876 32284 25676 32340
rect 25732 32284 25742 32340
rect 29138 32284 29148 32340
rect 29204 32284 29596 32340
rect 29652 32284 29662 32340
rect 38882 32284 38892 32340
rect 38948 32284 38958 32340
rect 41234 32284 41244 32340
rect 41300 32284 42028 32340
rect 42084 32284 42700 32340
rect 42756 32284 42766 32340
rect 50372 32284 54012 32340
rect 54068 32284 54078 32340
rect 38892 32228 38948 32284
rect 38892 32172 45724 32228
rect 45780 32172 45790 32228
rect 8355 32116 8365 32172
rect 8421 32116 8469 32172
rect 8525 32116 8573 32172
rect 8629 32116 8639 32172
rect 22662 32116 22672 32172
rect 22728 32116 22776 32172
rect 22832 32116 22880 32172
rect 22936 32116 22946 32172
rect 36969 32116 36979 32172
rect 37035 32116 37083 32172
rect 37139 32116 37187 32172
rect 37243 32116 37253 32172
rect 51276 32116 51286 32172
rect 51342 32116 51390 32172
rect 51446 32116 51494 32172
rect 51550 32116 51560 32172
rect 1586 32060 1596 32116
rect 1652 32060 3164 32116
rect 3220 32060 3230 32116
rect 15586 32060 15596 32116
rect 15652 32060 16268 32116
rect 16324 32060 16716 32116
rect 16772 32060 16782 32116
rect 37874 32060 37884 32116
rect 37940 32060 38780 32116
rect 38836 32060 39340 32116
rect 39396 32060 39406 32116
rect 42018 32060 42028 32116
rect 42084 32060 44044 32116
rect 44100 32060 44110 32116
rect 45612 32060 47180 32116
rect 47236 32060 47246 32116
rect 45612 32004 45668 32060
rect 2930 31948 2940 32004
rect 2996 31948 3836 32004
rect 3892 31948 5180 32004
rect 5236 31948 5246 32004
rect 7634 31948 7644 32004
rect 7700 31948 24332 32004
rect 24388 31948 24398 32004
rect 25666 31948 25676 32004
rect 25732 31948 26460 32004
rect 26516 31948 26526 32004
rect 26852 31948 27636 32004
rect 30146 31948 30156 32004
rect 30212 31948 45612 32004
rect 45668 31948 45678 32004
rect 46946 31948 46956 32004
rect 47012 31948 49308 32004
rect 49364 31948 49374 32004
rect 49522 31948 49532 32004
rect 49588 31948 50204 32004
rect 50260 31948 50876 32004
rect 50932 31948 53340 32004
rect 53396 31948 53406 32004
rect 26852 31892 26908 31948
rect 2818 31836 2828 31892
rect 2884 31836 3276 31892
rect 3332 31836 4620 31892
rect 4676 31836 4686 31892
rect 6514 31836 6524 31892
rect 6580 31836 7196 31892
rect 7252 31836 7262 31892
rect 7522 31836 7532 31892
rect 7588 31836 26908 31892
rect 27580 31780 27636 31948
rect 27906 31836 27916 31892
rect 27972 31836 33852 31892
rect 33908 31836 33918 31892
rect 34962 31836 34972 31892
rect 35028 31836 35812 31892
rect 36418 31836 36428 31892
rect 36484 31836 37772 31892
rect 37828 31836 39452 31892
rect 39508 31836 39518 31892
rect 41794 31836 41804 31892
rect 41860 31836 43708 31892
rect 43764 31836 43774 31892
rect 45490 31836 45500 31892
rect 45556 31836 46620 31892
rect 46676 31836 49084 31892
rect 49140 31836 49150 31892
rect 54898 31836 54908 31892
rect 54964 31836 55468 31892
rect 55524 31836 58156 31892
rect 58212 31836 58222 31892
rect 35756 31780 35812 31836
rect 1810 31724 1820 31780
rect 1876 31724 6076 31780
rect 6132 31724 6142 31780
rect 8418 31724 8428 31780
rect 8484 31724 10668 31780
rect 10724 31724 10734 31780
rect 13234 31724 13244 31780
rect 13300 31724 14252 31780
rect 14308 31724 16492 31780
rect 16548 31724 16558 31780
rect 17042 31724 17052 31780
rect 17108 31724 18284 31780
rect 18340 31724 18350 31780
rect 21522 31724 21532 31780
rect 21588 31724 26124 31780
rect 26180 31724 26190 31780
rect 26338 31724 26348 31780
rect 26404 31724 27356 31780
rect 27412 31724 27422 31780
rect 27580 31724 31724 31780
rect 31780 31724 31790 31780
rect 33282 31724 33292 31780
rect 33348 31724 33740 31780
rect 33796 31724 35532 31780
rect 35588 31724 35598 31780
rect 35756 31724 38780 31780
rect 38836 31724 38846 31780
rect 39666 31724 39676 31780
rect 39732 31724 39742 31780
rect 40562 31724 40572 31780
rect 40628 31724 45052 31780
rect 45108 31724 45118 31780
rect 45378 31724 45388 31780
rect 45444 31724 46284 31780
rect 46340 31724 48188 31780
rect 48244 31724 48860 31780
rect 48916 31724 48926 31780
rect 53554 31724 53564 31780
rect 53620 31724 56588 31780
rect 56644 31724 56654 31780
rect 56886 31724 56924 31780
rect 56980 31724 56990 31780
rect 0 31668 800 31696
rect 1820 31668 1876 31724
rect 0 31612 1876 31668
rect 3266 31612 3276 31668
rect 3332 31612 4732 31668
rect 4788 31612 5628 31668
rect 5684 31612 5694 31668
rect 8306 31612 8316 31668
rect 8372 31612 8988 31668
rect 9044 31612 9054 31668
rect 26852 31612 29148 31668
rect 29204 31612 29214 31668
rect 33394 31612 33404 31668
rect 33460 31612 34524 31668
rect 34580 31612 35980 31668
rect 36036 31612 36540 31668
rect 36596 31612 38892 31668
rect 38948 31612 38958 31668
rect 0 31584 800 31612
rect 5170 31500 5180 31556
rect 5236 31500 8876 31556
rect 8932 31500 10332 31556
rect 10388 31500 10398 31556
rect 10770 31500 10780 31556
rect 10836 31500 12908 31556
rect 12964 31500 12974 31556
rect 17938 31500 17948 31556
rect 18004 31500 18956 31556
rect 19012 31500 20188 31556
rect 20244 31500 20254 31556
rect 25666 31500 25676 31556
rect 25732 31500 26572 31556
rect 26628 31500 26638 31556
rect 26852 31444 26908 31612
rect 39676 31556 39732 31724
rect 41794 31612 41804 31668
rect 41860 31612 42588 31668
rect 42644 31612 42654 31668
rect 43138 31612 43148 31668
rect 43204 31612 46844 31668
rect 46900 31612 46910 31668
rect 27570 31500 27580 31556
rect 27636 31500 30212 31556
rect 31714 31500 31724 31556
rect 31780 31500 32508 31556
rect 32564 31500 32574 31556
rect 36642 31500 36652 31556
rect 36708 31500 38108 31556
rect 38164 31500 39732 31556
rect 17378 31388 17388 31444
rect 17444 31388 18060 31444
rect 18116 31388 20300 31444
rect 20356 31388 26908 31444
rect 15508 31332 15518 31388
rect 15574 31332 15622 31388
rect 15678 31332 15726 31388
rect 15782 31332 15792 31388
rect 27580 31220 27636 31500
rect 30156 31444 30212 31500
rect 30156 31388 34412 31444
rect 34468 31388 34478 31444
rect 29815 31332 29825 31388
rect 29881 31332 29929 31388
rect 29985 31332 30033 31388
rect 30089 31332 30099 31388
rect 44122 31332 44132 31388
rect 44188 31332 44236 31388
rect 44292 31332 44340 31388
rect 44396 31332 44406 31388
rect 58429 31332 58439 31388
rect 58495 31332 58543 31388
rect 58599 31332 58647 31388
rect 58703 31332 58713 31388
rect 2258 31164 2268 31220
rect 2324 31164 7980 31220
rect 8036 31164 8046 31220
rect 14802 31164 14812 31220
rect 14868 31164 15820 31220
rect 15876 31164 19012 31220
rect 19394 31164 19404 31220
rect 19460 31164 21644 31220
rect 21700 31164 21710 31220
rect 26674 31164 26684 31220
rect 26740 31164 27636 31220
rect 29362 31164 29372 31220
rect 29428 31164 31836 31220
rect 31892 31164 37548 31220
rect 37604 31164 37614 31220
rect 39218 31164 39228 31220
rect 39284 31164 40124 31220
rect 40180 31164 40908 31220
rect 40964 31164 40974 31220
rect 4946 31052 4956 31108
rect 5012 31052 6244 31108
rect 14914 31052 14924 31108
rect 14980 31052 16604 31108
rect 16660 31052 16670 31108
rect 6188 30996 6244 31052
rect 1698 30940 1708 30996
rect 1764 30940 5068 30996
rect 5124 30940 5134 30996
rect 6178 30940 6188 30996
rect 6244 30940 10108 30996
rect 10164 30940 10174 30996
rect 18956 30884 19012 31164
rect 26898 31052 26908 31108
rect 26964 31052 27692 31108
rect 27748 31052 27758 31108
rect 33282 31052 33292 31108
rect 33348 31052 36316 31108
rect 36372 31052 37324 31108
rect 37380 31052 37390 31108
rect 38612 31052 45948 31108
rect 46004 31052 46014 31108
rect 56914 31052 56924 31108
rect 56980 31052 58044 31108
rect 58100 31052 58110 31108
rect 23986 30940 23996 30996
rect 24052 30940 34076 30996
rect 34132 30940 34142 30996
rect 38612 30884 38668 31052
rect 42690 30940 42700 30996
rect 42756 30940 43932 30996
rect 43988 30940 43998 30996
rect 18956 30828 26908 30884
rect 28354 30828 28364 30884
rect 28420 30828 29372 30884
rect 29428 30828 29438 30884
rect 29810 30828 29820 30884
rect 29876 30828 30604 30884
rect 30660 30828 31500 30884
rect 31556 30828 38668 30884
rect 40338 30828 40348 30884
rect 40404 30828 41468 30884
rect 41524 30828 41534 30884
rect 48066 30828 48076 30884
rect 48132 30828 49308 30884
rect 49364 30828 49374 30884
rect 54450 30828 54460 30884
rect 54516 30828 55244 30884
rect 55300 30828 55310 30884
rect 26852 30772 26908 30828
rect 3154 30716 3164 30772
rect 3220 30716 4620 30772
rect 4676 30716 4686 30772
rect 20850 30716 20860 30772
rect 20916 30716 22428 30772
rect 22484 30716 22494 30772
rect 23314 30716 23324 30772
rect 23380 30716 24444 30772
rect 24500 30716 24510 30772
rect 26852 30716 28924 30772
rect 28980 30716 28990 30772
rect 32396 30660 32452 30828
rect 35186 30716 35196 30772
rect 35252 30716 41244 30772
rect 41300 30716 41310 30772
rect 44482 30716 44492 30772
rect 44548 30716 45500 30772
rect 45556 30716 45566 30772
rect 48178 30716 48188 30772
rect 48244 30716 50764 30772
rect 50820 30716 50830 30772
rect 23538 30604 23548 30660
rect 23604 30604 24556 30660
rect 24612 30604 24622 30660
rect 32386 30604 32396 30660
rect 32452 30604 32462 30660
rect 39330 30604 39340 30660
rect 39396 30604 43036 30660
rect 43092 30604 43102 30660
rect 0 30548 800 30576
rect 8355 30548 8365 30604
rect 8421 30548 8469 30604
rect 8525 30548 8573 30604
rect 8629 30548 8639 30604
rect 22662 30548 22672 30604
rect 22728 30548 22776 30604
rect 22832 30548 22880 30604
rect 22936 30548 22946 30604
rect 36969 30548 36979 30604
rect 37035 30548 37083 30604
rect 37139 30548 37187 30604
rect 37243 30548 37253 30604
rect 51276 30548 51286 30604
rect 51342 30548 51390 30604
rect 51446 30548 51494 30604
rect 51550 30548 51560 30604
rect 0 30492 1708 30548
rect 1764 30492 1774 30548
rect 2034 30492 2044 30548
rect 2100 30492 5180 30548
rect 5236 30492 5246 30548
rect 28242 30492 28252 30548
rect 28308 30492 29372 30548
rect 29428 30492 31836 30548
rect 31892 30492 31902 30548
rect 0 30464 800 30492
rect 2258 30380 2268 30436
rect 2324 30380 10332 30436
rect 10388 30380 10398 30436
rect 18610 30380 18620 30436
rect 18676 30380 19964 30436
rect 20020 30380 20030 30436
rect 28466 30380 28476 30436
rect 28532 30380 29484 30436
rect 29540 30380 30156 30436
rect 30212 30380 30222 30436
rect 44818 30380 44828 30436
rect 44884 30380 50652 30436
rect 50708 30380 50718 30436
rect 53666 30380 53676 30436
rect 53732 30380 57204 30436
rect 57148 30324 57204 30380
rect 2482 30268 2492 30324
rect 2548 30268 4956 30324
rect 5012 30268 5022 30324
rect 6738 30268 6748 30324
rect 6804 30268 8092 30324
rect 8148 30268 8158 30324
rect 18386 30268 18396 30324
rect 18452 30268 18900 30324
rect 21522 30268 21532 30324
rect 21588 30268 28420 30324
rect 31602 30268 31612 30324
rect 31668 30268 35980 30324
rect 36036 30268 36046 30324
rect 39788 30268 40292 30324
rect 41458 30268 41468 30324
rect 41524 30268 44604 30324
rect 44660 30268 44670 30324
rect 54450 30268 54460 30324
rect 54516 30268 56700 30324
rect 56756 30268 56766 30324
rect 57138 30268 57148 30324
rect 57204 30268 57214 30324
rect 18844 30212 18900 30268
rect 4498 30156 4508 30212
rect 4564 30156 5964 30212
rect 6020 30156 6030 30212
rect 9986 30156 9996 30212
rect 10052 30156 11340 30212
rect 11396 30156 11406 30212
rect 14914 30156 14924 30212
rect 14980 30156 17052 30212
rect 17108 30156 17118 30212
rect 18834 30156 18844 30212
rect 18900 30156 20188 30212
rect 20244 30156 20254 30212
rect 23538 30156 23548 30212
rect 23604 30156 26012 30212
rect 26068 30156 26078 30212
rect 28364 30100 28420 30268
rect 39788 30212 39844 30268
rect 28578 30156 28588 30212
rect 28644 30156 31388 30212
rect 31444 30156 31454 30212
rect 31938 30156 31948 30212
rect 32004 30156 39844 30212
rect 40002 30156 40012 30212
rect 40068 30156 40078 30212
rect 40012 30100 40068 30156
rect 1698 30044 1708 30100
rect 1764 30044 2492 30100
rect 2548 30044 2558 30100
rect 4722 30044 4732 30100
rect 4788 30044 6412 30100
rect 6468 30044 6478 30100
rect 8372 30044 10780 30100
rect 10836 30044 10846 30100
rect 15092 30044 26908 30100
rect 28364 30044 32060 30100
rect 32116 30044 32126 30100
rect 35522 30044 35532 30100
rect 35588 30044 36988 30100
rect 37044 30044 37054 30100
rect 37650 30044 37660 30100
rect 37716 30044 40068 30100
rect 40236 30100 40292 30268
rect 45714 30156 45724 30212
rect 45780 30156 47180 30212
rect 47236 30156 47246 30212
rect 49186 30156 49196 30212
rect 49252 30156 50428 30212
rect 50484 30156 50494 30212
rect 53778 30156 53788 30212
rect 53844 30156 55692 30212
rect 55748 30156 57372 30212
rect 57428 30156 57438 30212
rect 40236 30044 42812 30100
rect 42868 30044 42878 30100
rect 54114 30044 54124 30100
rect 54180 30044 55468 30100
rect 55524 30044 55534 30100
rect 55794 30044 55804 30100
rect 55860 30044 57596 30100
rect 57652 30044 57662 30100
rect 8372 29988 8428 30044
rect 2370 29932 2380 29988
rect 2436 29932 3052 29988
rect 3108 29932 3118 29988
rect 3938 29932 3948 29988
rect 4004 29932 8428 29988
rect 14700 29932 15036 29988
rect 15092 29932 15148 30044
rect 26852 29988 26908 30044
rect 37660 29988 37716 30044
rect 17042 29932 17052 29988
rect 17108 29932 17612 29988
rect 17668 29932 21868 29988
rect 21924 29932 21934 29988
rect 23986 29932 23996 29988
rect 24052 29932 24780 29988
rect 24836 29932 24846 29988
rect 26852 29932 29708 29988
rect 29764 29932 29774 29988
rect 37090 29932 37100 29988
rect 37156 29932 37716 29988
rect 42578 29932 42588 29988
rect 42644 29932 43484 29988
rect 43540 29932 52780 29988
rect 52836 29932 52846 29988
rect 52994 29932 53004 29988
rect 53060 29932 54236 29988
rect 54292 29932 54302 29988
rect 14700 29876 14756 29932
rect 3714 29820 3724 29876
rect 3780 29820 5516 29876
rect 5572 29820 5582 29876
rect 5730 29820 5740 29876
rect 5796 29820 7196 29876
rect 7252 29820 9660 29876
rect 9716 29820 9726 29876
rect 10210 29820 10220 29876
rect 10276 29820 11116 29876
rect 11172 29820 11182 29876
rect 14690 29820 14700 29876
rect 14756 29820 14766 29876
rect 18162 29820 18172 29876
rect 18228 29820 19404 29876
rect 19460 29820 19470 29876
rect 47954 29820 47964 29876
rect 48020 29820 48972 29876
rect 49028 29820 49038 29876
rect 5516 29652 5572 29820
rect 15508 29764 15518 29820
rect 15574 29764 15622 29820
rect 15678 29764 15726 29820
rect 15782 29764 15792 29820
rect 29815 29764 29825 29820
rect 29881 29764 29929 29820
rect 29985 29764 30033 29820
rect 30089 29764 30099 29820
rect 44122 29764 44132 29820
rect 44188 29764 44236 29820
rect 44292 29764 44340 29820
rect 44396 29764 44406 29820
rect 58429 29764 58439 29820
rect 58495 29764 58543 29820
rect 58599 29764 58647 29820
rect 58703 29764 58713 29820
rect 20850 29708 20860 29764
rect 20916 29708 21868 29764
rect 21924 29708 21934 29764
rect 28242 29708 28252 29764
rect 28308 29708 29596 29764
rect 29652 29708 29662 29764
rect 31938 29708 31948 29764
rect 32004 29708 33068 29764
rect 33124 29708 33134 29764
rect 5516 29596 8540 29652
rect 8596 29596 8606 29652
rect 12898 29596 12908 29652
rect 12964 29596 13804 29652
rect 13860 29596 20748 29652
rect 20804 29596 21196 29652
rect 21252 29596 21756 29652
rect 21812 29596 21822 29652
rect 24322 29596 24332 29652
rect 24388 29596 25676 29652
rect 25732 29596 25742 29652
rect 32386 29596 32396 29652
rect 32452 29596 32956 29652
rect 33012 29596 34636 29652
rect 34692 29596 34702 29652
rect 36194 29596 36204 29652
rect 36260 29596 36932 29652
rect 37762 29596 37772 29652
rect 37828 29596 38780 29652
rect 38836 29596 38846 29652
rect 42588 29596 44940 29652
rect 44996 29596 45500 29652
rect 45556 29596 45566 29652
rect 46386 29596 46396 29652
rect 46452 29596 48972 29652
rect 49028 29596 49038 29652
rect 56130 29596 56140 29652
rect 56196 29596 56924 29652
rect 56980 29596 56990 29652
rect 36876 29540 36932 29596
rect 42588 29540 42644 29596
rect 2930 29484 2940 29540
rect 2996 29484 9436 29540
rect 9492 29484 9502 29540
rect 15092 29484 36820 29540
rect 36876 29484 42644 29540
rect 42802 29484 42812 29540
rect 42868 29484 45724 29540
rect 45780 29484 45790 29540
rect 51650 29484 51660 29540
rect 51716 29484 54348 29540
rect 54404 29484 54414 29540
rect 55906 29484 55916 29540
rect 55972 29484 57932 29540
rect 57988 29484 57998 29540
rect 0 29428 800 29456
rect 15092 29428 15148 29484
rect 36764 29428 36820 29484
rect 0 29372 2380 29428
rect 2436 29372 2446 29428
rect 13346 29372 13356 29428
rect 13412 29372 15148 29428
rect 19730 29372 19740 29428
rect 19796 29372 23548 29428
rect 23604 29372 23772 29428
rect 23828 29372 23838 29428
rect 27570 29372 27580 29428
rect 27636 29372 29036 29428
rect 29092 29372 29102 29428
rect 30594 29372 30604 29428
rect 30660 29372 31612 29428
rect 31668 29372 31678 29428
rect 32162 29372 32172 29428
rect 32228 29372 33180 29428
rect 33236 29372 33246 29428
rect 35410 29372 35420 29428
rect 35476 29372 36540 29428
rect 36596 29372 36606 29428
rect 36764 29372 38668 29428
rect 44146 29372 44156 29428
rect 44212 29372 46284 29428
rect 46340 29372 46350 29428
rect 51762 29372 51772 29428
rect 51828 29372 53004 29428
rect 53060 29372 53228 29428
rect 53284 29372 54572 29428
rect 54628 29372 54638 29428
rect 0 29344 800 29372
rect 38612 29316 38668 29372
rect 1026 29260 1036 29316
rect 1092 29260 1932 29316
rect 1988 29260 5516 29316
rect 5572 29260 5582 29316
rect 7746 29260 7756 29316
rect 7812 29260 8204 29316
rect 8260 29260 8270 29316
rect 21298 29260 21308 29316
rect 21364 29260 22316 29316
rect 22372 29260 22382 29316
rect 24210 29260 24220 29316
rect 24276 29260 27916 29316
rect 27972 29260 27982 29316
rect 28802 29260 28812 29316
rect 28868 29260 29596 29316
rect 29652 29260 29662 29316
rect 35298 29260 35308 29316
rect 35364 29260 37324 29316
rect 37380 29260 37390 29316
rect 38612 29260 46060 29316
rect 46116 29260 46126 29316
rect 50306 29260 50316 29316
rect 50372 29260 51212 29316
rect 51268 29260 53340 29316
rect 53396 29260 54796 29316
rect 54852 29260 54862 29316
rect 2594 29148 2604 29204
rect 2660 29148 3052 29204
rect 3108 29148 3118 29204
rect 6076 29148 8316 29204
rect 8372 29148 9604 29204
rect 13010 29148 13020 29204
rect 13076 29148 13580 29204
rect 13636 29148 26908 29204
rect 33730 29148 33740 29204
rect 33796 29148 34524 29204
rect 34580 29148 34590 29204
rect 48178 29148 48188 29204
rect 48244 29148 49196 29204
rect 49252 29148 49532 29204
rect 49588 29148 49598 29204
rect 54002 29148 54012 29204
rect 54068 29148 55916 29204
rect 55972 29148 55982 29204
rect 6076 29092 6132 29148
rect 9548 29092 9604 29148
rect 26852 29092 26908 29148
rect 2118 29036 2156 29092
rect 2212 29036 2222 29092
rect 4946 29036 4956 29092
rect 5012 29036 6076 29092
rect 6132 29036 6142 29092
rect 9538 29036 9548 29092
rect 9604 29036 10108 29092
rect 10164 29036 10174 29092
rect 12786 29036 12796 29092
rect 12852 29036 13244 29092
rect 13300 29036 13310 29092
rect 23314 29036 23324 29092
rect 23380 29036 25116 29092
rect 25172 29036 25182 29092
rect 26852 29036 36820 29092
rect 53778 29036 53788 29092
rect 53844 29036 54236 29092
rect 54292 29036 54302 29092
rect 8355 28980 8365 29036
rect 8421 28980 8469 29036
rect 8525 28980 8573 29036
rect 8629 28980 8639 29036
rect 22662 28980 22672 29036
rect 22728 28980 22776 29036
rect 22832 28980 22880 29036
rect 22936 28980 22946 29036
rect 18162 28924 18172 28980
rect 18228 28924 19068 28980
rect 19124 28924 20076 28980
rect 20132 28924 20636 28980
rect 20692 28924 20702 28980
rect 23426 28924 23436 28980
rect 23492 28924 25900 28980
rect 25956 28924 27580 28980
rect 27636 28924 27646 28980
rect 31388 28924 36428 28980
rect 36484 28924 36494 28980
rect 31388 28868 31444 28924
rect 36764 28868 36820 29036
rect 36969 28980 36979 29036
rect 37035 28980 37083 29036
rect 37139 28980 37187 29036
rect 37243 28980 37253 29036
rect 51276 28980 51286 29036
rect 51342 28980 51390 29036
rect 51446 28980 51494 29036
rect 51550 28980 51560 29036
rect 41234 28924 41244 28980
rect 41300 28924 43596 28980
rect 43652 28924 43662 28980
rect 44034 28924 44044 28980
rect 44100 28924 44940 28980
rect 44996 28924 45006 28980
rect 1250 28812 1260 28868
rect 1316 28812 3724 28868
rect 3780 28812 3790 28868
rect 3938 28812 3948 28868
rect 4004 28812 4732 28868
rect 4788 28812 8316 28868
rect 8372 28812 8382 28868
rect 8642 28812 8652 28868
rect 8708 28812 31444 28868
rect 31602 28812 31612 28868
rect 31668 28812 34020 28868
rect 36764 28812 37100 28868
rect 37156 28812 37660 28868
rect 37716 28812 43372 28868
rect 43428 28812 44716 28868
rect 44772 28812 44782 28868
rect 49970 28812 49980 28868
rect 50036 28812 51548 28868
rect 51604 28812 52668 28868
rect 52724 28812 52734 28868
rect 54674 28812 54684 28868
rect 54740 28812 55692 28868
rect 55748 28812 57820 28868
rect 57876 28812 57886 28868
rect 10658 28700 10668 28756
rect 10724 28700 12796 28756
rect 12852 28700 12862 28756
rect 14466 28700 14476 28756
rect 14532 28700 20188 28756
rect 20244 28700 21476 28756
rect 21970 28700 21980 28756
rect 22036 28700 22988 28756
rect 23044 28700 24892 28756
rect 24948 28700 24958 28756
rect 25778 28700 25788 28756
rect 25844 28700 33292 28756
rect 33348 28700 33358 28756
rect 14476 28644 14532 28700
rect 3266 28588 3276 28644
rect 3332 28588 3724 28644
rect 3780 28588 3790 28644
rect 4722 28588 4732 28644
rect 4788 28588 5516 28644
rect 5572 28588 5582 28644
rect 5954 28588 5964 28644
rect 6020 28588 6748 28644
rect 6804 28588 6814 28644
rect 9426 28588 9436 28644
rect 9492 28588 9772 28644
rect 9828 28588 9838 28644
rect 11442 28588 11452 28644
rect 11508 28588 12012 28644
rect 12068 28588 12078 28644
rect 12226 28588 12236 28644
rect 12292 28588 14532 28644
rect 17714 28588 17724 28644
rect 17780 28588 18844 28644
rect 18900 28588 18910 28644
rect 3378 28476 3388 28532
rect 3444 28476 4396 28532
rect 4452 28476 4462 28532
rect 19730 28476 19740 28532
rect 19796 28476 20524 28532
rect 20580 28476 20590 28532
rect 21420 28420 21476 28700
rect 22530 28588 22540 28644
rect 22596 28588 23324 28644
rect 23380 28588 23390 28644
rect 23986 28588 23996 28644
rect 24052 28588 25452 28644
rect 25508 28588 25518 28644
rect 32946 28588 32956 28644
rect 33012 28588 33180 28644
rect 33236 28588 33740 28644
rect 33796 28588 33806 28644
rect 33964 28532 34020 28812
rect 35858 28700 35868 28756
rect 35924 28700 38668 28756
rect 39890 28700 39900 28756
rect 39956 28700 40796 28756
rect 40852 28700 40862 28756
rect 43922 28700 43932 28756
rect 43988 28700 45724 28756
rect 45780 28700 46396 28756
rect 46452 28700 46462 28756
rect 51874 28700 51884 28756
rect 51940 28700 52780 28756
rect 52836 28700 54012 28756
rect 54068 28700 54078 28756
rect 38612 28644 38668 28700
rect 38612 28588 39340 28644
rect 39396 28588 39406 28644
rect 39554 28588 39564 28644
rect 39620 28588 41580 28644
rect 41636 28588 41646 28644
rect 44258 28588 44268 28644
rect 44324 28588 45276 28644
rect 45332 28588 45342 28644
rect 51426 28588 51436 28644
rect 51492 28588 53228 28644
rect 53284 28588 53788 28644
rect 53844 28588 53854 28644
rect 55010 28588 55020 28644
rect 55076 28588 55804 28644
rect 55860 28588 56364 28644
rect 56420 28588 56430 28644
rect 22082 28476 22092 28532
rect 22148 28476 26908 28532
rect 26964 28476 26974 28532
rect 27122 28476 27132 28532
rect 27188 28476 28476 28532
rect 28532 28476 29260 28532
rect 29316 28476 29326 28532
rect 33964 28476 38668 28532
rect 40674 28476 40684 28532
rect 40740 28476 41244 28532
rect 41300 28476 41310 28532
rect 52098 28476 52108 28532
rect 52164 28476 54348 28532
rect 54404 28476 54414 28532
rect 56914 28476 56924 28532
rect 56980 28476 57372 28532
rect 57428 28476 58156 28532
rect 58212 28476 58222 28532
rect 1810 28364 1820 28420
rect 1876 28364 5292 28420
rect 5348 28364 5358 28420
rect 5842 28364 5852 28420
rect 5908 28364 11228 28420
rect 11284 28364 11294 28420
rect 11442 28364 11452 28420
rect 11508 28364 12124 28420
rect 12180 28364 12190 28420
rect 21410 28364 21420 28420
rect 21476 28364 22316 28420
rect 22372 28364 22382 28420
rect 24546 28364 24556 28420
rect 24612 28364 25788 28420
rect 25844 28364 25854 28420
rect 26852 28364 35756 28420
rect 35812 28364 36204 28420
rect 36260 28364 36270 28420
rect 37202 28364 37212 28420
rect 37268 28364 38220 28420
rect 38276 28364 38286 28420
rect 38612 28364 38668 28476
rect 38724 28364 38734 28420
rect 44818 28364 44828 28420
rect 44884 28364 45276 28420
rect 45332 28364 45342 28420
rect 0 28308 800 28336
rect 0 28252 1708 28308
rect 1764 28252 1774 28308
rect 0 28224 800 28252
rect 15508 28196 15518 28252
rect 15574 28196 15622 28252
rect 15678 28196 15726 28252
rect 15782 28196 15792 28252
rect 4050 28140 4060 28196
rect 4116 28140 4732 28196
rect 4788 28140 9324 28196
rect 9380 28140 9390 28196
rect 18498 28140 18508 28196
rect 18564 28140 23324 28196
rect 23380 28140 23390 28196
rect 10770 28028 10780 28084
rect 10836 28028 11900 28084
rect 11956 28028 11966 28084
rect 7298 27916 7308 27972
rect 7364 27916 13132 27972
rect 13188 27916 13198 27972
rect 18610 27916 18620 27972
rect 18676 27916 20188 27972
rect 20244 27916 20254 27972
rect 26852 27860 26908 28364
rect 45490 28252 45500 28308
rect 45556 28252 46284 28308
rect 46340 28252 46350 28308
rect 29815 28196 29825 28252
rect 29881 28196 29929 28252
rect 29985 28196 30033 28252
rect 30089 28196 30099 28252
rect 44122 28196 44132 28252
rect 44188 28196 44236 28252
rect 44292 28196 44340 28252
rect 44396 28196 44406 28252
rect 58429 28196 58439 28252
rect 58495 28196 58543 28252
rect 58599 28196 58647 28252
rect 58703 28196 58713 28252
rect 35410 28140 35420 28196
rect 35476 28140 35486 28196
rect 49298 28140 49308 28196
rect 49364 28140 52556 28196
rect 52612 28140 52622 28196
rect 35420 28084 35476 28140
rect 28802 28028 28812 28084
rect 28868 28028 35476 28084
rect 35532 28028 36316 28084
rect 36372 28028 36382 28084
rect 38770 28028 38780 28084
rect 38836 28028 41020 28084
rect 41076 28028 41086 28084
rect 51762 28028 51772 28084
rect 51828 28028 54236 28084
rect 54292 28028 54302 28084
rect 35532 27972 35588 28028
rect 27010 27916 27020 27972
rect 27076 27916 35588 27972
rect 35746 27916 35756 27972
rect 35812 27916 37212 27972
rect 37268 27916 37278 27972
rect 40226 27916 40236 27972
rect 40292 27916 40908 27972
rect 40964 27916 40974 27972
rect 41234 27916 41244 27972
rect 41300 27916 48132 27972
rect 50530 27916 50540 27972
rect 50596 27916 51884 27972
rect 51940 27916 51950 27972
rect 48076 27860 48132 27916
rect 8082 27804 8092 27860
rect 8148 27804 8428 27860
rect 8484 27804 8494 27860
rect 11442 27804 11452 27860
rect 11508 27804 13916 27860
rect 13972 27804 13982 27860
rect 18274 27804 18284 27860
rect 18340 27804 19404 27860
rect 19460 27804 19470 27860
rect 20066 27804 20076 27860
rect 20132 27804 20860 27860
rect 20916 27804 20926 27860
rect 21084 27804 26908 27860
rect 27346 27804 27356 27860
rect 27412 27804 27692 27860
rect 27748 27804 27758 27860
rect 34626 27804 34636 27860
rect 34692 27804 35644 27860
rect 35700 27804 38220 27860
rect 38276 27804 38286 27860
rect 43362 27804 43372 27860
rect 43428 27804 43820 27860
rect 43876 27804 43886 27860
rect 44258 27804 44268 27860
rect 44324 27804 45500 27860
rect 45556 27804 45566 27860
rect 45938 27804 45948 27860
rect 46004 27804 47852 27860
rect 47908 27804 47918 27860
rect 48066 27804 48076 27860
rect 48132 27804 48142 27860
rect 50306 27804 50316 27860
rect 50372 27804 50764 27860
rect 50820 27804 51436 27860
rect 51492 27804 51502 27860
rect 52994 27804 53004 27860
rect 53060 27804 55132 27860
rect 55188 27804 55198 27860
rect 14802 27692 14812 27748
rect 14868 27692 18956 27748
rect 19012 27692 19022 27748
rect 19842 27692 19852 27748
rect 19908 27692 20412 27748
rect 20468 27692 20478 27748
rect 21084 27636 21140 27804
rect 22306 27692 22316 27748
rect 22372 27692 22876 27748
rect 22932 27692 22942 27748
rect 24658 27692 24668 27748
rect 24724 27692 25228 27748
rect 25284 27692 25294 27748
rect 26002 27692 26012 27748
rect 26068 27692 28028 27748
rect 28084 27692 28094 27748
rect 28578 27692 28588 27748
rect 28644 27692 28654 27748
rect 31266 27692 31276 27748
rect 31332 27692 32172 27748
rect 32228 27692 42364 27748
rect 42420 27692 42430 27748
rect 43922 27692 43932 27748
rect 43988 27692 45052 27748
rect 45108 27692 45118 27748
rect 52098 27692 52108 27748
rect 52164 27692 52892 27748
rect 52948 27692 52958 27748
rect 53778 27692 53788 27748
rect 53844 27692 54572 27748
rect 54628 27692 54638 27748
rect 28588 27636 28644 27692
rect 14242 27580 14252 27636
rect 14308 27580 21140 27636
rect 22540 27580 25900 27636
rect 25956 27580 25966 27636
rect 26226 27580 26236 27636
rect 26292 27580 28644 27636
rect 34514 27580 34524 27636
rect 34580 27580 34590 27636
rect 34738 27580 34748 27636
rect 34804 27580 38668 27636
rect 43362 27580 43372 27636
rect 43428 27580 50204 27636
rect 50260 27580 50876 27636
rect 50932 27580 50942 27636
rect 51100 27580 52444 27636
rect 52500 27580 54796 27636
rect 54852 27580 54862 27636
rect 18050 27468 18060 27524
rect 18116 27468 22316 27524
rect 22372 27468 22382 27524
rect 8355 27412 8365 27468
rect 8421 27412 8469 27468
rect 8525 27412 8573 27468
rect 8629 27412 8639 27468
rect 22540 27412 22596 27580
rect 25442 27468 25452 27524
rect 25508 27468 27356 27524
rect 27412 27468 27422 27524
rect 28018 27468 28028 27524
rect 28084 27468 29372 27524
rect 29428 27468 29438 27524
rect 22662 27412 22672 27468
rect 22728 27412 22776 27468
rect 22832 27412 22880 27468
rect 22936 27412 22946 27468
rect 34524 27412 34580 27580
rect 38612 27524 38668 27580
rect 51100 27524 51156 27580
rect 38612 27468 45276 27524
rect 45332 27468 45342 27524
rect 46610 27468 46620 27524
rect 46676 27468 51156 27524
rect 36969 27412 36979 27468
rect 37035 27412 37083 27468
rect 37139 27412 37187 27468
rect 37243 27412 37253 27468
rect 51276 27412 51286 27468
rect 51342 27412 51390 27468
rect 51446 27412 51494 27468
rect 51550 27412 51560 27468
rect 19170 27356 19180 27412
rect 19236 27356 20300 27412
rect 20356 27356 20366 27412
rect 20524 27356 22596 27412
rect 23314 27356 23324 27412
rect 23380 27356 34860 27412
rect 34916 27356 34926 27412
rect 38612 27356 47516 27412
rect 47572 27356 47582 27412
rect 20524 27300 20580 27356
rect 38612 27300 38668 27356
rect 15698 27244 15708 27300
rect 15764 27244 20580 27300
rect 22082 27244 22092 27300
rect 22148 27244 22876 27300
rect 22932 27244 38668 27300
rect 46946 27244 46956 27300
rect 47012 27244 47740 27300
rect 47796 27244 47806 27300
rect 51874 27244 51884 27300
rect 51940 27244 52780 27300
rect 52836 27244 52846 27300
rect 55412 27244 57484 27300
rect 57540 27244 57550 27300
rect 0 27188 800 27216
rect 55412 27188 55468 27244
rect 0 27132 1820 27188
rect 1876 27132 1886 27188
rect 15922 27132 15932 27188
rect 15988 27132 17276 27188
rect 17332 27132 18172 27188
rect 18228 27132 18238 27188
rect 22194 27132 22204 27188
rect 22260 27132 22988 27188
rect 23044 27132 23054 27188
rect 23874 27132 23884 27188
rect 23940 27132 24892 27188
rect 24948 27132 24958 27188
rect 46834 27132 46844 27188
rect 46900 27132 47180 27188
rect 47236 27132 48412 27188
rect 48468 27132 48478 27188
rect 54786 27132 54796 27188
rect 54852 27132 55468 27188
rect 55804 27132 57316 27188
rect 0 27104 800 27132
rect 1820 27076 1876 27132
rect 55804 27076 55860 27132
rect 57260 27076 57316 27132
rect 1820 27020 2548 27076
rect 5282 27020 5292 27076
rect 5348 27020 5628 27076
rect 5684 27020 5694 27076
rect 11218 27020 11228 27076
rect 11284 27020 11788 27076
rect 11844 27020 11854 27076
rect 18610 27020 18620 27076
rect 18676 27020 19516 27076
rect 19572 27020 19582 27076
rect 22530 27020 22540 27076
rect 22596 27020 33740 27076
rect 33796 27020 34076 27076
rect 34132 27020 34142 27076
rect 38322 27020 38332 27076
rect 38388 27020 44940 27076
rect 44996 27020 45006 27076
rect 45490 27020 45500 27076
rect 45556 27020 45566 27076
rect 46274 27020 46284 27076
rect 46340 27020 47292 27076
rect 47348 27020 47852 27076
rect 47908 27020 47918 27076
rect 49298 27020 49308 27076
rect 49364 27020 49644 27076
rect 49700 27020 49710 27076
rect 52546 27020 52556 27076
rect 52612 27020 55860 27076
rect 56018 27020 56028 27076
rect 56084 27020 56094 27076
rect 57250 27020 57260 27076
rect 57316 27020 57326 27076
rect 2492 26740 2548 27020
rect 45500 26964 45556 27020
rect 56028 26964 56084 27020
rect 9202 26908 9212 26964
rect 9268 26908 9996 26964
rect 10052 26908 10332 26964
rect 10388 26908 10398 26964
rect 12002 26908 12012 26964
rect 12068 26908 12684 26964
rect 12740 26908 14028 26964
rect 14084 26908 14094 26964
rect 22642 26908 22652 26964
rect 22708 26908 23548 26964
rect 23604 26908 23614 26964
rect 24322 26908 24332 26964
rect 24388 26908 26236 26964
rect 26292 26908 26302 26964
rect 27906 26908 27916 26964
rect 27972 26908 29260 26964
rect 29316 26908 29326 26964
rect 30818 26908 30828 26964
rect 30884 26908 32060 26964
rect 32116 26908 32126 26964
rect 34962 26908 34972 26964
rect 35028 26908 35756 26964
rect 35812 26908 35822 26964
rect 42242 26908 42252 26964
rect 42308 26908 43260 26964
rect 43316 26908 43326 26964
rect 45500 26908 48188 26964
rect 48244 26908 48254 26964
rect 49522 26908 49532 26964
rect 49588 26908 50540 26964
rect 50596 26908 51884 26964
rect 51940 26908 51950 26964
rect 54114 26908 54124 26964
rect 54180 26908 56084 26964
rect 18834 26796 18844 26852
rect 18900 26796 19628 26852
rect 19684 26796 19694 26852
rect 20514 26796 20524 26852
rect 20580 26796 22316 26852
rect 22372 26796 22382 26852
rect 30034 26796 30044 26852
rect 30100 26796 38668 26852
rect 42018 26796 42028 26852
rect 42084 26796 43484 26852
rect 43540 26796 43550 26852
rect 50754 26796 50764 26852
rect 50820 26796 51548 26852
rect 51604 26796 51614 26852
rect 53890 26796 53900 26852
rect 53956 26796 57372 26852
rect 57428 26796 57438 26852
rect 2482 26684 2492 26740
rect 2548 26684 2558 26740
rect 15508 26628 15518 26684
rect 15574 26628 15622 26684
rect 15678 26628 15726 26684
rect 15782 26628 15792 26684
rect 29815 26628 29825 26684
rect 29881 26628 29929 26684
rect 29985 26628 30033 26684
rect 30089 26628 30099 26684
rect 7186 26572 7196 26628
rect 7252 26572 13468 26628
rect 13524 26572 13534 26628
rect 17938 26572 17948 26628
rect 18004 26572 20188 26628
rect 20244 26572 20748 26628
rect 20804 26572 20814 26628
rect 21858 26572 21868 26628
rect 21924 26572 22316 26628
rect 22372 26572 22382 26628
rect 23202 26572 23212 26628
rect 23268 26572 24892 26628
rect 24948 26572 25228 26628
rect 25284 26572 25294 26628
rect 33170 26572 33180 26628
rect 33236 26572 33964 26628
rect 34020 26572 34030 26628
rect 38612 26516 38668 26796
rect 44122 26628 44132 26684
rect 44188 26628 44236 26684
rect 44292 26628 44340 26684
rect 44396 26628 44406 26684
rect 58429 26628 58439 26684
rect 58495 26628 58543 26684
rect 58599 26628 58647 26684
rect 58703 26628 58713 26684
rect 47506 26572 47516 26628
rect 47572 26572 49308 26628
rect 49364 26572 49374 26628
rect 51650 26572 51660 26628
rect 51716 26572 51884 26628
rect 51940 26572 51950 26628
rect 53442 26572 53452 26628
rect 53508 26572 54012 26628
rect 54068 26572 55132 26628
rect 55188 26572 55198 26628
rect 7410 26460 7420 26516
rect 7476 26460 8988 26516
rect 9044 26460 9054 26516
rect 11974 26460 12012 26516
rect 12068 26460 12078 26516
rect 16370 26460 16380 26516
rect 16436 26460 26908 26516
rect 33282 26460 33292 26516
rect 33348 26460 33852 26516
rect 33908 26460 33918 26516
rect 34514 26460 34524 26516
rect 34580 26460 36204 26516
rect 36260 26460 37324 26516
rect 37380 26460 37390 26516
rect 38612 26460 56476 26516
rect 56532 26460 56542 26516
rect 26852 26404 26908 26460
rect 4610 26348 4620 26404
rect 4676 26348 7532 26404
rect 7588 26348 7598 26404
rect 26852 26348 30940 26404
rect 30996 26348 31006 26404
rect 33730 26348 33740 26404
rect 33796 26348 34300 26404
rect 34356 26348 34860 26404
rect 34916 26348 35308 26404
rect 35364 26348 35374 26404
rect 40114 26348 40124 26404
rect 40180 26348 41020 26404
rect 41076 26348 41086 26404
rect 44454 26348 44492 26404
rect 44548 26348 44558 26404
rect 46610 26348 46620 26404
rect 46676 26348 53340 26404
rect 53396 26348 54012 26404
rect 54068 26348 54078 26404
rect 3266 26236 3276 26292
rect 3332 26236 4676 26292
rect 4946 26236 4956 26292
rect 5012 26236 6076 26292
rect 6132 26236 6142 26292
rect 6514 26236 6524 26292
rect 6580 26236 8652 26292
rect 8708 26236 8718 26292
rect 19618 26236 19628 26292
rect 19684 26236 20300 26292
rect 20356 26236 20366 26292
rect 22866 26236 22876 26292
rect 22932 26236 23772 26292
rect 23828 26236 24220 26292
rect 24276 26236 24286 26292
rect 24658 26236 24668 26292
rect 24724 26236 25564 26292
rect 25620 26236 30492 26292
rect 30548 26236 30558 26292
rect 31602 26236 31612 26292
rect 31668 26236 32060 26292
rect 32116 26236 32284 26292
rect 32340 26236 32350 26292
rect 34962 26236 34972 26292
rect 35028 26236 37996 26292
rect 38052 26236 38332 26292
rect 38388 26236 38398 26292
rect 38546 26236 38556 26292
rect 38612 26236 40348 26292
rect 40404 26236 41132 26292
rect 41188 26236 41198 26292
rect 44594 26236 44604 26292
rect 44660 26236 45948 26292
rect 46004 26236 46014 26292
rect 49298 26236 49308 26292
rect 49364 26236 50428 26292
rect 50484 26236 50494 26292
rect 55906 26236 55916 26292
rect 55972 26236 57148 26292
rect 57204 26236 57214 26292
rect 0 25984 800 26096
rect 4620 26068 4676 26236
rect 8194 26124 8204 26180
rect 8260 26124 9772 26180
rect 9828 26124 10220 26180
rect 10276 26124 10286 26180
rect 15586 26124 15596 26180
rect 15652 26124 16492 26180
rect 16548 26124 17500 26180
rect 17556 26124 21532 26180
rect 21588 26124 21598 26180
rect 26852 26124 46956 26180
rect 47012 26124 47964 26180
rect 48020 26124 48030 26180
rect 52210 26124 52220 26180
rect 52276 26124 53228 26180
rect 53284 26124 54124 26180
rect 54180 26124 54190 26180
rect 55682 26124 55692 26180
rect 55748 26124 56700 26180
rect 56756 26124 56766 26180
rect 1474 26012 1484 26068
rect 1540 26012 4284 26068
rect 4340 26012 4350 26068
rect 4610 26012 4620 26068
rect 4676 26012 4686 26068
rect 26852 25956 26908 26124
rect 30482 26012 30492 26068
rect 30548 26012 47068 26068
rect 47124 26012 47134 26068
rect 24546 25900 24556 25956
rect 24612 25900 26908 25956
rect 37874 25900 37884 25956
rect 37940 25900 37996 25956
rect 38052 25900 38062 25956
rect 38210 25900 38220 25956
rect 38276 25900 38314 25956
rect 39106 25900 39116 25956
rect 39172 25900 50204 25956
rect 50260 25900 50270 25956
rect 8355 25844 8365 25900
rect 8421 25844 8469 25900
rect 8525 25844 8573 25900
rect 8629 25844 8639 25900
rect 22662 25844 22672 25900
rect 22728 25844 22776 25900
rect 22832 25844 22880 25900
rect 22936 25844 22946 25900
rect 36969 25844 36979 25900
rect 37035 25844 37083 25900
rect 37139 25844 37187 25900
rect 37243 25844 37253 25900
rect 51276 25844 51286 25900
rect 51342 25844 51390 25900
rect 51446 25844 51494 25900
rect 51550 25844 51560 25900
rect 21522 25788 21532 25844
rect 21588 25788 22428 25844
rect 22484 25788 22494 25844
rect 23090 25788 23100 25844
rect 23156 25788 32844 25844
rect 32900 25788 33180 25844
rect 33236 25788 33246 25844
rect 37874 25788 37884 25844
rect 37940 25788 38332 25844
rect 38388 25788 38398 25844
rect 2034 25676 2044 25732
rect 2100 25676 6188 25732
rect 6244 25676 6254 25732
rect 8530 25676 8540 25732
rect 8596 25676 13356 25732
rect 13412 25676 13422 25732
rect 13682 25676 13692 25732
rect 13748 25676 14364 25732
rect 14420 25676 26908 25732
rect 28130 25676 28140 25732
rect 28196 25676 28588 25732
rect 28644 25676 28654 25732
rect 36082 25676 36092 25732
rect 36148 25676 36988 25732
rect 37044 25676 37054 25732
rect 37314 25676 37324 25732
rect 37380 25676 38108 25732
rect 38164 25676 39340 25732
rect 39396 25676 39406 25732
rect 43586 25676 43596 25732
rect 43652 25676 43932 25732
rect 43988 25676 43998 25732
rect 48178 25676 48188 25732
rect 48244 25676 49084 25732
rect 49140 25676 49150 25732
rect 51202 25676 51212 25732
rect 51268 25676 51772 25732
rect 51828 25676 52780 25732
rect 52836 25676 52846 25732
rect 26852 25620 26908 25676
rect 4050 25564 4060 25620
rect 4116 25564 4844 25620
rect 4900 25564 8204 25620
rect 8260 25564 8270 25620
rect 11890 25564 11900 25620
rect 11956 25564 12460 25620
rect 12516 25564 12526 25620
rect 16370 25564 16380 25620
rect 16436 25564 17164 25620
rect 17220 25564 24556 25620
rect 24612 25564 24622 25620
rect 26852 25564 39116 25620
rect 39172 25564 39182 25620
rect 46162 25564 46172 25620
rect 46228 25564 47068 25620
rect 47124 25564 47134 25620
rect 47292 25564 51548 25620
rect 51604 25564 52892 25620
rect 52948 25564 52958 25620
rect 55906 25564 55916 25620
rect 55972 25564 57596 25620
rect 57652 25564 57662 25620
rect 47292 25508 47348 25564
rect 2034 25452 2044 25508
rect 2100 25452 10052 25508
rect 11974 25452 12012 25508
rect 12068 25452 12078 25508
rect 15026 25452 15036 25508
rect 15092 25452 15820 25508
rect 15876 25452 21308 25508
rect 21364 25452 25228 25508
rect 25284 25452 25294 25508
rect 27906 25452 27916 25508
rect 27972 25452 29148 25508
rect 29204 25452 29214 25508
rect 30146 25452 30156 25508
rect 30212 25452 30716 25508
rect 30772 25452 30782 25508
rect 31154 25452 31164 25508
rect 31220 25452 32172 25508
rect 32228 25452 32238 25508
rect 34850 25452 34860 25508
rect 34916 25452 35868 25508
rect 35924 25452 37772 25508
rect 37828 25452 38332 25508
rect 38388 25452 38398 25508
rect 38546 25452 38556 25508
rect 38612 25452 39452 25508
rect 39508 25452 40012 25508
rect 40068 25452 40078 25508
rect 43586 25452 43596 25508
rect 43652 25452 47348 25508
rect 47842 25452 47852 25508
rect 47908 25452 48636 25508
rect 48692 25452 48702 25508
rect 52108 25452 53340 25508
rect 53396 25452 53406 25508
rect 55122 25452 55132 25508
rect 55188 25452 55804 25508
rect 55860 25452 55870 25508
rect 9996 25284 10052 25452
rect 11218 25340 11228 25396
rect 11284 25340 11676 25396
rect 11732 25340 11742 25396
rect 16706 25340 16716 25396
rect 16772 25340 20524 25396
rect 20580 25340 21644 25396
rect 21700 25340 21710 25396
rect 22418 25340 22428 25396
rect 22484 25340 25788 25396
rect 25844 25340 25854 25396
rect 27570 25340 27580 25396
rect 27636 25340 27804 25396
rect 27860 25340 30268 25396
rect 30324 25340 30334 25396
rect 33170 25340 33180 25396
rect 33236 25340 34972 25396
rect 35028 25340 35038 25396
rect 37314 25340 37324 25396
rect 37380 25340 37548 25396
rect 37604 25340 37614 25396
rect 38322 25340 38332 25396
rect 38388 25340 39788 25396
rect 39844 25340 39854 25396
rect 45938 25340 45948 25396
rect 46004 25340 46508 25396
rect 46564 25340 46574 25396
rect 52108 25284 52164 25452
rect 53442 25340 53452 25396
rect 53508 25340 54236 25396
rect 54292 25340 54302 25396
rect 9986 25228 9996 25284
rect 10052 25228 10444 25284
rect 10500 25228 12796 25284
rect 12852 25228 12862 25284
rect 14018 25228 14028 25284
rect 14084 25228 23100 25284
rect 23156 25228 23166 25284
rect 27122 25228 27132 25284
rect 27188 25228 27916 25284
rect 27972 25228 30044 25284
rect 30100 25228 30110 25284
rect 32946 25228 32956 25284
rect 33012 25228 34412 25284
rect 34468 25228 34478 25284
rect 35970 25228 35980 25284
rect 36036 25228 37100 25284
rect 37156 25228 37548 25284
rect 37604 25228 37614 25284
rect 49186 25228 49196 25284
rect 49252 25228 52108 25284
rect 52164 25228 52174 25284
rect 53330 25228 53340 25284
rect 53396 25228 54124 25284
rect 54180 25228 54190 25284
rect 3378 25116 3388 25172
rect 3444 25116 3948 25172
rect 4004 25116 4014 25172
rect 16258 25116 16268 25172
rect 16324 25116 22876 25172
rect 22932 25116 22942 25172
rect 28802 25116 28812 25172
rect 28868 25116 29596 25172
rect 29652 25116 29662 25172
rect 30594 25116 30604 25172
rect 30660 25116 33852 25172
rect 33908 25116 33918 25172
rect 35634 25116 35644 25172
rect 35700 25116 36428 25172
rect 36484 25116 36494 25172
rect 40562 25116 40572 25172
rect 40628 25116 42476 25172
rect 42532 25116 42542 25172
rect 15508 25060 15518 25116
rect 15574 25060 15622 25116
rect 15678 25060 15726 25116
rect 15782 25060 15792 25116
rect 29815 25060 29825 25116
rect 29881 25060 29929 25116
rect 29985 25060 30033 25116
rect 30089 25060 30099 25116
rect 17500 25004 22316 25060
rect 22372 25004 22382 25060
rect 29138 25004 29148 25060
rect 29204 25004 29372 25060
rect 29428 25004 29438 25060
rect 0 24864 800 24976
rect 17500 24948 17556 25004
rect 33852 24948 33908 25116
rect 44122 25060 44132 25116
rect 44188 25060 44236 25116
rect 44292 25060 44340 25116
rect 44396 25060 44406 25116
rect 58429 25060 58439 25116
rect 58495 25060 58543 25116
rect 58599 25060 58647 25116
rect 58703 25060 58713 25116
rect 34066 25004 34076 25060
rect 34132 25004 41916 25060
rect 41972 25004 41982 25060
rect 2146 24892 2156 24948
rect 2212 24892 5796 24948
rect 15474 24892 15484 24948
rect 15540 24892 17556 24948
rect 18274 24892 18284 24948
rect 18340 24892 19180 24948
rect 19236 24892 19246 24948
rect 21970 24892 21980 24948
rect 22036 24892 24332 24948
rect 24388 24892 24398 24948
rect 27682 24892 27692 24948
rect 27748 24892 28476 24948
rect 28532 24892 33628 24948
rect 33684 24892 33694 24948
rect 33852 24892 36764 24948
rect 36820 24892 36830 24948
rect 37538 24892 37548 24948
rect 37604 24892 38892 24948
rect 38948 24892 43092 24948
rect 43922 24892 43932 24948
rect 43988 24892 45276 24948
rect 45332 24892 45836 24948
rect 45892 24892 45902 24948
rect 46610 24892 46620 24948
rect 46676 24892 48188 24948
rect 48244 24892 48254 24948
rect 50418 24892 50428 24948
rect 50484 24892 51548 24948
rect 51604 24892 51614 24948
rect 3164 24780 4060 24836
rect 4116 24780 4126 24836
rect 3164 24724 3220 24780
rect 5740 24724 5796 24892
rect 43036 24836 43092 24892
rect 8306 24780 8316 24836
rect 8372 24780 27020 24836
rect 27076 24780 27086 24836
rect 27570 24780 27580 24836
rect 27636 24780 30492 24836
rect 30548 24780 30558 24836
rect 31500 24780 37884 24836
rect 37940 24780 37950 24836
rect 38098 24780 38108 24836
rect 38164 24780 39228 24836
rect 39284 24780 39294 24836
rect 41906 24780 41916 24836
rect 41972 24780 42812 24836
rect 42868 24780 42878 24836
rect 43036 24780 49420 24836
rect 49476 24780 49486 24836
rect 50530 24780 50540 24836
rect 50596 24780 52220 24836
rect 52276 24780 52286 24836
rect 3154 24668 3164 24724
rect 3220 24668 3230 24724
rect 3938 24668 3948 24724
rect 4004 24668 4396 24724
rect 4452 24668 4462 24724
rect 5730 24668 5740 24724
rect 5796 24668 5806 24724
rect 15092 24668 15484 24724
rect 15540 24668 15550 24724
rect 19618 24668 19628 24724
rect 19684 24668 23772 24724
rect 23828 24668 23838 24724
rect 28018 24668 28028 24724
rect 28084 24668 29260 24724
rect 29316 24668 29326 24724
rect 29698 24668 29708 24724
rect 29764 24668 30940 24724
rect 30996 24668 31006 24724
rect 3276 24556 3388 24612
rect 3444 24556 3454 24612
rect 7634 24556 7644 24612
rect 7700 24556 8092 24612
rect 8148 24556 8652 24612
rect 8708 24556 8718 24612
rect 15026 24556 15036 24612
rect 15092 24556 15148 24668
rect 31500 24612 31556 24780
rect 32162 24668 32172 24724
rect 32228 24668 33404 24724
rect 33460 24668 33470 24724
rect 37090 24668 37100 24724
rect 37156 24668 38444 24724
rect 38500 24668 38510 24724
rect 38612 24668 38892 24724
rect 38948 24668 38958 24724
rect 41234 24668 41244 24724
rect 41300 24668 42924 24724
rect 42980 24668 42990 24724
rect 44034 24668 44044 24724
rect 44100 24668 44492 24724
rect 44548 24668 44558 24724
rect 45042 24668 45052 24724
rect 45108 24668 46060 24724
rect 46116 24668 46396 24724
rect 46452 24668 46956 24724
rect 47012 24668 47022 24724
rect 50418 24668 50428 24724
rect 50484 24668 52556 24724
rect 52612 24668 52622 24724
rect 53106 24668 53116 24724
rect 53172 24668 54684 24724
rect 54740 24668 54750 24724
rect 24658 24556 24668 24612
rect 24724 24556 25340 24612
rect 25396 24556 26124 24612
rect 26180 24556 26190 24612
rect 30706 24556 30716 24612
rect 30772 24556 31500 24612
rect 31556 24556 31566 24612
rect 36194 24556 36204 24612
rect 36260 24556 37548 24612
rect 37604 24556 37614 24612
rect 38070 24556 38108 24612
rect 38164 24556 38174 24612
rect 3276 24500 3332 24556
rect 38612 24500 38668 24668
rect 38770 24556 38780 24612
rect 38836 24556 40012 24612
rect 40068 24556 40078 24612
rect 2482 24444 2492 24500
rect 2548 24444 3332 24500
rect 4050 24444 4060 24500
rect 4116 24444 6412 24500
rect 6468 24444 6478 24500
rect 18274 24444 18284 24500
rect 18340 24444 19740 24500
rect 19796 24444 25004 24500
rect 25060 24444 25070 24500
rect 29810 24444 29820 24500
rect 29876 24444 30268 24500
rect 30324 24444 38668 24500
rect 44492 24500 44548 24668
rect 47618 24556 47628 24612
rect 47684 24556 49084 24612
rect 49140 24556 49150 24612
rect 57250 24556 57260 24612
rect 57316 24556 58156 24612
rect 58212 24556 58222 24612
rect 44492 24444 45052 24500
rect 45108 24444 45118 24500
rect 54674 24444 54684 24500
rect 54740 24444 56924 24500
rect 56980 24444 56990 24500
rect 38182 24332 38220 24388
rect 38276 24332 38286 24388
rect 38892 24332 43932 24388
rect 43988 24332 44716 24388
rect 44772 24332 44782 24388
rect 8355 24276 8365 24332
rect 8421 24276 8469 24332
rect 8525 24276 8573 24332
rect 8629 24276 8639 24332
rect 22662 24276 22672 24332
rect 22728 24276 22776 24332
rect 22832 24276 22880 24332
rect 22936 24276 22946 24332
rect 36969 24276 36979 24332
rect 37035 24276 37083 24332
rect 37139 24276 37187 24332
rect 37243 24276 37253 24332
rect 38892 24276 38948 24332
rect 51276 24276 51286 24332
rect 51342 24276 51390 24332
rect 51446 24276 51494 24332
rect 51550 24276 51560 24332
rect 1698 24220 1708 24276
rect 1764 24220 3276 24276
rect 3332 24220 3342 24276
rect 10994 24220 11004 24276
rect 11060 24220 13468 24276
rect 13524 24220 13534 24276
rect 23202 24220 23212 24276
rect 23268 24220 31948 24276
rect 32004 24220 32014 24276
rect 37874 24220 37884 24276
rect 37940 24220 38948 24276
rect 39106 24220 39116 24276
rect 39172 24220 49756 24276
rect 49812 24220 49822 24276
rect 2258 24108 2268 24164
rect 2324 24108 3164 24164
rect 3220 24108 3230 24164
rect 6290 24108 6300 24164
rect 6356 24108 7532 24164
rect 7588 24108 7598 24164
rect 10210 24108 10220 24164
rect 10276 24108 11116 24164
rect 11172 24108 11182 24164
rect 13346 24108 13356 24164
rect 13412 24108 35644 24164
rect 35700 24108 46508 24164
rect 46564 24108 46574 24164
rect 47618 24108 47628 24164
rect 47684 24108 48636 24164
rect 48692 24108 49308 24164
rect 49364 24108 49374 24164
rect 51986 24108 51996 24164
rect 52052 24108 53116 24164
rect 53172 24108 53182 24164
rect 2156 23996 4620 24052
rect 4676 23996 4686 24052
rect 17714 23996 17724 24052
rect 17780 23996 18508 24052
rect 18564 23996 18574 24052
rect 19618 23996 19628 24052
rect 19684 23996 21420 24052
rect 21476 23996 21486 24052
rect 27010 23996 27020 24052
rect 27076 23996 27580 24052
rect 27636 23996 27646 24052
rect 36082 23996 36092 24052
rect 36148 23996 37548 24052
rect 37604 23996 37614 24052
rect 37986 23996 37996 24052
rect 38052 23996 38444 24052
rect 38500 23996 38510 24052
rect 43586 23996 43596 24052
rect 43652 23996 43932 24052
rect 43988 23996 43998 24052
rect 44828 23996 45164 24052
rect 45220 23996 45230 24052
rect 0 23744 800 23856
rect 2156 23716 2212 23996
rect 44828 23940 44884 23996
rect 46508 23940 46564 24108
rect 50418 23996 50428 24052
rect 50484 23996 53340 24052
rect 53396 23996 53406 24052
rect 7634 23884 7644 23940
rect 7700 23884 8204 23940
rect 8260 23884 8270 23940
rect 21074 23884 21084 23940
rect 21140 23884 23212 23940
rect 23268 23884 23278 23940
rect 28578 23884 28588 23940
rect 28644 23884 29596 23940
rect 29652 23884 31724 23940
rect 31780 23884 31892 23940
rect 32386 23884 32396 23940
rect 32452 23884 32956 23940
rect 33012 23884 35308 23940
rect 35364 23884 35374 23940
rect 38546 23884 38556 23940
rect 38612 23884 39900 23940
rect 39956 23884 39966 23940
rect 43698 23884 43708 23940
rect 43764 23884 44884 23940
rect 45042 23884 45052 23940
rect 45108 23884 45836 23940
rect 45892 23884 45902 23940
rect 46508 23884 50596 23940
rect 2604 23772 3388 23828
rect 3444 23772 3454 23828
rect 6962 23772 6972 23828
rect 7028 23772 7868 23828
rect 7924 23772 7934 23828
rect 11890 23772 11900 23828
rect 11956 23772 12012 23828
rect 12068 23772 12572 23828
rect 12628 23772 12638 23828
rect 21410 23772 21420 23828
rect 21476 23772 28812 23828
rect 28868 23772 28878 23828
rect 2146 23660 2156 23716
rect 2212 23660 2222 23716
rect 2604 23604 2660 23772
rect 31836 23716 31892 23884
rect 32050 23772 32060 23828
rect 32116 23772 33068 23828
rect 33124 23772 33134 23828
rect 35858 23772 35868 23828
rect 35924 23772 37100 23828
rect 37156 23772 39004 23828
rect 39060 23772 46900 23828
rect 47394 23772 47404 23828
rect 47460 23772 48356 23828
rect 46844 23716 46900 23772
rect 48300 23716 48356 23772
rect 50540 23716 50596 23884
rect 51314 23772 51324 23828
rect 51380 23772 52892 23828
rect 52948 23772 52958 23828
rect 56242 23772 56252 23828
rect 56308 23772 57036 23828
rect 57092 23772 57102 23828
rect 2818 23660 2828 23716
rect 2884 23660 4508 23716
rect 4564 23660 4574 23716
rect 12002 23660 12012 23716
rect 12068 23660 12124 23716
rect 12180 23660 12190 23716
rect 17378 23660 17388 23716
rect 17444 23660 19740 23716
rect 19796 23660 19806 23716
rect 20290 23660 20300 23716
rect 20356 23660 21308 23716
rect 21364 23660 21374 23716
rect 24546 23660 24556 23716
rect 24612 23660 25228 23716
rect 25284 23660 25294 23716
rect 26852 23660 27692 23716
rect 27748 23660 27758 23716
rect 28018 23660 28028 23716
rect 28084 23660 31388 23716
rect 31444 23660 31454 23716
rect 31836 23660 32284 23716
rect 32340 23660 32350 23716
rect 37510 23660 37548 23716
rect 37604 23660 37614 23716
rect 37958 23660 37996 23716
rect 38052 23660 38062 23716
rect 39778 23660 39788 23716
rect 39844 23660 42700 23716
rect 42756 23660 44548 23716
rect 44706 23660 44716 23716
rect 44772 23660 45948 23716
rect 46004 23660 46014 23716
rect 46834 23660 46844 23716
rect 46900 23660 47964 23716
rect 48020 23660 48030 23716
rect 48290 23660 48300 23716
rect 48356 23660 49868 23716
rect 49924 23660 49934 23716
rect 50082 23660 50092 23716
rect 50148 23660 50428 23716
rect 50530 23660 50540 23716
rect 50596 23660 50634 23716
rect 50754 23660 50764 23716
rect 50820 23660 51548 23716
rect 51604 23660 52780 23716
rect 52836 23660 52846 23716
rect 56466 23660 56476 23716
rect 56532 23660 57260 23716
rect 57316 23660 57326 23716
rect 26852 23604 26908 23660
rect 44492 23604 44548 23660
rect 50372 23604 50428 23660
rect 2258 23548 2268 23604
rect 2324 23548 2604 23604
rect 2660 23548 2670 23604
rect 24434 23548 24444 23604
rect 24500 23548 26908 23604
rect 27906 23548 27916 23604
rect 27972 23548 29260 23604
rect 29316 23548 29326 23604
rect 39666 23548 39676 23604
rect 39732 23548 40908 23604
rect 40964 23548 41692 23604
rect 41748 23548 41758 23604
rect 44492 23548 45724 23604
rect 45780 23548 49756 23604
rect 49812 23548 49822 23604
rect 50372 23548 51324 23604
rect 51380 23548 51390 23604
rect 15508 23492 15518 23548
rect 15574 23492 15622 23548
rect 15678 23492 15726 23548
rect 15782 23492 15792 23548
rect 29815 23492 29825 23548
rect 29881 23492 29929 23548
rect 29985 23492 30033 23548
rect 30089 23492 30099 23548
rect 44122 23492 44132 23548
rect 44188 23492 44236 23548
rect 44292 23492 44340 23548
rect 44396 23492 44406 23548
rect 58429 23492 58439 23548
rect 58495 23492 58543 23548
rect 58599 23492 58647 23548
rect 58703 23492 58713 23548
rect 1922 23436 1932 23492
rect 1988 23436 9772 23492
rect 9828 23436 9838 23492
rect 30156 23436 33292 23492
rect 33348 23436 33852 23492
rect 33908 23436 33918 23492
rect 34066 23436 34076 23492
rect 34132 23436 35868 23492
rect 35924 23436 35934 23492
rect 38546 23436 38556 23492
rect 38612 23436 43484 23492
rect 43540 23436 43820 23492
rect 43876 23436 43886 23492
rect 44706 23436 44716 23492
rect 44772 23436 44828 23492
rect 44884 23436 44894 23492
rect 45238 23436 45276 23492
rect 45332 23436 45342 23492
rect 15698 23324 15708 23380
rect 15764 23324 16604 23380
rect 16660 23324 16670 23380
rect 27010 23324 27020 23380
rect 27076 23324 28028 23380
rect 28084 23324 28924 23380
rect 28980 23324 28990 23380
rect 30156 23268 30212 23436
rect 30594 23324 30604 23380
rect 30660 23324 31724 23380
rect 31780 23324 31790 23380
rect 33506 23324 33516 23380
rect 33572 23324 34636 23380
rect 34692 23324 34702 23380
rect 38210 23324 38220 23380
rect 38276 23324 39564 23380
rect 39620 23324 39630 23380
rect 39890 23324 39900 23380
rect 39956 23324 42812 23380
rect 42868 23324 43260 23380
rect 43316 23324 49308 23380
rect 49364 23324 50204 23380
rect 50260 23324 50270 23380
rect 9174 23212 9212 23268
rect 9268 23212 9278 23268
rect 12226 23212 12236 23268
rect 12292 23212 13692 23268
rect 13748 23212 13758 23268
rect 13906 23212 13916 23268
rect 13972 23212 14028 23268
rect 14084 23212 17444 23268
rect 17388 23156 17444 23212
rect 26852 23212 30212 23268
rect 30482 23212 30492 23268
rect 30548 23212 31500 23268
rect 31556 23212 34580 23268
rect 34850 23212 34860 23268
rect 34916 23212 37884 23268
rect 37940 23212 37950 23268
rect 45266 23212 45276 23268
rect 45332 23212 45612 23268
rect 45668 23212 45678 23268
rect 46498 23212 46508 23268
rect 46564 23212 47180 23268
rect 47236 23212 48188 23268
rect 48244 23212 49084 23268
rect 49140 23212 49150 23268
rect 49634 23212 49644 23268
rect 49700 23212 50652 23268
rect 50708 23212 50718 23268
rect 26852 23156 26908 23212
rect 34524 23156 34580 23212
rect 12786 23100 12796 23156
rect 12852 23100 13356 23156
rect 13412 23100 13422 23156
rect 14130 23100 14140 23156
rect 14196 23100 15932 23156
rect 15988 23100 15998 23156
rect 17378 23100 17388 23156
rect 17444 23100 17454 23156
rect 23090 23100 23100 23156
rect 23156 23100 24332 23156
rect 24388 23100 26908 23156
rect 30146 23100 30156 23156
rect 30212 23100 30828 23156
rect 30884 23100 33180 23156
rect 33236 23100 34300 23156
rect 34356 23100 34366 23156
rect 34524 23100 38556 23156
rect 38612 23100 38622 23156
rect 39554 23100 39564 23156
rect 39620 23100 42924 23156
rect 42980 23100 42990 23156
rect 45266 23100 45276 23156
rect 45332 23100 45388 23156
rect 45444 23100 45454 23156
rect 48066 23100 48076 23156
rect 48132 23100 54348 23156
rect 54404 23100 54414 23156
rect 56018 23100 56028 23156
rect 56084 23100 56924 23156
rect 56980 23100 56990 23156
rect 2482 22988 2492 23044
rect 2548 22988 3052 23044
rect 3108 22988 3118 23044
rect 3378 22988 3388 23044
rect 3444 22988 3724 23044
rect 3780 22988 3790 23044
rect 3938 22988 3948 23044
rect 4004 22988 4620 23044
rect 4676 22988 4686 23044
rect 12674 22988 12684 23044
rect 12740 22988 15036 23044
rect 15092 22988 15102 23044
rect 25330 22988 25340 23044
rect 25396 22988 27804 23044
rect 27860 22988 27870 23044
rect 28028 22988 30268 23044
rect 30324 22988 31836 23044
rect 31892 22988 31902 23044
rect 36418 22988 36428 23044
rect 36484 22988 38332 23044
rect 38388 22988 46956 23044
rect 47012 22988 47404 23044
rect 47460 22988 47470 23044
rect 48178 22988 48188 23044
rect 48244 22988 48524 23044
rect 48580 22988 48860 23044
rect 48916 22988 48926 23044
rect 49746 22988 49756 23044
rect 49812 22988 54460 23044
rect 54516 22988 54908 23044
rect 54964 22988 54974 23044
rect 28028 22932 28084 22988
rect 6738 22876 6748 22932
rect 6804 22876 9212 22932
rect 9268 22876 9278 22932
rect 13766 22876 13804 22932
rect 13860 22876 13870 22932
rect 27346 22876 27356 22932
rect 27412 22876 28084 22932
rect 29250 22876 29260 22932
rect 29316 22876 31164 22932
rect 31220 22876 31612 22932
rect 31668 22876 31678 22932
rect 32022 22876 32060 22932
rect 32116 22876 32126 22932
rect 35298 22876 35308 22932
rect 35364 22876 37212 22932
rect 37268 22876 37278 22932
rect 37436 22876 38220 22932
rect 38276 22876 38286 22932
rect 40450 22876 40460 22932
rect 40516 22876 41692 22932
rect 41748 22876 42588 22932
rect 42644 22876 42654 22932
rect 44370 22876 44380 22932
rect 44436 22876 54236 22932
rect 54292 22876 55020 22932
rect 55076 22876 55086 22932
rect 37436 22820 37492 22876
rect 7298 22764 7308 22820
rect 7364 22764 7532 22820
rect 7588 22764 8092 22820
rect 8148 22764 8158 22820
rect 9324 22764 14252 22820
rect 14308 22764 14700 22820
rect 14756 22764 15148 22820
rect 25228 22764 35196 22820
rect 0 22624 800 22736
rect 8355 22708 8365 22764
rect 8421 22708 8469 22764
rect 8525 22708 8573 22764
rect 8629 22708 8639 22764
rect 9324 22708 9380 22764
rect 15092 22708 15148 22764
rect 22662 22708 22672 22764
rect 22728 22708 22776 22764
rect 22832 22708 22880 22764
rect 22936 22708 22946 22764
rect 25228 22708 25284 22764
rect 9314 22652 9324 22708
rect 9380 22652 9390 22708
rect 10882 22652 10892 22708
rect 10948 22652 14924 22708
rect 14980 22652 14990 22708
rect 15092 22652 15260 22708
rect 15316 22652 15326 22708
rect 25218 22652 25228 22708
rect 25284 22652 25294 22708
rect 27234 22652 27244 22708
rect 27300 22652 30604 22708
rect 30660 22652 30670 22708
rect 31266 22652 31276 22708
rect 31332 22652 33292 22708
rect 33348 22652 33358 22708
rect 35252 22596 35308 22820
rect 37314 22764 37324 22820
rect 37380 22764 37492 22820
rect 37762 22764 37772 22820
rect 37828 22764 38780 22820
rect 38836 22764 38846 22820
rect 46722 22764 46732 22820
rect 46788 22764 48972 22820
rect 49028 22764 49038 22820
rect 36969 22708 36979 22764
rect 37035 22708 37083 22764
rect 37139 22708 37187 22764
rect 37243 22708 37253 22764
rect 51276 22708 51286 22764
rect 51342 22708 51390 22764
rect 51446 22708 51494 22764
rect 51550 22708 51560 22764
rect 37958 22652 37996 22708
rect 38052 22652 38062 22708
rect 40226 22652 40236 22708
rect 40292 22652 48076 22708
rect 48132 22652 50428 22708
rect 50484 22652 50494 22708
rect 55458 22652 55468 22708
rect 55524 22652 55534 22708
rect 55468 22596 55524 22652
rect 4610 22540 4620 22596
rect 4676 22540 7756 22596
rect 7812 22540 7822 22596
rect 13906 22540 13916 22596
rect 13972 22540 15932 22596
rect 15988 22540 15998 22596
rect 21186 22540 21196 22596
rect 21252 22540 23100 22596
rect 23156 22540 23166 22596
rect 24210 22540 24220 22596
rect 24276 22540 27356 22596
rect 27412 22540 27422 22596
rect 30930 22540 30940 22596
rect 30996 22540 34748 22596
rect 34804 22540 34814 22596
rect 35252 22540 36988 22596
rect 37044 22540 37054 22596
rect 37762 22540 37772 22596
rect 37828 22540 39228 22596
rect 39284 22540 39294 22596
rect 55010 22540 55020 22596
rect 55076 22540 56700 22596
rect 56756 22540 56766 22596
rect 34748 22484 34804 22540
rect 7158 22428 7196 22484
rect 7252 22428 7262 22484
rect 15092 22428 16268 22484
rect 16324 22428 16334 22484
rect 26786 22428 26796 22484
rect 26852 22428 30828 22484
rect 30884 22428 30894 22484
rect 31938 22428 31948 22484
rect 32004 22428 32508 22484
rect 32564 22428 32574 22484
rect 34748 22428 35308 22484
rect 35364 22428 35644 22484
rect 35700 22428 35710 22484
rect 36194 22428 36204 22484
rect 36260 22428 36764 22484
rect 36820 22428 39676 22484
rect 39732 22428 39742 22484
rect 44034 22428 44044 22484
rect 44100 22428 44492 22484
rect 44548 22428 46396 22484
rect 46452 22428 46462 22484
rect 47394 22428 47404 22484
rect 47460 22428 48412 22484
rect 48468 22428 48478 22484
rect 15092 22372 15148 22428
rect 4498 22316 4508 22372
rect 4564 22316 8764 22372
rect 8820 22316 8830 22372
rect 13010 22316 13020 22372
rect 13076 22316 15148 22372
rect 20402 22316 20412 22372
rect 20468 22316 21532 22372
rect 21588 22316 22092 22372
rect 22148 22316 22158 22372
rect 22418 22316 22428 22372
rect 22484 22316 22876 22372
rect 22932 22316 25228 22372
rect 25284 22316 25294 22372
rect 28578 22316 28588 22372
rect 28644 22316 29260 22372
rect 29316 22316 29326 22372
rect 32386 22316 32396 22372
rect 32452 22316 33404 22372
rect 33460 22316 33470 22372
rect 34514 22316 34524 22372
rect 34580 22316 38444 22372
rect 38500 22316 39900 22372
rect 39956 22316 39966 22372
rect 44370 22316 44380 22372
rect 44436 22316 45500 22372
rect 45556 22316 45724 22372
rect 45780 22316 45790 22372
rect 48962 22316 48972 22372
rect 49028 22316 52892 22372
rect 52948 22316 52958 22372
rect 57250 22316 57260 22372
rect 57316 22316 57596 22372
rect 57652 22316 57662 22372
rect 2594 22204 2604 22260
rect 2660 22204 3724 22260
rect 3780 22204 3790 22260
rect 4722 22204 4732 22260
rect 4788 22204 5964 22260
rect 6020 22204 6030 22260
rect 10098 22204 10108 22260
rect 10164 22204 11340 22260
rect 11396 22204 12684 22260
rect 12740 22204 13692 22260
rect 13748 22204 13758 22260
rect 14578 22204 14588 22260
rect 14644 22204 15932 22260
rect 15988 22204 15998 22260
rect 18946 22204 18956 22260
rect 19012 22204 19404 22260
rect 19460 22204 21084 22260
rect 21140 22204 21150 22260
rect 23986 22204 23996 22260
rect 24052 22204 24892 22260
rect 24948 22204 26012 22260
rect 26068 22204 27580 22260
rect 27636 22204 30604 22260
rect 30660 22204 30670 22260
rect 31378 22204 31388 22260
rect 31444 22204 33964 22260
rect 34020 22204 36316 22260
rect 36372 22204 37660 22260
rect 37716 22204 37726 22260
rect 37874 22204 37884 22260
rect 37940 22204 38108 22260
rect 38164 22204 38174 22260
rect 39218 22204 39228 22260
rect 39284 22204 41356 22260
rect 41412 22204 41422 22260
rect 45154 22204 45164 22260
rect 45220 22204 45836 22260
rect 45892 22204 45902 22260
rect 46050 22204 46060 22260
rect 46116 22204 46620 22260
rect 46676 22204 46686 22260
rect 47394 22204 47404 22260
rect 47460 22204 47964 22260
rect 48020 22204 49308 22260
rect 49364 22204 49374 22260
rect 50418 22204 50428 22260
rect 50484 22204 51996 22260
rect 52052 22204 52444 22260
rect 52500 22204 52510 22260
rect 13346 22092 13356 22148
rect 13412 22092 13804 22148
rect 13860 22092 14140 22148
rect 14196 22092 14206 22148
rect 14354 22092 14364 22148
rect 14420 22092 14430 22148
rect 15026 22092 15036 22148
rect 15092 22092 18172 22148
rect 18228 22092 18238 22148
rect 20066 22092 20076 22148
rect 20132 22092 24220 22148
rect 24276 22092 24286 22148
rect 24434 22092 24444 22148
rect 24500 22092 25340 22148
rect 25396 22092 28588 22148
rect 28644 22092 29036 22148
rect 29092 22092 29102 22148
rect 29596 22092 31668 22148
rect 31910 22092 31948 22148
rect 32004 22092 32014 22148
rect 32610 22092 32620 22148
rect 32676 22092 35308 22148
rect 35364 22092 35756 22148
rect 35812 22092 35822 22148
rect 38108 22092 39004 22148
rect 39060 22092 40236 22148
rect 40292 22092 40302 22148
rect 40674 22092 40684 22148
rect 40740 22092 41468 22148
rect 41524 22092 41692 22148
rect 41748 22092 41758 22148
rect 43932 22092 47068 22148
rect 47170 22092 47180 22148
rect 47236 22092 47852 22148
rect 47908 22092 47918 22148
rect 50194 22092 50204 22148
rect 50260 22092 51324 22148
rect 51380 22092 53116 22148
rect 53172 22092 53182 22148
rect 14364 22036 14420 22092
rect 29596 22036 29652 22092
rect 31612 22036 31668 22092
rect 38108 22036 38164 22092
rect 43932 22036 43988 22092
rect 2790 21980 2828 22036
rect 2884 21980 2894 22036
rect 3332 21980 9772 22036
rect 9828 21980 9838 22036
rect 13990 21980 14028 22036
rect 14084 21980 14094 22036
rect 14364 21980 15428 22036
rect 15932 21980 16716 22036
rect 16772 21980 16782 22036
rect 21634 21980 21644 22036
rect 21700 21980 22092 22036
rect 22148 21980 22158 22036
rect 25778 21980 25788 22036
rect 25844 21980 26124 22036
rect 26180 21980 29652 22036
rect 31602 21980 31612 22036
rect 31668 21980 31678 22036
rect 31836 21980 36428 22036
rect 36484 21980 36494 22036
rect 38098 21980 38108 22036
rect 38164 21980 38174 22036
rect 38612 21980 43988 22036
rect 3332 21924 3388 21980
rect 4284 21924 4340 21980
rect 1586 21868 1596 21924
rect 1652 21868 3388 21924
rect 4274 21868 4284 21924
rect 4340 21868 4350 21924
rect 8978 21868 8988 21924
rect 9044 21868 9324 21924
rect 9380 21868 9390 21924
rect 15372 21812 15428 21980
rect 15508 21924 15518 21980
rect 15574 21924 15622 21980
rect 15678 21924 15726 21980
rect 15782 21924 15792 21980
rect 15932 21812 15988 21980
rect 29815 21924 29825 21980
rect 29881 21924 29929 21980
rect 29985 21924 30033 21980
rect 30089 21924 30099 21980
rect 20178 21868 20188 21924
rect 20244 21868 23604 21924
rect 25106 21868 25116 21924
rect 25172 21868 25900 21924
rect 25956 21868 26684 21924
rect 26740 21868 26750 21924
rect 23548 21812 23604 21868
rect 31836 21812 31892 21980
rect 38612 21924 38668 21980
rect 44122 21924 44132 21980
rect 44188 21924 44236 21980
rect 44292 21924 44340 21980
rect 44396 21924 44406 21980
rect 33730 21868 33740 21924
rect 33796 21868 34412 21924
rect 34468 21868 38668 21924
rect 1810 21756 1820 21812
rect 1876 21756 4844 21812
rect 4900 21756 5628 21812
rect 5684 21756 5694 21812
rect 9090 21756 9100 21812
rect 9156 21756 10668 21812
rect 10724 21756 10734 21812
rect 13458 21756 13468 21812
rect 13524 21756 13916 21812
rect 13972 21756 14420 21812
rect 14690 21756 14700 21812
rect 14756 21756 15148 21812
rect 15372 21756 15988 21812
rect 17826 21756 17836 21812
rect 17892 21756 21644 21812
rect 21700 21756 22764 21812
rect 22820 21756 22830 21812
rect 23548 21756 31892 21812
rect 32498 21756 32508 21812
rect 32564 21756 32844 21812
rect 32900 21756 32910 21812
rect 33478 21756 33516 21812
rect 33572 21756 33582 21812
rect 33842 21756 33852 21812
rect 33908 21756 38444 21812
rect 38500 21756 38668 21812
rect 39666 21756 39676 21812
rect 39732 21756 46172 21812
rect 46228 21756 46452 21812
rect 14364 21700 14420 21756
rect 15092 21700 15148 21756
rect 2482 21644 2492 21700
rect 2548 21644 14140 21700
rect 14196 21644 14206 21700
rect 14354 21644 14364 21700
rect 14420 21644 14430 21700
rect 15092 21644 15372 21700
rect 15428 21644 15596 21700
rect 15652 21644 15662 21700
rect 16034 21644 16044 21700
rect 16100 21644 16492 21700
rect 16548 21644 17500 21700
rect 17556 21644 17566 21700
rect 18498 21644 18508 21700
rect 18564 21644 19068 21700
rect 19124 21644 19134 21700
rect 22418 21644 22428 21700
rect 22484 21644 34524 21700
rect 34580 21644 34590 21700
rect 35410 21644 35420 21700
rect 35476 21644 35486 21700
rect 37426 21644 37436 21700
rect 37492 21644 37996 21700
rect 38052 21644 38062 21700
rect 38612 21644 38668 21756
rect 46396 21700 46452 21756
rect 47012 21700 47068 22092
rect 50306 21980 50316 22036
rect 50372 21980 50708 22036
rect 50652 21812 50708 21980
rect 58429 21924 58439 21980
rect 58495 21924 58543 21980
rect 58599 21924 58647 21980
rect 58703 21924 58713 21980
rect 50866 21868 50876 21924
rect 50932 21868 51324 21924
rect 51380 21868 52220 21924
rect 52276 21868 52286 21924
rect 50652 21756 50988 21812
rect 51044 21756 51054 21812
rect 54338 21756 54348 21812
rect 54404 21756 55692 21812
rect 55748 21756 55758 21812
rect 38724 21644 38734 21700
rect 40338 21644 40348 21700
rect 40404 21644 46060 21700
rect 46116 21644 46126 21700
rect 46386 21644 46396 21700
rect 46452 21644 46462 21700
rect 47012 21644 47516 21700
rect 47572 21644 47582 21700
rect 48066 21644 48076 21700
rect 48132 21644 49756 21700
rect 49812 21644 50652 21700
rect 50708 21644 50718 21700
rect 53666 21644 53676 21700
rect 53732 21644 55916 21700
rect 55972 21644 55982 21700
rect 0 21504 800 21616
rect 35420 21588 35476 21644
rect 2492 21532 3388 21588
rect 3444 21532 4620 21588
rect 4676 21532 10444 21588
rect 10500 21532 10510 21588
rect 15474 21532 15484 21588
rect 15540 21532 16604 21588
rect 16660 21532 29372 21588
rect 29428 21532 30268 21588
rect 30324 21532 30940 21588
rect 30996 21532 31006 21588
rect 31490 21532 31500 21588
rect 31556 21532 31948 21588
rect 32004 21532 32620 21588
rect 32676 21532 32686 21588
rect 32834 21532 32844 21588
rect 32900 21532 33628 21588
rect 33684 21532 33694 21588
rect 35420 21532 39228 21588
rect 39284 21532 39294 21588
rect 39442 21532 39452 21588
rect 39508 21532 40124 21588
rect 40180 21532 40908 21588
rect 40964 21532 40974 21588
rect 42914 21532 42924 21588
rect 42980 21532 44492 21588
rect 44548 21532 44558 21588
rect 2492 21364 2548 21532
rect 46060 21476 46116 21644
rect 47516 21588 47572 21644
rect 47058 21532 47068 21588
rect 47124 21532 47162 21588
rect 47516 21532 48132 21588
rect 48262 21532 48300 21588
rect 48356 21532 48366 21588
rect 50652 21532 51100 21588
rect 51156 21532 51166 21588
rect 55234 21532 55244 21588
rect 55300 21532 57372 21588
rect 57428 21532 58044 21588
rect 58100 21532 58110 21588
rect 48076 21476 48132 21532
rect 3154 21420 3164 21476
rect 3220 21420 3388 21476
rect 13346 21420 13356 21476
rect 13412 21420 21028 21476
rect 25218 21420 25228 21476
rect 25284 21420 26236 21476
rect 26292 21420 26302 21476
rect 28018 21420 28028 21476
rect 28084 21420 29148 21476
rect 29204 21420 29214 21476
rect 29586 21420 29596 21476
rect 29652 21420 30492 21476
rect 30548 21420 30558 21476
rect 32022 21420 32060 21476
rect 32116 21420 32126 21476
rect 32498 21420 32508 21476
rect 32564 21420 39340 21476
rect 39396 21420 44828 21476
rect 44884 21420 44894 21476
rect 46060 21420 47852 21476
rect 47908 21420 47918 21476
rect 48066 21420 48076 21476
rect 48132 21420 48142 21476
rect 2258 21308 2268 21364
rect 2324 21308 2548 21364
rect 3332 21364 3388 21420
rect 20972 21364 21028 21420
rect 3332 21308 3836 21364
rect 3892 21308 8540 21364
rect 8596 21308 8606 21364
rect 9986 21308 9996 21364
rect 10052 21308 10892 21364
rect 10948 21308 10958 21364
rect 15026 21308 15036 21364
rect 15092 21308 18396 21364
rect 18452 21308 18462 21364
rect 20972 21308 35252 21364
rect 35410 21308 35420 21364
rect 35476 21308 37436 21364
rect 37492 21308 37502 21364
rect 43138 21308 43148 21364
rect 43204 21308 45948 21364
rect 46004 21308 46014 21364
rect 46834 21308 46844 21364
rect 46900 21308 48412 21364
rect 48468 21308 48478 21364
rect 35196 21252 35252 21308
rect 50652 21252 50708 21532
rect 1474 21196 1484 21252
rect 1540 21196 4732 21252
rect 4788 21196 4798 21252
rect 15474 21196 15484 21252
rect 15540 21196 16380 21252
rect 16436 21196 16446 21252
rect 19170 21196 19180 21252
rect 19236 21196 19964 21252
rect 20020 21196 20030 21252
rect 26338 21196 26348 21252
rect 26404 21196 31164 21252
rect 31220 21196 31230 21252
rect 33142 21196 33180 21252
rect 33236 21196 33246 21252
rect 35196 21196 35644 21252
rect 35700 21196 36092 21252
rect 36148 21196 36158 21252
rect 37762 21196 37772 21252
rect 37828 21196 46732 21252
rect 46788 21196 46798 21252
rect 47618 21196 47628 21252
rect 47684 21196 50092 21252
rect 50148 21196 50158 21252
rect 50642 21196 50652 21252
rect 50708 21196 50718 21252
rect 8355 21140 8365 21196
rect 8421 21140 8469 21196
rect 8525 21140 8573 21196
rect 8629 21140 8639 21196
rect 22662 21140 22672 21196
rect 22728 21140 22776 21196
rect 22832 21140 22880 21196
rect 22936 21140 22946 21196
rect 2818 21084 2828 21140
rect 2884 21084 3164 21140
rect 3220 21084 3230 21140
rect 16258 21084 16268 21140
rect 16324 21084 20300 21140
rect 20356 21084 20366 21140
rect 28018 21084 28028 21140
rect 28084 21084 31948 21140
rect 32004 21084 32172 21140
rect 32228 21084 33516 21140
rect 33572 21084 33852 21140
rect 33908 21084 33918 21140
rect 36092 21028 36148 21196
rect 36969 21140 36979 21196
rect 37035 21140 37083 21196
rect 37139 21140 37187 21196
rect 37243 21140 37253 21196
rect 51276 21140 51286 21196
rect 51342 21140 51390 21196
rect 51446 21140 51494 21196
rect 51550 21140 51560 21196
rect 37650 21084 37660 21140
rect 37716 21084 37996 21140
rect 38052 21084 38062 21140
rect 45938 21084 45948 21140
rect 46004 21084 47180 21140
rect 47236 21084 47246 21140
rect 11732 20972 18956 21028
rect 19012 20972 19022 21028
rect 19506 20972 19516 21028
rect 19572 20972 34636 21028
rect 34692 20972 34702 21028
rect 36092 20972 38836 21028
rect 41458 20972 41468 21028
rect 41524 20972 41916 21028
rect 41972 20972 41982 21028
rect 47842 20972 47852 21028
rect 47908 20972 51548 21028
rect 51604 20972 51614 21028
rect 4162 20860 4172 20916
rect 4228 20860 4620 20916
rect 4676 20860 5292 20916
rect 5348 20860 5358 20916
rect 10658 20860 10668 20916
rect 10724 20860 11452 20916
rect 11508 20860 11518 20916
rect 11732 20804 11788 20972
rect 16146 20860 16156 20916
rect 16212 20860 17388 20916
rect 17444 20860 17454 20916
rect 19730 20860 19740 20916
rect 19796 20860 20972 20916
rect 21028 20860 25228 20916
rect 25284 20860 25294 20916
rect 30482 20860 30492 20916
rect 30548 20860 34972 20916
rect 35028 20860 37436 20916
rect 37492 20860 37502 20916
rect 38780 20804 38836 20972
rect 41234 20860 41244 20916
rect 41300 20860 44380 20916
rect 44436 20860 44446 20916
rect 48962 20860 48972 20916
rect 49028 20860 49084 20916
rect 49140 20860 49150 20916
rect 50866 20860 50876 20916
rect 50932 20860 51212 20916
rect 51268 20860 51278 20916
rect 11330 20748 11340 20804
rect 11396 20748 11788 20804
rect 13692 20748 16268 20804
rect 16324 20748 16334 20804
rect 16594 20748 16604 20804
rect 16660 20748 16670 20804
rect 21410 20748 21420 20804
rect 21476 20748 21980 20804
rect 22036 20748 22046 20804
rect 28466 20748 28476 20804
rect 28532 20748 30156 20804
rect 30212 20748 30222 20804
rect 32722 20748 32732 20804
rect 32788 20748 33516 20804
rect 33572 20748 33582 20804
rect 36418 20748 36428 20804
rect 36484 20748 38108 20804
rect 38164 20748 38174 20804
rect 38780 20748 50428 20804
rect 50484 20748 50494 20804
rect 50642 20748 50652 20804
rect 50708 20748 54124 20804
rect 54180 20748 54190 20804
rect 2482 20636 2492 20692
rect 2548 20636 3276 20692
rect 3332 20636 3342 20692
rect 13692 20580 13748 20748
rect 14914 20636 14924 20692
rect 14980 20636 15932 20692
rect 15988 20636 15998 20692
rect 16604 20580 16660 20748
rect 21298 20636 21308 20692
rect 21364 20636 23772 20692
rect 23828 20636 29260 20692
rect 29316 20636 29326 20692
rect 30706 20636 30716 20692
rect 30772 20636 31052 20692
rect 31108 20636 31118 20692
rect 32134 20636 32172 20692
rect 32228 20636 32238 20692
rect 33842 20636 33852 20692
rect 33908 20636 35420 20692
rect 35476 20636 35486 20692
rect 37986 20636 37996 20692
rect 38052 20636 39452 20692
rect 39508 20636 42028 20692
rect 42084 20636 42094 20692
rect 46050 20636 46060 20692
rect 46116 20636 46620 20692
rect 46676 20636 47628 20692
rect 47684 20636 47694 20692
rect 52882 20636 52892 20692
rect 52948 20636 54460 20692
rect 54516 20636 54526 20692
rect 9762 20524 9772 20580
rect 9828 20524 13692 20580
rect 13748 20524 13758 20580
rect 13906 20524 13916 20580
rect 13972 20524 16660 20580
rect 32498 20524 32508 20580
rect 32564 20524 40460 20580
rect 40516 20524 40796 20580
rect 40852 20524 40862 20580
rect 41570 20524 41580 20580
rect 41636 20524 42924 20580
rect 42980 20524 42990 20580
rect 46162 20524 46172 20580
rect 46228 20524 53564 20580
rect 53620 20524 53630 20580
rect 55682 20524 55692 20580
rect 55748 20524 56812 20580
rect 56868 20524 56878 20580
rect 0 20384 800 20496
rect 1698 20412 1708 20468
rect 1764 20412 2044 20468
rect 2100 20412 2110 20468
rect 4498 20412 4508 20468
rect 4564 20412 10332 20468
rect 10388 20412 10398 20468
rect 18498 20412 18508 20468
rect 18564 20412 19740 20468
rect 19796 20412 19806 20468
rect 36194 20412 36204 20468
rect 36260 20412 36764 20468
rect 36820 20412 36830 20468
rect 49186 20412 49196 20468
rect 49252 20412 50204 20468
rect 50260 20412 50270 20468
rect 50418 20412 50428 20468
rect 50484 20412 50876 20468
rect 50932 20412 51996 20468
rect 52052 20412 52062 20468
rect 54786 20412 54796 20468
rect 54852 20412 56140 20468
rect 56196 20412 56700 20468
rect 56756 20412 56766 20468
rect 15508 20356 15518 20412
rect 15574 20356 15622 20412
rect 15678 20356 15726 20412
rect 15782 20356 15792 20412
rect 29815 20356 29825 20412
rect 29881 20356 29929 20412
rect 29985 20356 30033 20412
rect 30089 20356 30099 20412
rect 44122 20356 44132 20412
rect 44188 20356 44236 20412
rect 44292 20356 44340 20412
rect 44396 20356 44406 20412
rect 58429 20356 58439 20412
rect 58495 20356 58543 20412
rect 58599 20356 58647 20412
rect 58703 20356 58713 20412
rect 12114 20300 12124 20356
rect 12180 20300 14924 20356
rect 14980 20300 14990 20356
rect 18050 20300 18060 20356
rect 18116 20300 19516 20356
rect 19572 20300 19582 20356
rect 36082 20300 36092 20356
rect 36148 20300 36652 20356
rect 36708 20300 36718 20356
rect 48850 20300 48860 20356
rect 48916 20300 50316 20356
rect 50372 20300 50382 20356
rect 3714 20188 3724 20244
rect 3780 20188 5180 20244
rect 5236 20188 5246 20244
rect 5506 20188 5516 20244
rect 5572 20188 8988 20244
rect 9044 20188 9054 20244
rect 15922 20188 15932 20244
rect 15988 20188 17500 20244
rect 17556 20188 18172 20244
rect 18228 20188 18238 20244
rect 19282 20188 19292 20244
rect 19348 20188 26012 20244
rect 26068 20188 26078 20244
rect 29698 20188 29708 20244
rect 29764 20188 31388 20244
rect 31444 20188 34636 20244
rect 34692 20188 44940 20244
rect 44996 20188 45006 20244
rect 49410 20188 49420 20244
rect 49476 20188 53116 20244
rect 53172 20188 53182 20244
rect 3378 20076 3388 20132
rect 3444 20076 4396 20132
rect 4452 20076 4462 20132
rect 4946 20076 4956 20132
rect 5012 20076 7420 20132
rect 7476 20076 7486 20132
rect 11106 20076 11116 20132
rect 11172 20076 11788 20132
rect 11844 20076 12572 20132
rect 12628 20076 12638 20132
rect 16492 20076 17612 20132
rect 17668 20076 22092 20132
rect 22148 20076 23100 20132
rect 23156 20076 23166 20132
rect 24658 20076 24668 20132
rect 24724 20076 26348 20132
rect 26404 20076 26414 20132
rect 28102 20076 28140 20132
rect 28196 20076 28206 20132
rect 30706 20076 30716 20132
rect 30772 20076 32508 20132
rect 32564 20076 32574 20132
rect 35186 20076 35196 20132
rect 35252 20076 37884 20132
rect 37940 20076 37950 20132
rect 43922 20076 43932 20132
rect 43988 20076 44716 20132
rect 44772 20076 44782 20132
rect 45378 20076 45388 20132
rect 45444 20076 47852 20132
rect 47908 20076 49644 20132
rect 49700 20076 50316 20132
rect 50372 20076 50382 20132
rect 51202 20076 51212 20132
rect 51268 20076 51996 20132
rect 52052 20076 52780 20132
rect 52836 20076 52846 20132
rect 52994 20076 53004 20132
rect 53060 20076 55804 20132
rect 55860 20076 57036 20132
rect 57092 20076 57102 20132
rect 16492 20020 16548 20076
rect 700 19964 1708 20020
rect 1764 19964 5068 20020
rect 5124 19964 5134 20020
rect 9090 19964 9100 20020
rect 9156 19964 10780 20020
rect 10836 19964 11452 20020
rect 11508 19964 11518 20020
rect 15092 19964 16548 20020
rect 16706 19964 16716 20020
rect 16772 19964 28028 20020
rect 28084 19964 28094 20020
rect 28354 19964 28364 20020
rect 28420 19964 28700 20020
rect 28756 19964 30156 20020
rect 30212 19964 30222 20020
rect 31938 19964 31948 20020
rect 32004 19964 33180 20020
rect 33236 19964 35308 20020
rect 35364 19964 35374 20020
rect 36204 19964 38444 20020
rect 38500 19964 38510 20020
rect 38770 19964 38780 20020
rect 38836 19964 39676 20020
rect 39732 19964 39742 20020
rect 42354 19964 42364 20020
rect 42420 19964 43260 20020
rect 43316 19964 43326 20020
rect 44034 19964 44044 20020
rect 44100 19964 46508 20020
rect 46564 19964 46574 20020
rect 48066 19964 48076 20020
rect 48132 19964 48972 20020
rect 49028 19964 49038 20020
rect 49746 19964 49756 20020
rect 49812 19964 52556 20020
rect 52612 19964 52622 20020
rect 700 19572 756 19964
rect 15092 19908 15148 19964
rect 36204 19908 36260 19964
rect 2034 19852 2044 19908
rect 2100 19852 2604 19908
rect 2660 19852 2670 19908
rect 11106 19852 11116 19908
rect 11172 19852 11900 19908
rect 11956 19852 12460 19908
rect 12516 19852 12526 19908
rect 13682 19852 13692 19908
rect 13748 19852 14588 19908
rect 14644 19852 15148 19908
rect 18946 19852 18956 19908
rect 19012 19852 20188 19908
rect 20244 19852 20636 19908
rect 20692 19852 20702 19908
rect 24322 19852 24332 19908
rect 24388 19852 25676 19908
rect 25732 19852 25742 19908
rect 28130 19852 28140 19908
rect 28196 19852 33460 19908
rect 36194 19852 36204 19908
rect 36260 19852 36270 19908
rect 37538 19852 37548 19908
rect 37604 19852 39228 19908
rect 39284 19852 39294 19908
rect 46022 19852 46060 19908
rect 46116 19852 46126 19908
rect 47394 19852 47404 19908
rect 47460 19852 53788 19908
rect 53844 19852 53854 19908
rect 56018 19852 56028 19908
rect 56084 19852 56588 19908
rect 56644 19852 56654 19908
rect 33404 19796 33460 19852
rect 3714 19740 3724 19796
rect 3780 19740 4060 19796
rect 4116 19740 4126 19796
rect 6738 19740 6748 19796
rect 6804 19740 8652 19796
rect 8708 19740 13468 19796
rect 13524 19740 13534 19796
rect 17826 19740 17836 19796
rect 17892 19740 19180 19796
rect 19236 19740 19246 19796
rect 32274 19740 32284 19796
rect 32340 19740 33068 19796
rect 33124 19740 33134 19796
rect 33404 19740 40348 19796
rect 40404 19740 40684 19796
rect 40740 19740 40750 19796
rect 43922 19740 43932 19796
rect 43988 19740 52108 19796
rect 52164 19740 52174 19796
rect 32722 19628 32732 19684
rect 32788 19628 34636 19684
rect 34692 19628 34702 19684
rect 37650 19628 37660 19684
rect 37716 19628 38668 19684
rect 38724 19628 38734 19684
rect 39330 19628 39340 19684
rect 39396 19628 41020 19684
rect 41076 19628 48748 19684
rect 48804 19628 48814 19684
rect 50418 19628 50428 19684
rect 50484 19628 50540 19684
rect 50596 19628 50606 19684
rect 8355 19572 8365 19628
rect 8421 19572 8469 19628
rect 8525 19572 8573 19628
rect 8629 19572 8639 19628
rect 22662 19572 22672 19628
rect 22728 19572 22776 19628
rect 22832 19572 22880 19628
rect 22936 19572 22946 19628
rect 36969 19572 36979 19628
rect 37035 19572 37083 19628
rect 37139 19572 37187 19628
rect 37243 19572 37253 19628
rect 51276 19572 51286 19628
rect 51342 19572 51390 19628
rect 51446 19572 51494 19628
rect 51550 19572 51560 19628
rect 700 19516 980 19572
rect 7410 19516 7420 19572
rect 7476 19516 7756 19572
rect 7812 19516 7822 19572
rect 10322 19516 10332 19572
rect 10388 19516 10780 19572
rect 10836 19516 10846 19572
rect 19842 19516 19852 19572
rect 19908 19516 20188 19572
rect 20244 19516 21532 19572
rect 21588 19516 21598 19572
rect 31938 19516 31948 19572
rect 32004 19516 32844 19572
rect 32900 19516 32910 19572
rect 38546 19516 38556 19572
rect 38612 19516 40124 19572
rect 40180 19516 47180 19572
rect 47236 19516 47246 19572
rect 49522 19516 49532 19572
rect 49588 19516 49980 19572
rect 50036 19516 50046 19572
rect 0 19348 800 19376
rect 924 19348 980 19516
rect 10332 19460 10388 19516
rect 8082 19404 8092 19460
rect 8148 19404 10388 19460
rect 11732 19404 29764 19460
rect 29922 19404 29932 19460
rect 29988 19404 32732 19460
rect 32788 19404 32798 19460
rect 33058 19404 33068 19460
rect 33124 19404 34412 19460
rect 34468 19404 34478 19460
rect 48962 19404 48972 19460
rect 49028 19404 50204 19460
rect 50260 19404 50270 19460
rect 53890 19404 53900 19460
rect 53956 19404 55916 19460
rect 55972 19404 56812 19460
rect 56868 19404 56878 19460
rect 11732 19348 11788 19404
rect 29708 19348 29764 19404
rect 0 19292 980 19348
rect 2706 19292 2716 19348
rect 2772 19292 3612 19348
rect 3668 19292 3678 19348
rect 8194 19292 8204 19348
rect 8260 19292 9212 19348
rect 9268 19292 11788 19348
rect 12786 19292 12796 19348
rect 12852 19292 17164 19348
rect 17220 19292 17230 19348
rect 22866 19292 22876 19348
rect 22932 19292 23996 19348
rect 24052 19292 29260 19348
rect 29316 19292 29326 19348
rect 29708 19292 35308 19348
rect 35364 19292 35374 19348
rect 35970 19292 35980 19348
rect 36036 19292 37996 19348
rect 38052 19292 38062 19348
rect 40450 19292 40460 19348
rect 40516 19292 45164 19348
rect 45220 19292 47404 19348
rect 47460 19292 47470 19348
rect 50530 19292 50540 19348
rect 50596 19292 51548 19348
rect 51604 19292 52668 19348
rect 52724 19292 52734 19348
rect 0 19264 800 19292
rect 1698 19180 1708 19236
rect 1764 19180 1932 19236
rect 1988 19180 5740 19236
rect 5796 19180 5806 19236
rect 6514 19180 6524 19236
rect 6580 19180 7196 19236
rect 7252 19180 7262 19236
rect 12674 19180 12684 19236
rect 12740 19180 17276 19236
rect 17332 19180 18956 19236
rect 19012 19180 19022 19236
rect 20066 19180 20076 19236
rect 20132 19180 20972 19236
rect 21028 19180 21038 19236
rect 22754 19180 22764 19236
rect 22820 19180 23772 19236
rect 23828 19180 23838 19236
rect 28466 19180 28476 19236
rect 28532 19180 29036 19236
rect 29092 19180 29102 19236
rect 33058 19180 33068 19236
rect 33124 19180 34524 19236
rect 34580 19180 34590 19236
rect 34738 19180 34748 19236
rect 34804 19180 37660 19236
rect 37716 19180 37726 19236
rect 41794 19180 41804 19236
rect 41860 19180 43260 19236
rect 43316 19180 43326 19236
rect 46946 19180 46956 19236
rect 47012 19180 47852 19236
rect 47908 19180 47918 19236
rect 48178 19180 48188 19236
rect 48244 19180 51772 19236
rect 51828 19180 52892 19236
rect 52948 19180 52958 19236
rect 55010 19180 55020 19236
rect 55076 19180 55692 19236
rect 55748 19180 55758 19236
rect 3602 19068 3612 19124
rect 3668 19068 6300 19124
rect 6356 19068 6366 19124
rect 8306 19068 8316 19124
rect 8372 19068 8988 19124
rect 9044 19068 9054 19124
rect 10434 19068 10444 19124
rect 10500 19068 11452 19124
rect 11508 19068 11518 19124
rect 12786 19068 12796 19124
rect 12852 19068 15820 19124
rect 15876 19068 17612 19124
rect 17668 19068 17678 19124
rect 26674 19068 26684 19124
rect 26740 19068 26908 19124
rect 26964 19068 26974 19124
rect 28130 19068 28140 19124
rect 28196 19068 29484 19124
rect 29540 19068 33180 19124
rect 33236 19068 33246 19124
rect 35252 19068 35644 19124
rect 35700 19068 35756 19124
rect 35812 19068 35822 19124
rect 36082 19068 36092 19124
rect 36148 19068 36158 19124
rect 37762 19068 37772 19124
rect 37828 19068 44828 19124
rect 44884 19068 44894 19124
rect 46722 19068 46732 19124
rect 46788 19068 47292 19124
rect 47348 19068 47358 19124
rect 47628 19068 48636 19124
rect 48692 19068 49420 19124
rect 49476 19068 49486 19124
rect 49746 19068 49756 19124
rect 49812 19068 50316 19124
rect 50372 19068 50382 19124
rect 26684 19012 26740 19068
rect 6066 18956 6076 19012
rect 6132 18956 7532 19012
rect 7588 18956 7598 19012
rect 13794 18956 13804 19012
rect 13860 18956 14364 19012
rect 14420 18956 14430 19012
rect 15092 18956 15484 19012
rect 15540 18956 15932 19012
rect 15988 18956 16492 19012
rect 16548 18956 16558 19012
rect 17154 18956 17164 19012
rect 17220 18956 17724 19012
rect 17780 18956 17790 19012
rect 18722 18956 18732 19012
rect 18788 18956 19404 19012
rect 19460 18956 23772 19012
rect 23828 18956 23838 19012
rect 25442 18956 25452 19012
rect 25508 18956 26348 19012
rect 26404 18956 26740 19012
rect 26852 18956 30604 19012
rect 30660 18956 30670 19012
rect 3490 18844 3500 18900
rect 3556 18844 4284 18900
rect 4340 18844 4350 18900
rect 15092 18676 15148 18956
rect 26852 18900 26908 18956
rect 35252 18900 35308 19068
rect 36092 19012 36148 19068
rect 36092 18956 38668 19012
rect 41346 18956 41356 19012
rect 41412 18956 42028 19012
rect 42084 18956 42094 19012
rect 43932 18956 45556 19012
rect 45714 18956 45724 19012
rect 45780 18956 46060 19012
rect 46116 18956 46126 19012
rect 19506 18844 19516 18900
rect 19572 18844 26908 18900
rect 30258 18844 30268 18900
rect 30324 18844 35308 18900
rect 35522 18844 35532 18900
rect 35588 18844 36428 18900
rect 36484 18844 36494 18900
rect 15508 18788 15518 18844
rect 15574 18788 15622 18844
rect 15678 18788 15726 18844
rect 15782 18788 15792 18844
rect 29815 18788 29825 18844
rect 29881 18788 29929 18844
rect 29985 18788 30033 18844
rect 30089 18788 30099 18844
rect 38612 18788 38668 18956
rect 43932 18788 43988 18956
rect 45500 18900 45556 18956
rect 47628 18900 47684 19068
rect 47852 18956 48860 19012
rect 48916 18956 49532 19012
rect 49588 18956 49598 19012
rect 47852 18900 47908 18956
rect 45500 18844 47684 18900
rect 47842 18844 47852 18900
rect 47908 18844 47918 18900
rect 49046 18844 49084 18900
rect 49140 18844 49150 18900
rect 44122 18788 44132 18844
rect 44188 18788 44236 18844
rect 44292 18788 44340 18844
rect 44396 18788 44406 18844
rect 58429 18788 58439 18844
rect 58495 18788 58543 18844
rect 58599 18788 58647 18844
rect 58703 18788 58713 18844
rect 16818 18732 16828 18788
rect 16884 18732 17500 18788
rect 17556 18732 19068 18788
rect 19124 18732 26908 18788
rect 34178 18732 34188 18788
rect 34244 18732 37548 18788
rect 37604 18732 37614 18788
rect 38612 18732 43988 18788
rect 47954 18732 47964 18788
rect 48020 18732 48188 18788
rect 48244 18732 48254 18788
rect 2482 18620 2492 18676
rect 2548 18620 3500 18676
rect 3556 18620 3566 18676
rect 7522 18620 7532 18676
rect 7588 18620 8652 18676
rect 8708 18620 8718 18676
rect 13570 18620 13580 18676
rect 13636 18620 15148 18676
rect 24658 18620 24668 18676
rect 24724 18620 25788 18676
rect 25844 18620 25854 18676
rect 26852 18564 26908 18732
rect 32274 18620 32284 18676
rect 32340 18620 33292 18676
rect 33348 18620 33358 18676
rect 35298 18620 35308 18676
rect 35364 18620 36316 18676
rect 36372 18620 36382 18676
rect 36726 18620 36764 18676
rect 36820 18620 36830 18676
rect 37874 18620 37884 18676
rect 37940 18620 38780 18676
rect 38836 18620 38846 18676
rect 42690 18620 42700 18676
rect 42756 18620 44492 18676
rect 44548 18620 44558 18676
rect 12898 18508 12908 18564
rect 12964 18508 23212 18564
rect 23268 18508 23278 18564
rect 24770 18508 24780 18564
rect 24836 18508 26684 18564
rect 26740 18508 26750 18564
rect 26852 18508 48188 18564
rect 48244 18508 48254 18564
rect 49522 18508 49532 18564
rect 49588 18508 50428 18564
rect 50484 18508 50494 18564
rect 4834 18396 4844 18452
rect 4900 18396 5516 18452
rect 5572 18396 6524 18452
rect 6580 18396 6590 18452
rect 9202 18396 9212 18452
rect 9268 18396 9436 18452
rect 9492 18396 10332 18452
rect 10388 18396 10398 18452
rect 10546 18396 10556 18452
rect 10612 18396 11452 18452
rect 11508 18396 11518 18452
rect 13234 18396 13244 18452
rect 13300 18396 17948 18452
rect 18004 18396 18014 18452
rect 20626 18396 20636 18452
rect 20692 18396 22204 18452
rect 22260 18396 29260 18452
rect 29316 18396 29326 18452
rect 29810 18396 29820 18452
rect 29876 18396 30716 18452
rect 30772 18396 30782 18452
rect 32386 18396 32396 18452
rect 32452 18396 33068 18452
rect 33124 18396 34636 18452
rect 34692 18396 34702 18452
rect 36866 18396 36876 18452
rect 36932 18396 36942 18452
rect 37314 18396 37324 18452
rect 37380 18396 38332 18452
rect 38388 18396 38398 18452
rect 42018 18396 42028 18452
rect 42084 18396 44380 18452
rect 44436 18396 44446 18452
rect 47170 18396 47180 18452
rect 47236 18396 47964 18452
rect 48020 18396 48030 18452
rect 50194 18396 50204 18452
rect 50260 18396 50428 18452
rect 50754 18396 50764 18452
rect 50820 18396 55132 18452
rect 55188 18396 55198 18452
rect 36876 18340 36932 18396
rect 50372 18340 50428 18396
rect 6402 18284 6412 18340
rect 6468 18284 7308 18340
rect 7364 18284 12348 18340
rect 12404 18284 16940 18340
rect 16996 18284 17006 18340
rect 18050 18284 18060 18340
rect 18116 18284 18126 18340
rect 21298 18284 21308 18340
rect 21364 18284 21980 18340
rect 22036 18284 22046 18340
rect 28018 18284 28028 18340
rect 28084 18284 28476 18340
rect 28532 18284 30380 18340
rect 30436 18284 30446 18340
rect 35858 18284 35868 18340
rect 35924 18284 38668 18340
rect 42886 18284 42924 18340
rect 42980 18284 42990 18340
rect 43250 18284 43260 18340
rect 43316 18284 44156 18340
rect 44212 18284 45164 18340
rect 45220 18284 45230 18340
rect 50372 18284 54796 18340
rect 54852 18284 55580 18340
rect 55636 18284 55646 18340
rect 56018 18284 56028 18340
rect 56084 18284 56812 18340
rect 56868 18284 56878 18340
rect 0 18228 800 18256
rect 18060 18228 18116 18284
rect 0 18172 1708 18228
rect 1764 18172 1774 18228
rect 6178 18172 6188 18228
rect 6244 18172 7644 18228
rect 7700 18172 7710 18228
rect 7868 18172 12684 18228
rect 12740 18172 12750 18228
rect 18060 18172 26908 18228
rect 27906 18172 27916 18228
rect 27972 18172 30604 18228
rect 30660 18172 31276 18228
rect 31332 18172 31342 18228
rect 36978 18172 36988 18228
rect 37044 18172 37604 18228
rect 0 18144 800 18172
rect 7868 18116 7924 18172
rect 26852 18116 26908 18172
rect 5170 18060 5180 18116
rect 5236 18060 7924 18116
rect 10434 18060 10444 18116
rect 10500 18060 10892 18116
rect 10948 18060 12908 18116
rect 12964 18060 13468 18116
rect 13524 18060 13534 18116
rect 26852 18060 30156 18116
rect 30212 18060 30222 18116
rect 33730 18060 33740 18116
rect 33796 18060 34860 18116
rect 34916 18060 34926 18116
rect 8355 18004 8365 18060
rect 8421 18004 8469 18060
rect 8525 18004 8573 18060
rect 8629 18004 8639 18060
rect 22662 18004 22672 18060
rect 22728 18004 22776 18060
rect 22832 18004 22880 18060
rect 22936 18004 22946 18060
rect 36969 18004 36979 18060
rect 37035 18004 37083 18060
rect 37139 18004 37187 18060
rect 37243 18004 37253 18060
rect 37548 18004 37604 18172
rect 38612 18116 38668 18284
rect 40114 18172 40124 18228
rect 40180 18172 46844 18228
rect 46900 18172 49308 18228
rect 49364 18172 50092 18228
rect 50148 18172 50158 18228
rect 38612 18060 45724 18116
rect 45780 18060 45790 18116
rect 51276 18004 51286 18060
rect 51342 18004 51390 18060
rect 51446 18004 51494 18060
rect 51550 18004 51560 18060
rect 2818 17948 2828 18004
rect 2884 17948 3500 18004
rect 3556 17948 3566 18004
rect 14802 17948 14812 18004
rect 14868 17948 15260 18004
rect 15316 17948 15326 18004
rect 33842 17948 33852 18004
rect 33908 17948 35868 18004
rect 35924 17948 35934 18004
rect 37538 17948 37548 18004
rect 37604 17948 37614 18004
rect 45154 17948 45164 18004
rect 45220 17948 47068 18004
rect 47124 17948 47134 18004
rect 47478 17948 47516 18004
rect 47572 17948 47582 18004
rect 15026 17836 15036 17892
rect 15092 17836 16604 17892
rect 16660 17836 16670 17892
rect 22306 17836 22316 17892
rect 22372 17836 23548 17892
rect 23604 17836 23614 17892
rect 29138 17836 29148 17892
rect 29204 17836 30044 17892
rect 30100 17836 30110 17892
rect 34290 17836 34300 17892
rect 34356 17836 38668 17892
rect 41122 17836 41132 17892
rect 41188 17836 41468 17892
rect 41524 17836 41534 17892
rect 42914 17836 42924 17892
rect 42980 17836 44716 17892
rect 44772 17836 44782 17892
rect 47404 17836 55692 17892
rect 55748 17836 55758 17892
rect 38612 17780 38668 17836
rect 47404 17780 47460 17836
rect 7158 17724 7196 17780
rect 7252 17724 7980 17780
rect 8036 17724 8046 17780
rect 9538 17724 9548 17780
rect 9604 17724 10220 17780
rect 10276 17724 11788 17780
rect 11844 17724 11854 17780
rect 12562 17724 12572 17780
rect 12628 17724 13356 17780
rect 13412 17724 13422 17780
rect 16706 17724 16716 17780
rect 16772 17724 19292 17780
rect 19348 17724 19628 17780
rect 19684 17724 20188 17780
rect 20244 17724 20254 17780
rect 23650 17724 23660 17780
rect 23716 17724 24220 17780
rect 24276 17724 33740 17780
rect 33796 17724 33806 17780
rect 35074 17724 35084 17780
rect 35140 17724 37100 17780
rect 37156 17724 37166 17780
rect 37314 17724 37324 17780
rect 37380 17724 38108 17780
rect 38164 17724 38174 17780
rect 38612 17724 39340 17780
rect 39396 17724 39406 17780
rect 40338 17724 40348 17780
rect 40404 17724 43148 17780
rect 43204 17724 43214 17780
rect 43820 17724 47460 17780
rect 54450 17724 54460 17780
rect 54516 17724 55244 17780
rect 55300 17724 55310 17780
rect 43820 17668 43876 17724
rect 1698 17612 1708 17668
rect 1764 17612 6412 17668
rect 6468 17612 6478 17668
rect 8530 17612 8540 17668
rect 8596 17612 10668 17668
rect 10724 17612 10734 17668
rect 11442 17612 11452 17668
rect 11508 17612 12124 17668
rect 12180 17612 12190 17668
rect 13010 17612 13020 17668
rect 13076 17612 14028 17668
rect 14084 17612 14094 17668
rect 20514 17612 20524 17668
rect 20580 17612 21308 17668
rect 21364 17612 21374 17668
rect 27906 17612 27916 17668
rect 27972 17612 29148 17668
rect 29204 17612 29214 17668
rect 32722 17612 32732 17668
rect 32788 17612 34412 17668
rect 34468 17612 34478 17668
rect 34738 17612 34748 17668
rect 34804 17612 35532 17668
rect 35588 17612 35598 17668
rect 43810 17612 43820 17668
rect 43876 17612 43886 17668
rect 45938 17612 45948 17668
rect 46004 17612 53116 17668
rect 53172 17612 53182 17668
rect 55570 17612 55580 17668
rect 55636 17612 57148 17668
rect 57204 17612 57214 17668
rect 3490 17500 3500 17556
rect 3556 17500 3948 17556
rect 4004 17500 9772 17556
rect 9828 17500 9838 17556
rect 13542 17500 13580 17556
rect 13636 17500 13646 17556
rect 14242 17500 14252 17556
rect 14308 17500 15260 17556
rect 15316 17500 16492 17556
rect 16548 17500 16558 17556
rect 20402 17500 20412 17556
rect 20468 17500 21532 17556
rect 21588 17500 21598 17556
rect 24546 17500 24556 17556
rect 24612 17500 26796 17556
rect 26852 17500 26862 17556
rect 35606 17500 35644 17556
rect 35700 17500 35710 17556
rect 47842 17500 47852 17556
rect 47908 17500 48748 17556
rect 48804 17500 48814 17556
rect 49074 17500 49084 17556
rect 49140 17500 54684 17556
rect 54740 17500 54750 17556
rect 57026 17500 57036 17556
rect 57092 17500 57708 17556
rect 57764 17500 57774 17556
rect 3714 17388 3724 17444
rect 3780 17388 4172 17444
rect 4228 17388 5628 17444
rect 5684 17388 5694 17444
rect 10994 17388 11004 17444
rect 11060 17388 14028 17444
rect 14084 17388 14094 17444
rect 15092 17388 16268 17444
rect 16324 17388 16334 17444
rect 18050 17388 18060 17444
rect 18116 17388 18126 17444
rect 25890 17388 25900 17444
rect 25956 17388 31052 17444
rect 31108 17388 33068 17444
rect 33124 17388 33134 17444
rect 34402 17388 34412 17444
rect 34468 17388 34972 17444
rect 35028 17388 48972 17444
rect 49028 17388 49532 17444
rect 49588 17388 50092 17444
rect 50148 17388 50158 17444
rect 50978 17388 50988 17444
rect 51044 17388 55580 17444
rect 55636 17388 55646 17444
rect 56018 17388 56028 17444
rect 56084 17388 57932 17444
rect 57988 17388 57998 17444
rect 5628 17332 5684 17388
rect 15092 17332 15148 17388
rect 2034 17276 2044 17332
rect 2100 17276 2828 17332
rect 2884 17276 2894 17332
rect 5628 17276 15148 17332
rect 16006 17276 16044 17332
rect 16100 17276 16110 17332
rect 15508 17220 15518 17276
rect 15574 17220 15622 17276
rect 15678 17220 15726 17276
rect 15782 17220 15792 17276
rect 18060 17220 18116 17388
rect 30818 17276 30828 17332
rect 30884 17276 31388 17332
rect 31444 17276 31454 17332
rect 31714 17276 31724 17332
rect 31780 17276 35084 17332
rect 35140 17276 35150 17332
rect 47954 17276 47964 17332
rect 48020 17276 50764 17332
rect 50820 17276 50830 17332
rect 29815 17220 29825 17276
rect 29881 17220 29929 17276
rect 29985 17220 30033 17276
rect 30089 17220 30099 17276
rect 44122 17220 44132 17276
rect 44188 17220 44236 17276
rect 44292 17220 44340 17276
rect 44396 17220 44406 17276
rect 58429 17220 58439 17276
rect 58495 17220 58543 17276
rect 58599 17220 58647 17276
rect 58703 17220 58713 17276
rect 7746 17164 7756 17220
rect 7812 17164 8988 17220
rect 9044 17164 9436 17220
rect 9492 17164 9502 17220
rect 18060 17164 26908 17220
rect 26964 17164 26974 17220
rect 30594 17164 30604 17220
rect 30660 17164 32172 17220
rect 32228 17164 43036 17220
rect 43092 17164 43102 17220
rect 45266 17164 45276 17220
rect 45332 17164 45948 17220
rect 46004 17164 47740 17220
rect 47796 17164 47806 17220
rect 50418 17164 50428 17220
rect 50484 17164 50876 17220
rect 50932 17164 50942 17220
rect 0 17108 800 17136
rect 43036 17108 43092 17164
rect 0 17052 2604 17108
rect 2660 17052 2670 17108
rect 9090 17052 9100 17108
rect 9156 17052 10108 17108
rect 10164 17052 13356 17108
rect 13412 17052 13422 17108
rect 14466 17052 14476 17108
rect 14532 17052 18172 17108
rect 18228 17052 18238 17108
rect 20850 17052 20860 17108
rect 20916 17052 23100 17108
rect 23156 17052 23166 17108
rect 23314 17052 23324 17108
rect 23380 17052 33180 17108
rect 33236 17052 33246 17108
rect 33730 17052 33740 17108
rect 33796 17052 34748 17108
rect 34804 17052 35868 17108
rect 35924 17052 35934 17108
rect 43036 17052 46508 17108
rect 46564 17052 46956 17108
rect 47012 17052 47022 17108
rect 49858 17052 49868 17108
rect 49924 17052 51212 17108
rect 51268 17052 51278 17108
rect 55906 17052 55916 17108
rect 55972 17052 57148 17108
rect 57204 17052 57214 17108
rect 0 17024 800 17052
rect 2706 16940 2716 16996
rect 2772 16940 6972 16996
rect 7028 16940 7038 16996
rect 8866 16940 8876 16996
rect 8932 16940 9548 16996
rect 9604 16940 10892 16996
rect 10948 16940 13244 16996
rect 13300 16940 13310 16996
rect 13794 16940 13804 16996
rect 13860 16940 15260 16996
rect 15316 16940 15326 16996
rect 15698 16940 15708 16996
rect 15764 16940 17836 16996
rect 17892 16940 17902 16996
rect 20962 16940 20972 16996
rect 21028 16940 23436 16996
rect 23492 16940 25340 16996
rect 25396 16940 25406 16996
rect 26852 16940 30492 16996
rect 30548 16940 31724 16996
rect 31780 16940 31790 16996
rect 33394 16940 33404 16996
rect 33460 16940 33852 16996
rect 33908 16940 34636 16996
rect 34692 16940 38668 16996
rect 38724 16940 38734 16996
rect 40226 16940 40236 16996
rect 40292 16940 41244 16996
rect 41300 16940 45724 16996
rect 45780 16940 46172 16996
rect 46228 16940 46732 16996
rect 46788 16940 46798 16996
rect 47282 16940 47292 16996
rect 47348 16940 47852 16996
rect 47908 16940 49980 16996
rect 50036 16940 50046 16996
rect 1810 16828 1820 16884
rect 1876 16828 3052 16884
rect 3108 16828 6300 16884
rect 6356 16828 6366 16884
rect 13122 16828 13132 16884
rect 13188 16828 14700 16884
rect 14756 16828 14766 16884
rect 14924 16828 15372 16884
rect 15428 16828 15438 16884
rect 15922 16828 15932 16884
rect 15988 16828 16268 16884
rect 16324 16828 16334 16884
rect 16594 16828 16604 16884
rect 16660 16828 17052 16884
rect 17108 16828 18060 16884
rect 18116 16828 18126 16884
rect 21186 16828 21196 16884
rect 21252 16828 21868 16884
rect 21924 16828 21934 16884
rect 24770 16828 24780 16884
rect 24836 16828 25676 16884
rect 25732 16828 25742 16884
rect 14924 16772 14980 16828
rect 26852 16772 26908 16940
rect 29474 16828 29484 16884
rect 29540 16828 30716 16884
rect 30772 16828 30782 16884
rect 32386 16828 32396 16884
rect 32452 16828 33964 16884
rect 34020 16828 34412 16884
rect 34468 16828 34478 16884
rect 36194 16828 36204 16884
rect 36260 16828 36652 16884
rect 36708 16828 36718 16884
rect 36866 16828 36876 16884
rect 36932 16828 38108 16884
rect 38164 16828 38174 16884
rect 39554 16828 39564 16884
rect 39620 16828 40908 16884
rect 40964 16828 41132 16884
rect 41188 16828 41198 16884
rect 42018 16828 42028 16884
rect 42084 16828 42700 16884
rect 42756 16828 42812 16884
rect 42868 16828 42878 16884
rect 46834 16828 46844 16884
rect 46900 16828 47628 16884
rect 47684 16828 47694 16884
rect 53554 16828 53564 16884
rect 53620 16828 54348 16884
rect 54404 16828 54908 16884
rect 54964 16828 54974 16884
rect 55122 16828 55132 16884
rect 55188 16828 55692 16884
rect 55748 16828 56812 16884
rect 56868 16828 56878 16884
rect 1362 16716 1372 16772
rect 1428 16716 2156 16772
rect 2212 16716 2222 16772
rect 7634 16716 7644 16772
rect 7700 16716 8988 16772
rect 9044 16716 9054 16772
rect 9762 16716 9772 16772
rect 9828 16716 10556 16772
rect 10612 16716 10622 16772
rect 14018 16716 14028 16772
rect 14084 16716 14812 16772
rect 14868 16716 14980 16772
rect 20290 16716 20300 16772
rect 20356 16716 23324 16772
rect 23380 16716 23390 16772
rect 25442 16716 25452 16772
rect 25508 16716 26908 16772
rect 29922 16716 29932 16772
rect 29988 16716 32284 16772
rect 32340 16716 32350 16772
rect 36390 16716 36428 16772
rect 36484 16716 36494 16772
rect 36754 16716 36764 16772
rect 36820 16716 40796 16772
rect 40852 16716 40862 16772
rect 41458 16716 41468 16772
rect 41524 16716 42252 16772
rect 42308 16716 42318 16772
rect 43922 16716 43932 16772
rect 43988 16716 45164 16772
rect 45220 16716 46956 16772
rect 47012 16716 47022 16772
rect 47506 16716 47516 16772
rect 47572 16716 48748 16772
rect 48804 16716 48814 16772
rect 48972 16716 50652 16772
rect 50708 16716 50718 16772
rect 51874 16716 51884 16772
rect 51940 16716 52892 16772
rect 52948 16716 52958 16772
rect 7186 16604 7196 16660
rect 7252 16604 8204 16660
rect 8260 16604 8270 16660
rect 9538 16604 9548 16660
rect 9604 16604 9884 16660
rect 9940 16604 9950 16660
rect 21746 16604 21756 16660
rect 21812 16604 22092 16660
rect 22148 16604 27356 16660
rect 27412 16604 27422 16660
rect 28466 16604 28476 16660
rect 28532 16604 34076 16660
rect 34132 16604 34142 16660
rect 35970 16604 35980 16660
rect 36036 16604 44940 16660
rect 44996 16604 45612 16660
rect 45668 16604 45678 16660
rect 46498 16604 46508 16660
rect 46564 16604 48748 16660
rect 48804 16604 48814 16660
rect 48972 16548 49028 16716
rect 49186 16604 49196 16660
rect 49252 16604 52780 16660
rect 52836 16604 53340 16660
rect 53396 16604 53406 16660
rect 18610 16492 18620 16548
rect 18676 16492 19740 16548
rect 19796 16492 20300 16548
rect 20356 16492 20366 16548
rect 24098 16492 24108 16548
rect 24164 16492 25340 16548
rect 25396 16492 25406 16548
rect 40898 16492 40908 16548
rect 40964 16492 49028 16548
rect 8355 16436 8365 16492
rect 8421 16436 8469 16492
rect 8525 16436 8573 16492
rect 8629 16436 8639 16492
rect 22662 16436 22672 16492
rect 22728 16436 22776 16492
rect 22832 16436 22880 16492
rect 22936 16436 22946 16492
rect 36969 16436 36979 16492
rect 37035 16436 37083 16492
rect 37139 16436 37187 16492
rect 37243 16436 37253 16492
rect 51276 16436 51286 16492
rect 51342 16436 51390 16492
rect 51446 16436 51494 16492
rect 51550 16436 51560 16492
rect 29362 16380 29372 16436
rect 29428 16380 34748 16436
rect 34804 16380 34814 16436
rect 46946 16380 46956 16436
rect 47012 16380 48860 16436
rect 48916 16380 50316 16436
rect 50372 16380 50382 16436
rect 4946 16268 4956 16324
rect 5012 16268 6300 16324
rect 6356 16268 6366 16324
rect 8652 16268 9604 16324
rect 10658 16268 10668 16324
rect 10724 16268 24444 16324
rect 24500 16268 24510 16324
rect 30034 16268 30044 16324
rect 30100 16268 31500 16324
rect 31556 16268 31566 16324
rect 36306 16268 36316 16324
rect 36372 16268 38220 16324
rect 38276 16268 38286 16324
rect 42354 16268 42364 16324
rect 42420 16268 42924 16324
rect 42980 16268 42990 16324
rect 44146 16268 44156 16324
rect 44212 16268 51548 16324
rect 51604 16268 51614 16324
rect 8652 16212 8708 16268
rect 9548 16212 9604 16268
rect 3490 16156 3500 16212
rect 3556 16156 8708 16212
rect 8866 16156 8876 16212
rect 8932 16156 9324 16212
rect 9380 16156 9390 16212
rect 9548 16156 13580 16212
rect 13636 16156 14364 16212
rect 14420 16156 14430 16212
rect 17714 16156 17724 16212
rect 17780 16156 24332 16212
rect 24388 16156 24398 16212
rect 25106 16156 25116 16212
rect 25172 16156 25182 16212
rect 28802 16156 28812 16212
rect 28868 16156 30716 16212
rect 30772 16156 30782 16212
rect 36082 16156 36092 16212
rect 36148 16156 38108 16212
rect 38164 16156 40908 16212
rect 40964 16156 40974 16212
rect 47058 16156 47068 16212
rect 47124 16156 48412 16212
rect 48468 16156 48860 16212
rect 48916 16156 49308 16212
rect 49364 16156 49374 16212
rect 4610 16044 4620 16100
rect 4676 16044 6748 16100
rect 6804 16044 8540 16100
rect 8596 16044 9212 16100
rect 9268 16044 9278 16100
rect 11330 16044 11340 16100
rect 11396 16044 12572 16100
rect 12628 16044 12638 16100
rect 20850 16044 20860 16100
rect 20916 16044 21756 16100
rect 21812 16044 21822 16100
rect 23286 16044 23324 16100
rect 23380 16044 23390 16100
rect 0 15988 800 16016
rect 25116 15988 25172 16156
rect 26898 16044 26908 16100
rect 26964 16044 27580 16100
rect 27636 16044 28252 16100
rect 28308 16044 28318 16100
rect 29698 16044 29708 16100
rect 29764 16044 30380 16100
rect 30436 16044 30446 16100
rect 36418 16044 36428 16100
rect 36484 16044 36988 16100
rect 37044 16044 37054 16100
rect 38210 16044 38220 16100
rect 38276 16044 38892 16100
rect 38948 16044 38958 16100
rect 39890 16044 39900 16100
rect 39956 16044 40460 16100
rect 40516 16044 45276 16100
rect 45332 16044 46172 16100
rect 46228 16044 46238 16100
rect 48178 16044 48188 16100
rect 48244 16044 48636 16100
rect 48692 16044 49532 16100
rect 49588 16044 50652 16100
rect 50708 16044 50718 16100
rect 0 15932 1708 15988
rect 1764 15932 5068 15988
rect 5124 15932 5134 15988
rect 7746 15932 7756 15988
rect 7812 15932 8204 15988
rect 8260 15932 8764 15988
rect 8820 15932 10668 15988
rect 10724 15932 10734 15988
rect 12226 15932 12236 15988
rect 12292 15932 14028 15988
rect 14084 15932 14924 15988
rect 14980 15932 14990 15988
rect 16930 15932 16940 15988
rect 16996 15932 22036 15988
rect 22194 15932 22204 15988
rect 22260 15932 23660 15988
rect 23716 15932 23726 15988
rect 25116 15932 31724 15988
rect 31780 15932 31790 15988
rect 32050 15932 32060 15988
rect 32116 15932 32844 15988
rect 32900 15932 32910 15988
rect 36530 15932 36540 15988
rect 36596 15932 37212 15988
rect 37268 15932 37278 15988
rect 0 15904 800 15932
rect 21980 15876 22036 15932
rect 6066 15820 6076 15876
rect 6132 15820 8316 15876
rect 8372 15820 8382 15876
rect 8978 15820 8988 15876
rect 9044 15820 11452 15876
rect 11508 15820 11518 15876
rect 18386 15820 18396 15876
rect 18452 15820 18956 15876
rect 19012 15820 19022 15876
rect 19506 15820 19516 15876
rect 19572 15820 20076 15876
rect 20132 15820 21084 15876
rect 21140 15820 21150 15876
rect 21980 15820 24780 15876
rect 24836 15820 25340 15876
rect 25396 15820 25406 15876
rect 26338 15820 26348 15876
rect 26404 15820 27244 15876
rect 27300 15820 27310 15876
rect 29810 15820 29820 15876
rect 29876 15820 30828 15876
rect 30884 15820 30894 15876
rect 31938 15820 31948 15876
rect 32004 15820 32508 15876
rect 32564 15820 32956 15876
rect 33012 15820 38668 15876
rect 38724 15820 38734 15876
rect 39900 15764 39956 16044
rect 45714 15932 45724 15988
rect 45780 15932 46284 15988
rect 46340 15932 47964 15988
rect 48020 15932 48030 15988
rect 49186 15932 49196 15988
rect 49252 15932 49980 15988
rect 50036 15932 50046 15988
rect 45490 15820 45500 15876
rect 45556 15820 46060 15876
rect 46116 15820 46126 15876
rect 47478 15820 47516 15876
rect 47572 15820 47582 15876
rect 21634 15708 21644 15764
rect 21700 15708 29652 15764
rect 33394 15708 33404 15764
rect 33460 15708 39956 15764
rect 15508 15652 15518 15708
rect 15574 15652 15622 15708
rect 15678 15652 15726 15708
rect 15782 15652 15792 15708
rect 10210 15596 10220 15652
rect 10276 15596 11508 15652
rect 28102 15596 28140 15652
rect 28196 15596 28206 15652
rect 11452 15540 11508 15596
rect 29596 15540 29652 15708
rect 29815 15652 29825 15708
rect 29881 15652 29929 15708
rect 29985 15652 30033 15708
rect 30089 15652 30099 15708
rect 44122 15652 44132 15708
rect 44188 15652 44236 15708
rect 44292 15652 44340 15708
rect 44396 15652 44406 15708
rect 58429 15652 58439 15708
rect 58495 15652 58543 15708
rect 58599 15652 58647 15708
rect 58703 15652 58713 15708
rect 32274 15596 32284 15652
rect 32340 15596 32620 15652
rect 32676 15596 32956 15652
rect 33012 15596 33628 15652
rect 33684 15596 40908 15652
rect 40964 15596 40974 15652
rect 45126 15596 45164 15652
rect 45220 15596 45230 15652
rect 11442 15484 11452 15540
rect 11508 15484 12684 15540
rect 12740 15484 12750 15540
rect 15474 15484 15484 15540
rect 15540 15484 16044 15540
rect 16100 15484 16110 15540
rect 16370 15484 16380 15540
rect 16436 15484 17164 15540
rect 17220 15484 17230 15540
rect 17602 15484 17612 15540
rect 17668 15484 19628 15540
rect 19684 15484 19694 15540
rect 26114 15484 26124 15540
rect 26180 15484 28084 15540
rect 29596 15484 35756 15540
rect 35812 15484 35822 15540
rect 39554 15484 39564 15540
rect 39620 15484 41020 15540
rect 41076 15484 44268 15540
rect 44324 15484 44334 15540
rect 44594 15484 44604 15540
rect 44660 15484 45724 15540
rect 45780 15484 45790 15540
rect 46386 15484 46396 15540
rect 46452 15484 46956 15540
rect 47012 15484 47022 15540
rect 55906 15484 55916 15540
rect 55972 15484 57484 15540
rect 57540 15484 57550 15540
rect 28028 15428 28084 15484
rect 4946 15372 4956 15428
rect 5012 15372 5516 15428
rect 5572 15372 6524 15428
rect 6580 15372 6590 15428
rect 10098 15372 10108 15428
rect 10164 15372 10780 15428
rect 10836 15372 10846 15428
rect 16706 15372 16716 15428
rect 16772 15372 18396 15428
rect 18452 15372 18462 15428
rect 21410 15372 21420 15428
rect 21476 15372 22540 15428
rect 22596 15372 27580 15428
rect 27636 15372 27646 15428
rect 28018 15372 28028 15428
rect 28084 15372 29596 15428
rect 29652 15372 29662 15428
rect 30706 15372 30716 15428
rect 30772 15372 31276 15428
rect 31332 15372 31342 15428
rect 33506 15372 33516 15428
rect 33572 15372 34748 15428
rect 34804 15372 34814 15428
rect 40002 15372 40012 15428
rect 40068 15372 41804 15428
rect 41860 15372 46620 15428
rect 46676 15372 46686 15428
rect 48178 15372 48188 15428
rect 48244 15372 50428 15428
rect 50484 15372 50494 15428
rect 52434 15372 52444 15428
rect 52500 15372 53228 15428
rect 53284 15372 53294 15428
rect 55122 15372 55132 15428
rect 55188 15372 56028 15428
rect 56084 15372 56094 15428
rect 5954 15260 5964 15316
rect 6020 15260 8204 15316
rect 8260 15260 9324 15316
rect 9380 15260 9390 15316
rect 9762 15260 9772 15316
rect 9828 15260 15036 15316
rect 15092 15260 15102 15316
rect 23202 15260 23212 15316
rect 23268 15260 24108 15316
rect 24164 15260 24174 15316
rect 25442 15260 25452 15316
rect 25508 15260 26908 15316
rect 27906 15260 27916 15316
rect 27972 15260 29372 15316
rect 29428 15260 29438 15316
rect 32274 15260 32284 15316
rect 32340 15260 32844 15316
rect 32900 15260 33404 15316
rect 33460 15260 33470 15316
rect 33954 15260 33964 15316
rect 34020 15260 40684 15316
rect 40740 15260 40750 15316
rect 41234 15260 41244 15316
rect 41300 15260 42140 15316
rect 42196 15260 42206 15316
rect 42364 15260 46060 15316
rect 46116 15260 46732 15316
rect 46788 15260 47292 15316
rect 47348 15260 47358 15316
rect 49074 15260 49084 15316
rect 49140 15260 51548 15316
rect 51604 15260 52892 15316
rect 52948 15260 52958 15316
rect 26852 15204 26908 15260
rect 33964 15204 34020 15260
rect 5170 15148 5180 15204
rect 5236 15148 8652 15204
rect 8708 15148 9548 15204
rect 9604 15148 9614 15204
rect 10658 15148 10668 15204
rect 10724 15148 11564 15204
rect 11620 15148 11630 15204
rect 12338 15148 12348 15204
rect 12404 15148 13804 15204
rect 13860 15148 13870 15204
rect 14578 15148 14588 15204
rect 14644 15148 14924 15204
rect 14980 15148 17724 15204
rect 17780 15148 17790 15204
rect 22754 15148 22764 15204
rect 22820 15148 23100 15204
rect 23156 15148 23166 15204
rect 25106 15148 25116 15204
rect 25172 15148 26012 15204
rect 26068 15148 26078 15204
rect 26852 15148 27356 15204
rect 27412 15148 34020 15204
rect 40684 15204 40740 15260
rect 42364 15204 42420 15260
rect 40684 15148 42420 15204
rect 42476 15148 43820 15204
rect 43876 15148 43886 15204
rect 51650 15148 51660 15204
rect 51716 15148 52556 15204
rect 52612 15148 52622 15204
rect 52770 15148 52780 15204
rect 52836 15148 54796 15204
rect 54852 15148 55804 15204
rect 55860 15148 55870 15204
rect 56130 15148 56140 15204
rect 56196 15148 57708 15204
rect 57764 15148 57774 15204
rect 12114 15092 12124 15148
rect 12180 15092 12190 15148
rect 42476 15092 42532 15148
rect 1036 15036 1820 15092
rect 1876 15036 5628 15092
rect 5684 15036 5694 15092
rect 7298 15036 7308 15092
rect 7364 15036 7980 15092
rect 8036 15036 8046 15092
rect 8204 15036 9772 15092
rect 9828 15036 9838 15092
rect 12124 15036 12684 15092
rect 12740 15036 12750 15092
rect 14018 15036 14028 15092
rect 14084 15036 14700 15092
rect 14756 15036 14766 15092
rect 18610 15036 18620 15092
rect 18676 15036 27804 15092
rect 27860 15036 27870 15092
rect 42466 15036 42476 15092
rect 42532 15036 42542 15092
rect 46946 15036 46956 15092
rect 47012 15036 48636 15092
rect 48692 15036 48702 15092
rect 0 14868 800 14896
rect 1036 14868 1092 15036
rect 2370 14924 2380 14980
rect 2436 14924 6636 14980
rect 6692 14924 6702 14980
rect 8204 14868 8260 15036
rect 8950 14924 8988 14980
rect 9044 14924 9054 14980
rect 20178 14924 20188 14980
rect 20244 14924 21644 14980
rect 21700 14924 21710 14980
rect 23426 14924 23436 14980
rect 23492 14924 35644 14980
rect 35700 14924 35710 14980
rect 39330 14924 39340 14980
rect 39396 14924 49868 14980
rect 49924 14924 50652 14980
rect 50708 14924 50718 14980
rect 8355 14868 8365 14924
rect 8421 14868 8469 14924
rect 8525 14868 8573 14924
rect 8629 14868 8639 14924
rect 22662 14868 22672 14924
rect 22728 14868 22776 14924
rect 22832 14868 22880 14924
rect 22936 14868 22946 14924
rect 36969 14868 36979 14924
rect 37035 14868 37083 14924
rect 37139 14868 37187 14924
rect 37243 14868 37253 14924
rect 51276 14868 51286 14924
rect 51342 14868 51390 14924
rect 51446 14868 51494 14924
rect 51550 14868 51560 14924
rect 0 14812 1092 14868
rect 4284 14812 8260 14868
rect 8764 14812 10556 14868
rect 10612 14812 10622 14868
rect 23090 14812 23100 14868
rect 23156 14812 25900 14868
rect 25956 14812 28588 14868
rect 28644 14812 28654 14868
rect 0 14784 800 14812
rect 3500 14700 3948 14756
rect 4004 14700 4014 14756
rect 3500 14644 3556 14700
rect 4284 14644 4340 14812
rect 8764 14756 8820 14812
rect 4498 14700 4508 14756
rect 4564 14700 8820 14756
rect 8978 14700 8988 14756
rect 9044 14700 9884 14756
rect 9940 14700 11228 14756
rect 11284 14700 11294 14756
rect 26898 14700 26908 14756
rect 26964 14700 26974 14756
rect 27794 14700 27804 14756
rect 27860 14700 37324 14756
rect 37380 14700 38556 14756
rect 38612 14700 38622 14756
rect 38882 14700 38892 14756
rect 38948 14700 40236 14756
rect 40292 14700 40302 14756
rect 50372 14700 51100 14756
rect 51156 14700 51166 14756
rect 26908 14644 26964 14700
rect 50372 14644 50428 14700
rect 3490 14588 3500 14644
rect 3556 14588 3566 14644
rect 4050 14588 4060 14644
rect 4116 14588 4284 14644
rect 4340 14588 4350 14644
rect 5516 14588 6972 14644
rect 7028 14588 8092 14644
rect 8148 14588 8158 14644
rect 14578 14588 14588 14644
rect 14644 14588 15932 14644
rect 15988 14588 17052 14644
rect 17108 14588 17118 14644
rect 21746 14588 21756 14644
rect 21812 14588 26124 14644
rect 26180 14588 26572 14644
rect 26628 14588 26638 14644
rect 26908 14588 33908 14644
rect 36194 14588 36204 14644
rect 36260 14588 43932 14644
rect 43988 14588 43998 14644
rect 45490 14588 45500 14644
rect 45556 14588 46620 14644
rect 46676 14588 46956 14644
rect 47012 14588 47022 14644
rect 50194 14588 50204 14644
rect 50260 14588 50428 14644
rect 54898 14588 54908 14644
rect 54964 14588 56140 14644
rect 56196 14588 56206 14644
rect 3378 14476 3388 14532
rect 3444 14476 4396 14532
rect 4452 14476 4844 14532
rect 4900 14476 4910 14532
rect 5516 14420 5572 14588
rect 33852 14532 33908 14588
rect 5730 14476 5740 14532
rect 5796 14476 7644 14532
rect 7700 14476 7710 14532
rect 7858 14476 7868 14532
rect 7924 14476 9884 14532
rect 9940 14476 9950 14532
rect 10210 14476 10220 14532
rect 10276 14476 10668 14532
rect 10724 14476 11564 14532
rect 11620 14476 11630 14532
rect 11778 14476 11788 14532
rect 11844 14476 12124 14532
rect 12180 14476 12190 14532
rect 14690 14476 14700 14532
rect 14756 14476 18284 14532
rect 18340 14476 18350 14532
rect 21298 14476 21308 14532
rect 21364 14476 22652 14532
rect 22708 14476 22718 14532
rect 23090 14476 23100 14532
rect 23156 14476 24556 14532
rect 24612 14476 25452 14532
rect 25508 14476 25518 14532
rect 25676 14476 30492 14532
rect 30548 14476 30558 14532
rect 33852 14476 37100 14532
rect 37156 14476 37660 14532
rect 37716 14476 37726 14532
rect 38658 14476 38668 14532
rect 38724 14476 39340 14532
rect 39396 14476 39406 14532
rect 39666 14476 39676 14532
rect 39732 14476 39742 14532
rect 40338 14476 40348 14532
rect 40404 14476 41132 14532
rect 41188 14476 41198 14532
rect 44258 14476 44268 14532
rect 44324 14476 46172 14532
rect 46228 14476 46238 14532
rect 48066 14476 48076 14532
rect 48132 14476 48748 14532
rect 48804 14476 48814 14532
rect 51986 14476 51996 14532
rect 52052 14476 55804 14532
rect 55860 14476 56252 14532
rect 56308 14476 56318 14532
rect 25676 14420 25732 14476
rect 1138 14364 1148 14420
rect 1204 14364 2716 14420
rect 2772 14364 2782 14420
rect 4946 14364 4956 14420
rect 5012 14364 5572 14420
rect 7298 14364 7308 14420
rect 7364 14364 8764 14420
rect 8820 14364 8830 14420
rect 10994 14364 11004 14420
rect 11060 14364 12572 14420
rect 12628 14364 12638 14420
rect 14102 14364 14140 14420
rect 14196 14364 15036 14420
rect 15092 14364 15102 14420
rect 15250 14364 15260 14420
rect 15316 14364 15932 14420
rect 15988 14364 16268 14420
rect 16324 14364 16334 14420
rect 21186 14364 21196 14420
rect 21252 14364 25732 14420
rect 26562 14364 26572 14420
rect 26628 14364 27916 14420
rect 27972 14364 28476 14420
rect 28532 14364 28542 14420
rect 34962 14364 34972 14420
rect 35028 14364 35196 14420
rect 35252 14364 39228 14420
rect 39284 14364 39294 14420
rect 39676 14308 39732 14476
rect 48290 14364 48300 14420
rect 48356 14364 48860 14420
rect 48916 14364 48926 14420
rect 1474 14252 1484 14308
rect 1540 14252 2044 14308
rect 2100 14252 2110 14308
rect 3826 14252 3836 14308
rect 3892 14252 4508 14308
rect 4564 14252 4574 14308
rect 6066 14252 6076 14308
rect 6132 14252 7980 14308
rect 8036 14252 8046 14308
rect 10098 14252 10108 14308
rect 10164 14252 11340 14308
rect 11396 14252 13692 14308
rect 13748 14252 13758 14308
rect 16370 14252 16380 14308
rect 16436 14252 17612 14308
rect 17668 14252 17678 14308
rect 20626 14252 20636 14308
rect 20692 14252 22988 14308
rect 23044 14252 23054 14308
rect 24658 14252 24668 14308
rect 24724 14252 25228 14308
rect 25284 14252 25294 14308
rect 26450 14252 26460 14308
rect 26516 14252 28252 14308
rect 28308 14252 28318 14308
rect 28578 14252 28588 14308
rect 28644 14252 29932 14308
rect 29988 14252 29998 14308
rect 31602 14252 31612 14308
rect 31668 14252 32508 14308
rect 32564 14252 32574 14308
rect 33058 14252 33068 14308
rect 33124 14252 34076 14308
rect 34132 14252 34142 14308
rect 34626 14252 34636 14308
rect 34692 14252 35644 14308
rect 35700 14252 35710 14308
rect 38770 14252 38780 14308
rect 38836 14252 39732 14308
rect 48178 14252 48188 14308
rect 48244 14252 49644 14308
rect 49700 14252 49710 14308
rect 25228 14196 25284 14252
rect 16146 14140 16156 14196
rect 16212 14140 20188 14196
rect 20244 14140 20254 14196
rect 25228 14140 26684 14196
rect 26740 14140 26750 14196
rect 42774 14140 42812 14196
rect 42868 14140 42878 14196
rect 48290 14140 48300 14196
rect 48356 14140 52444 14196
rect 52500 14140 52510 14196
rect 57250 14140 57260 14196
rect 57316 14140 57820 14196
rect 57876 14140 57886 14196
rect 15508 14084 15518 14140
rect 15574 14084 15622 14140
rect 15678 14084 15726 14140
rect 15782 14084 15792 14140
rect 29815 14084 29825 14140
rect 29881 14084 29929 14140
rect 29985 14084 30033 14140
rect 30089 14084 30099 14140
rect 44122 14084 44132 14140
rect 44188 14084 44236 14140
rect 44292 14084 44340 14140
rect 44396 14084 44406 14140
rect 58429 14084 58439 14140
rect 58495 14084 58543 14140
rect 58599 14084 58647 14140
rect 58703 14084 58713 14140
rect 3332 14028 4508 14084
rect 4564 14028 4574 14084
rect 6402 14028 6412 14084
rect 6468 14028 7644 14084
rect 7700 14028 7710 14084
rect 25778 14028 25788 14084
rect 25844 14028 26348 14084
rect 26404 14028 27356 14084
rect 27412 14028 27422 14084
rect 32162 14028 32172 14084
rect 32228 14028 35420 14084
rect 35476 14028 35486 14084
rect 3332 13972 3388 14028
rect 2006 13916 2044 13972
rect 2100 13916 3388 13972
rect 3490 13916 3500 13972
rect 3556 13916 3594 13972
rect 5628 13916 16604 13972
rect 16660 13916 16670 13972
rect 23538 13916 23548 13972
rect 23604 13916 25228 13972
rect 25284 13916 29148 13972
rect 29204 13916 30268 13972
rect 30324 13916 30716 13972
rect 30772 13916 30782 13972
rect 33730 13916 33740 13972
rect 33796 13916 34412 13972
rect 34468 13916 34478 13972
rect 2146 13804 2156 13860
rect 2212 13804 2548 13860
rect 2706 13804 2716 13860
rect 2772 13804 3724 13860
rect 3780 13804 3790 13860
rect 0 13748 800 13776
rect 2492 13748 2548 13804
rect 5628 13748 5684 13916
rect 7298 13804 7308 13860
rect 7364 13804 10556 13860
rect 10612 13804 10622 13860
rect 11554 13804 11564 13860
rect 11620 13804 13356 13860
rect 13412 13804 13422 13860
rect 22194 13804 22204 13860
rect 22260 13804 23884 13860
rect 23940 13804 24668 13860
rect 24724 13804 24734 13860
rect 29362 13804 29372 13860
rect 29428 13804 30156 13860
rect 30212 13804 30940 13860
rect 30996 13804 31006 13860
rect 32172 13804 35420 13860
rect 35476 13804 35486 13860
rect 36418 13804 36428 13860
rect 36484 13804 37436 13860
rect 37492 13804 37502 13860
rect 42914 13804 42924 13860
rect 42980 13804 43484 13860
rect 43540 13804 43550 13860
rect 44930 13804 44940 13860
rect 44996 13804 45276 13860
rect 45332 13804 47292 13860
rect 47348 13804 50428 13860
rect 50484 13804 50494 13860
rect 52994 13804 53004 13860
rect 53060 13804 54908 13860
rect 54964 13804 54974 13860
rect 32172 13748 32228 13804
rect 0 13692 2268 13748
rect 2324 13692 2334 13748
rect 2492 13692 2940 13748
rect 2996 13692 5684 13748
rect 5842 13692 5852 13748
rect 5908 13692 9548 13748
rect 9604 13692 9614 13748
rect 12786 13692 12796 13748
rect 12852 13692 13692 13748
rect 13748 13692 13758 13748
rect 15138 13692 15148 13748
rect 15204 13692 16268 13748
rect 16324 13692 16334 13748
rect 16594 13692 16604 13748
rect 16660 13692 18956 13748
rect 19012 13692 19022 13748
rect 23426 13692 23436 13748
rect 23492 13692 24220 13748
rect 24276 13692 24286 13748
rect 26852 13692 32228 13748
rect 32284 13692 33628 13748
rect 33684 13692 34244 13748
rect 0 13664 800 13692
rect 26852 13636 26908 13692
rect 32284 13636 32340 13692
rect 34188 13636 34244 13692
rect 5282 13580 5292 13636
rect 5348 13580 6300 13636
rect 6356 13580 6366 13636
rect 7074 13580 7084 13636
rect 7140 13580 8092 13636
rect 8148 13580 10108 13636
rect 10164 13580 10174 13636
rect 11554 13580 11564 13636
rect 11620 13580 14700 13636
rect 14756 13580 14766 13636
rect 17938 13580 17948 13636
rect 18004 13580 18676 13636
rect 20514 13580 20524 13636
rect 20580 13580 20972 13636
rect 21028 13580 21420 13636
rect 21476 13580 26908 13636
rect 30930 13580 30940 13636
rect 30996 13580 32060 13636
rect 32116 13580 32126 13636
rect 32274 13580 32284 13636
rect 32340 13580 32350 13636
rect 32498 13580 32508 13636
rect 32564 13580 33404 13636
rect 33460 13580 33964 13636
rect 34020 13580 34030 13636
rect 34178 13580 34188 13636
rect 34244 13580 34254 13636
rect 39778 13580 39788 13636
rect 39844 13580 41132 13636
rect 41188 13580 41198 13636
rect 43474 13580 43484 13636
rect 43540 13580 47516 13636
rect 47572 13580 47582 13636
rect 48290 13580 48300 13636
rect 48356 13580 50316 13636
rect 50372 13580 50382 13636
rect 51762 13580 51772 13636
rect 51828 13580 53340 13636
rect 53396 13580 53406 13636
rect 18620 13524 18676 13580
rect 4844 13468 5852 13524
rect 5908 13468 8428 13524
rect 8484 13468 8494 13524
rect 9090 13468 9100 13524
rect 9156 13468 9772 13524
rect 9828 13468 9838 13524
rect 10882 13468 10892 13524
rect 10948 13468 11228 13524
rect 11284 13468 11294 13524
rect 14354 13468 14364 13524
rect 14420 13468 16828 13524
rect 16884 13468 18172 13524
rect 18228 13468 18238 13524
rect 18610 13468 18620 13524
rect 18676 13468 21868 13524
rect 21924 13468 21934 13524
rect 24434 13468 24444 13524
rect 24500 13468 24780 13524
rect 24836 13468 24846 13524
rect 31490 13468 31500 13524
rect 31556 13468 32396 13524
rect 32452 13468 33292 13524
rect 33348 13468 33358 13524
rect 39330 13468 39340 13524
rect 39396 13468 40012 13524
rect 40068 13468 42476 13524
rect 42532 13468 42542 13524
rect 43922 13468 43932 13524
rect 43988 13468 45612 13524
rect 45668 13468 45678 13524
rect 4844 13412 4900 13468
rect 15820 13412 15876 13468
rect 41356 13412 41412 13468
rect 4834 13356 4844 13412
rect 4900 13356 4910 13412
rect 7970 13356 7980 13412
rect 8036 13356 8046 13412
rect 12338 13356 12348 13412
rect 12404 13356 12460 13412
rect 12516 13356 12526 13412
rect 15810 13356 15820 13412
rect 15876 13356 15886 13412
rect 16370 13356 16380 13412
rect 16436 13356 17500 13412
rect 17556 13356 17566 13412
rect 23314 13356 23324 13412
rect 23380 13356 24892 13412
rect 24948 13356 24958 13412
rect 30370 13356 30380 13412
rect 30436 13356 31724 13412
rect 31780 13356 31790 13412
rect 41346 13356 41356 13412
rect 41412 13356 41422 13412
rect 46274 13356 46284 13412
rect 46340 13356 48188 13412
rect 48244 13356 49420 13412
rect 49476 13356 49486 13412
rect 7980 13188 8036 13356
rect 8355 13300 8365 13356
rect 8421 13300 8469 13356
rect 8525 13300 8573 13356
rect 8629 13300 8639 13356
rect 16380 13300 16436 13356
rect 22662 13300 22672 13356
rect 22728 13300 22776 13356
rect 22832 13300 22880 13356
rect 22936 13300 22946 13356
rect 36969 13300 36979 13356
rect 37035 13300 37083 13356
rect 37139 13300 37187 13356
rect 37243 13300 37253 13356
rect 51276 13300 51286 13356
rect 51342 13300 51390 13356
rect 51446 13300 51494 13356
rect 51550 13300 51560 13356
rect 12114 13244 12124 13300
rect 12180 13244 12572 13300
rect 12628 13244 13804 13300
rect 13860 13244 16436 13300
rect 23426 13244 23436 13300
rect 23492 13244 32788 13300
rect 43586 13244 43596 13300
rect 43652 13244 44268 13300
rect 44324 13244 47852 13300
rect 47908 13244 48860 13300
rect 48916 13244 48926 13300
rect 57362 13244 57372 13300
rect 57428 13244 58044 13300
rect 58100 13244 58110 13300
rect 32732 13188 32788 13244
rect 7980 13132 8316 13188
rect 8372 13132 8382 13188
rect 11218 13132 11228 13188
rect 11284 13132 15372 13188
rect 15428 13132 15438 13188
rect 22082 13132 22092 13188
rect 22148 13132 26908 13188
rect 26964 13132 30156 13188
rect 30212 13132 31388 13188
rect 31444 13132 31454 13188
rect 32732 13132 50428 13188
rect 57474 13132 57484 13188
rect 57540 13132 57820 13188
rect 57876 13132 57886 13188
rect 50372 13076 50428 13132
rect 15092 13020 16156 13076
rect 16212 13020 16222 13076
rect 16594 13020 16604 13076
rect 16660 13020 17164 13076
rect 17220 13020 17230 13076
rect 21074 13020 21084 13076
rect 21140 13020 23436 13076
rect 23492 13020 23502 13076
rect 23660 13020 41916 13076
rect 41972 13020 41982 13076
rect 44706 13020 44716 13076
rect 44772 13020 45164 13076
rect 45220 13020 48300 13076
rect 48356 13020 48366 13076
rect 50372 13020 55468 13076
rect 55524 13020 55534 13076
rect 15092 12964 15148 13020
rect 23660 12964 23716 13020
rect 3042 12908 3052 12964
rect 3108 12908 4228 12964
rect 4172 12852 4228 12908
rect 5516 12908 15148 12964
rect 21746 12908 21756 12964
rect 21812 12908 23716 12964
rect 24658 12908 24668 12964
rect 24724 12908 25676 12964
rect 25732 12908 25742 12964
rect 26226 12908 26236 12964
rect 26292 12908 27132 12964
rect 27188 12908 27198 12964
rect 31154 12908 31164 12964
rect 31220 12908 34860 12964
rect 34916 12908 34926 12964
rect 37650 12908 37660 12964
rect 37716 12908 38556 12964
rect 38612 12908 38622 12964
rect 46022 12908 46060 12964
rect 46116 12908 46126 12964
rect 46386 12908 46396 12964
rect 46452 12908 46844 12964
rect 46900 12908 46910 12964
rect 49522 12908 49532 12964
rect 49588 12908 50540 12964
rect 50596 12908 50764 12964
rect 50820 12908 50830 12964
rect 1250 12796 1260 12852
rect 1316 12796 2380 12852
rect 2436 12796 2446 12852
rect 3490 12796 3500 12852
rect 3556 12796 3566 12852
rect 3714 12796 3724 12852
rect 3780 12796 3818 12852
rect 4162 12796 4172 12852
rect 4228 12796 4238 12852
rect 3500 12740 3556 12796
rect 5516 12740 5572 12908
rect 5730 12796 5740 12852
rect 5796 12796 6636 12852
rect 6692 12796 7868 12852
rect 7924 12796 7934 12852
rect 9202 12796 9212 12852
rect 9268 12796 11676 12852
rect 11732 12796 11742 12852
rect 15092 12796 15596 12852
rect 15652 12796 16492 12852
rect 16548 12796 16558 12852
rect 25106 12796 25116 12852
rect 25172 12796 25900 12852
rect 25956 12796 25966 12852
rect 30930 12796 30940 12852
rect 30996 12796 33964 12852
rect 34020 12796 34972 12852
rect 35028 12796 35038 12852
rect 40002 12796 40012 12852
rect 40068 12796 41132 12852
rect 41188 12796 41198 12852
rect 46162 12796 46172 12852
rect 46228 12796 51100 12852
rect 51156 12796 51166 12852
rect 15092 12740 15148 12796
rect 3042 12684 3052 12740
rect 3108 12684 4844 12740
rect 4900 12684 5572 12740
rect 6738 12684 6748 12740
rect 6804 12684 8988 12740
rect 9044 12684 10892 12740
rect 10948 12684 11228 12740
rect 11284 12684 11294 12740
rect 13010 12684 13020 12740
rect 13076 12684 14252 12740
rect 14308 12684 15148 12740
rect 15698 12684 15708 12740
rect 15764 12684 17612 12740
rect 17668 12684 17678 12740
rect 20626 12684 20636 12740
rect 20692 12684 22204 12740
rect 22260 12684 22270 12740
rect 22418 12684 22428 12740
rect 22484 12684 23884 12740
rect 23940 12684 23950 12740
rect 27458 12684 27468 12740
rect 27524 12684 28028 12740
rect 28084 12684 28094 12740
rect 29586 12684 29596 12740
rect 29652 12684 30604 12740
rect 30660 12684 30670 12740
rect 0 12628 800 12656
rect 0 12572 1708 12628
rect 1764 12572 1774 12628
rect 5506 12572 5516 12628
rect 5572 12572 13468 12628
rect 13524 12572 13534 12628
rect 16482 12572 16492 12628
rect 16548 12572 19740 12628
rect 19796 12572 19806 12628
rect 21858 12572 21868 12628
rect 21924 12572 23436 12628
rect 23492 12572 29372 12628
rect 29428 12572 29438 12628
rect 31826 12572 31836 12628
rect 31892 12572 34860 12628
rect 34916 12572 34926 12628
rect 0 12544 800 12572
rect 15508 12516 15518 12572
rect 15574 12516 15622 12572
rect 15678 12516 15726 12572
rect 15782 12516 15792 12572
rect 29815 12516 29825 12572
rect 29881 12516 29929 12572
rect 29985 12516 30033 12572
rect 30089 12516 30099 12572
rect 44122 12516 44132 12572
rect 44188 12516 44236 12572
rect 44292 12516 44340 12572
rect 44396 12516 44406 12572
rect 46172 12516 46228 12796
rect 58429 12516 58439 12572
rect 58495 12516 58543 12572
rect 58599 12516 58647 12572
rect 58703 12516 58713 12572
rect 9538 12460 9548 12516
rect 9604 12460 9614 12516
rect 17836 12460 26796 12516
rect 9548 12404 9604 12460
rect 4722 12348 4732 12404
rect 4788 12348 8092 12404
rect 8148 12348 9604 12404
rect 11890 12348 11900 12404
rect 11956 12348 12572 12404
rect 12628 12348 12638 12404
rect 13794 12348 13804 12404
rect 13860 12348 15820 12404
rect 15876 12348 15886 12404
rect 17836 12292 17892 12460
rect 26852 12404 26908 12516
rect 27010 12460 27020 12516
rect 27076 12460 29204 12516
rect 19730 12348 19740 12404
rect 19796 12348 20636 12404
rect 20692 12348 20702 12404
rect 26852 12348 28924 12404
rect 28980 12348 28990 12404
rect 29148 12292 29204 12460
rect 44828 12460 45164 12516
rect 45220 12460 46228 12516
rect 44828 12404 44884 12460
rect 44034 12348 44044 12404
rect 44100 12348 44884 12404
rect 45042 12348 45052 12404
rect 45108 12348 47180 12404
rect 47236 12348 47246 12404
rect 3714 12236 3724 12292
rect 3780 12236 5180 12292
rect 5236 12236 5246 12292
rect 15586 12236 15596 12292
rect 15652 12236 17836 12292
rect 17892 12236 17902 12292
rect 18050 12236 18060 12292
rect 18116 12236 19852 12292
rect 19908 12236 19918 12292
rect 21970 12236 21980 12292
rect 22036 12236 22428 12292
rect 22484 12236 22494 12292
rect 24546 12236 24556 12292
rect 24612 12236 25340 12292
rect 25396 12236 25406 12292
rect 27122 12236 27132 12292
rect 27188 12236 27804 12292
rect 27860 12236 27870 12292
rect 29148 12236 33236 12292
rect 40114 12236 40124 12292
rect 40180 12236 41132 12292
rect 41188 12236 41198 12292
rect 44706 12236 44716 12292
rect 44772 12236 45388 12292
rect 45444 12236 45454 12292
rect 45602 12236 45612 12292
rect 45668 12236 46452 12292
rect 46834 12236 46844 12292
rect 46900 12236 51212 12292
rect 51268 12236 52108 12292
rect 52164 12236 52174 12292
rect 55234 12236 55244 12292
rect 55300 12236 56140 12292
rect 56196 12236 56206 12292
rect 56578 12236 56588 12292
rect 56644 12236 57148 12292
rect 57204 12236 57214 12292
rect 15250 12124 15260 12180
rect 15316 12124 16828 12180
rect 16884 12124 17388 12180
rect 17444 12124 17454 12180
rect 18620 12124 20188 12180
rect 20244 12124 20254 12180
rect 23538 12124 23548 12180
rect 23604 12124 24332 12180
rect 24388 12124 24398 12180
rect 25890 12124 25900 12180
rect 25956 12124 27916 12180
rect 27972 12124 27982 12180
rect 28242 12124 28252 12180
rect 28308 12124 29484 12180
rect 29540 12124 29550 12180
rect 30706 12124 30716 12180
rect 30772 12124 31388 12180
rect 31444 12124 31454 12180
rect 18620 12068 18676 12124
rect 30716 12068 30772 12124
rect 33180 12068 33236 12236
rect 46396 12180 46452 12236
rect 35634 12124 35644 12180
rect 35700 12124 36764 12180
rect 36820 12124 37660 12180
rect 37716 12124 37726 12180
rect 45266 12124 45276 12180
rect 45332 12124 45836 12180
rect 45892 12124 45902 12180
rect 46386 12124 46396 12180
rect 46452 12124 46462 12180
rect 5170 12012 5180 12068
rect 5236 12012 5740 12068
rect 5796 12012 5806 12068
rect 14802 12012 14812 12068
rect 14868 12012 16604 12068
rect 16660 12012 18676 12068
rect 18834 12012 18844 12068
rect 18900 12012 20860 12068
rect 20916 12012 20926 12068
rect 24434 12012 24444 12068
rect 24500 12012 26124 12068
rect 26180 12012 26190 12068
rect 26450 12012 26460 12068
rect 26516 12012 27020 12068
rect 27076 12012 27086 12068
rect 27570 12012 27580 12068
rect 27636 12012 28364 12068
rect 28420 12012 30772 12068
rect 33170 12012 33180 12068
rect 33236 12012 33964 12068
rect 34020 12012 34412 12068
rect 34468 12012 34860 12068
rect 34916 12012 34926 12068
rect 36306 12012 36316 12068
rect 36372 12012 37884 12068
rect 37940 12012 37950 12068
rect 39330 12012 39340 12068
rect 39396 12012 41020 12068
rect 41076 12012 41086 12068
rect 42914 12012 42924 12068
rect 42980 12012 43820 12068
rect 43876 12012 44380 12068
rect 44436 12012 46172 12068
rect 46228 12012 47068 12068
rect 47124 12012 47134 12068
rect 47394 12012 47404 12068
rect 47460 12012 51100 12068
rect 51156 12012 51772 12068
rect 51828 12012 51838 12068
rect 55570 12012 55580 12068
rect 55636 12012 56812 12068
rect 56868 12012 57372 12068
rect 57428 12012 57438 12068
rect 9090 11900 9100 11956
rect 9156 11900 12404 11956
rect 18162 11900 18172 11956
rect 18228 11900 19964 11956
rect 20020 11900 20030 11956
rect 20290 11900 20300 11956
rect 20356 11900 21756 11956
rect 21812 11900 23212 11956
rect 23268 11900 23278 11956
rect 26226 11900 26236 11956
rect 26292 11900 32004 11956
rect 32162 11900 32172 11956
rect 32228 11900 33068 11956
rect 33124 11900 33852 11956
rect 33908 11900 33918 11956
rect 45378 11900 45388 11956
rect 45444 11900 45612 11956
rect 45668 11900 45678 11956
rect 45826 11900 45836 11956
rect 45892 11900 46340 11956
rect 46498 11900 46508 11956
rect 46564 11900 47180 11956
rect 47236 11900 47246 11956
rect 50754 11900 50764 11956
rect 50820 11900 51436 11956
rect 51492 11900 52332 11956
rect 52388 11900 52398 11956
rect 54898 11900 54908 11956
rect 54964 11900 57204 11956
rect 12348 11844 12404 11900
rect 31948 11844 32004 11900
rect 46284 11844 46340 11900
rect 57148 11844 57204 11900
rect 5058 11788 5068 11844
rect 5124 11788 5516 11844
rect 5572 11788 5582 11844
rect 11554 11788 11564 11844
rect 11620 11788 11844 11844
rect 12338 11788 12348 11844
rect 12404 11788 12414 11844
rect 18610 11788 18620 11844
rect 18676 11788 18956 11844
rect 19012 11788 19908 11844
rect 20066 11788 20076 11844
rect 20132 11788 22540 11844
rect 22596 11788 22606 11844
rect 26898 11788 26908 11844
rect 26964 11788 27692 11844
rect 27748 11788 27758 11844
rect 31948 11788 32508 11844
rect 32564 11788 32574 11844
rect 39218 11788 39228 11844
rect 39284 11788 42476 11844
rect 42532 11788 42542 11844
rect 46022 11788 46060 11844
rect 46116 11788 46126 11844
rect 46284 11788 46620 11844
rect 46676 11788 46686 11844
rect 56130 11788 56140 11844
rect 56196 11788 56812 11844
rect 56868 11788 56878 11844
rect 57138 11788 57148 11844
rect 57204 11788 57820 11844
rect 57876 11788 57886 11844
rect 8355 11732 8365 11788
rect 8421 11732 8469 11788
rect 8525 11732 8573 11788
rect 8629 11732 8639 11788
rect 11788 11732 11844 11788
rect 19852 11732 19908 11788
rect 22662 11732 22672 11788
rect 22728 11732 22776 11788
rect 22832 11732 22880 11788
rect 22936 11732 22946 11788
rect 36969 11732 36979 11788
rect 37035 11732 37083 11788
rect 37139 11732 37187 11788
rect 37243 11732 37253 11788
rect 41244 11732 41300 11788
rect 51276 11732 51286 11788
rect 51342 11732 51390 11788
rect 51446 11732 51494 11788
rect 51550 11732 51560 11788
rect 1708 11676 1932 11732
rect 1988 11676 1998 11732
rect 6290 11676 6300 11732
rect 6356 11676 7084 11732
rect 7140 11676 7644 11732
rect 7700 11676 7710 11732
rect 11788 11676 14364 11732
rect 14420 11676 14430 11732
rect 16930 11676 16940 11732
rect 16996 11676 19068 11732
rect 19124 11676 19134 11732
rect 19852 11676 20300 11732
rect 20356 11676 20366 11732
rect 23100 11676 32788 11732
rect 34066 11676 34076 11732
rect 34132 11676 34300 11732
rect 34356 11676 34366 11732
rect 41234 11676 41244 11732
rect 41300 11676 41310 11732
rect 42018 11676 42028 11732
rect 42084 11676 43596 11732
rect 43652 11676 43662 11732
rect 45714 11676 45724 11732
rect 45780 11676 46284 11732
rect 46340 11676 46350 11732
rect 49410 11676 49420 11732
rect 49476 11676 50092 11732
rect 50148 11676 50652 11732
rect 50708 11676 50718 11732
rect 0 11508 800 11536
rect 0 11452 980 11508
rect 0 11424 800 11452
rect 924 11396 980 11452
rect 1708 11396 1764 11676
rect 23100 11620 23156 11676
rect 32732 11620 32788 11676
rect 3602 11564 3612 11620
rect 3668 11564 4732 11620
rect 4788 11564 10444 11620
rect 10500 11564 10510 11620
rect 14130 11564 14140 11620
rect 14196 11564 14206 11620
rect 20178 11564 20188 11620
rect 20244 11564 20748 11620
rect 20804 11564 23156 11620
rect 27010 11564 27020 11620
rect 27076 11564 28588 11620
rect 28644 11564 29820 11620
rect 29876 11564 31500 11620
rect 31556 11564 31566 11620
rect 32732 11564 48748 11620
rect 48804 11564 48814 11620
rect 1922 11452 1932 11508
rect 1988 11452 3052 11508
rect 3108 11452 4060 11508
rect 4116 11452 9268 11508
rect 9212 11396 9268 11452
rect 14140 11396 14196 11564
rect 17938 11452 17948 11508
rect 18004 11452 19740 11508
rect 19796 11452 20524 11508
rect 20580 11452 20590 11508
rect 20850 11452 20860 11508
rect 20916 11452 22036 11508
rect 26002 11452 26012 11508
rect 26068 11452 26684 11508
rect 26740 11452 26750 11508
rect 27010 11452 27020 11508
rect 27076 11452 29596 11508
rect 29652 11452 30380 11508
rect 30436 11452 30446 11508
rect 30930 11452 30940 11508
rect 30996 11452 31836 11508
rect 31892 11452 31902 11508
rect 32386 11452 32396 11508
rect 32452 11452 33628 11508
rect 33684 11452 33694 11508
rect 37986 11452 37996 11508
rect 38052 11452 39564 11508
rect 39620 11452 39630 11508
rect 46946 11452 46956 11508
rect 47012 11452 47964 11508
rect 48020 11452 48030 11508
rect 21980 11396 22036 11452
rect 924 11340 2156 11396
rect 2212 11340 2222 11396
rect 2482 11340 2492 11396
rect 2548 11340 2558 11396
rect 3378 11340 3388 11396
rect 3444 11340 5628 11396
rect 5684 11340 5964 11396
rect 6020 11340 6636 11396
rect 6692 11340 6702 11396
rect 9202 11340 9212 11396
rect 9268 11340 9884 11396
rect 9940 11340 9950 11396
rect 12338 11340 12348 11396
rect 12404 11340 14196 11396
rect 14354 11340 14364 11396
rect 14420 11340 16940 11396
rect 16996 11340 17006 11396
rect 17826 11340 17836 11396
rect 17892 11340 19964 11396
rect 20020 11340 21308 11396
rect 21364 11340 21374 11396
rect 21970 11340 21980 11396
rect 22036 11340 22764 11396
rect 22820 11340 22830 11396
rect 24546 11340 24556 11396
rect 24612 11340 25228 11396
rect 25284 11340 25294 11396
rect 26898 11340 26908 11396
rect 26964 11340 26974 11396
rect 27122 11340 27132 11396
rect 27188 11340 28140 11396
rect 28196 11340 28206 11396
rect 31154 11340 31164 11396
rect 31220 11340 33404 11396
rect 33460 11340 33470 11396
rect 34850 11340 34860 11396
rect 34916 11340 38780 11396
rect 38836 11340 38846 11396
rect 45938 11340 45948 11396
rect 46004 11340 48188 11396
rect 48244 11340 48254 11396
rect 49746 11340 49756 11396
rect 49812 11340 50540 11396
rect 50596 11340 50606 11396
rect 2492 11284 2548 11340
rect 2492 11228 3612 11284
rect 3668 11228 3678 11284
rect 4498 11228 4508 11284
rect 4564 11228 5740 11284
rect 5796 11228 6748 11284
rect 6804 11228 7868 11284
rect 7924 11228 7934 11284
rect 14140 11172 14196 11340
rect 26908 11284 26964 11340
rect 22194 11228 22204 11284
rect 22260 11228 22876 11284
rect 22932 11228 22942 11284
rect 25666 11228 25676 11284
rect 25732 11228 28476 11284
rect 28532 11228 28542 11284
rect 29698 11228 29708 11284
rect 29764 11228 30716 11284
rect 30772 11228 32060 11284
rect 32116 11228 32126 11284
rect 32844 11172 32900 11340
rect 35746 11228 35756 11284
rect 35812 11228 37324 11284
rect 37380 11228 37390 11284
rect 43250 11228 43260 11284
rect 43316 11228 43932 11284
rect 43988 11228 45164 11284
rect 45220 11228 45230 11284
rect 45714 11228 45724 11284
rect 45780 11228 46396 11284
rect 46452 11228 46462 11284
rect 3266 11116 3276 11172
rect 3332 11116 3948 11172
rect 4004 11116 4014 11172
rect 5842 11116 5852 11172
rect 5908 11116 6412 11172
rect 6468 11116 6478 11172
rect 14140 11116 18284 11172
rect 18340 11116 18350 11172
rect 18722 11116 18732 11172
rect 18788 11116 19292 11172
rect 19348 11116 26908 11172
rect 27346 11116 27356 11172
rect 27412 11116 28364 11172
rect 28420 11116 28430 11172
rect 29474 11116 29484 11172
rect 29540 11116 30940 11172
rect 30996 11116 31006 11172
rect 32834 11116 32844 11172
rect 32900 11116 32910 11172
rect 34262 11116 34300 11172
rect 34356 11116 34366 11172
rect 35270 11116 35308 11172
rect 35364 11116 35374 11172
rect 26852 11060 26908 11116
rect 5394 11004 5404 11060
rect 5460 11004 7756 11060
rect 7812 11004 8316 11060
rect 8372 11004 8382 11060
rect 26852 11004 29204 11060
rect 30370 11004 30380 11060
rect 30436 11004 31724 11060
rect 31780 11004 31790 11060
rect 32610 11004 32620 11060
rect 32676 11004 34524 11060
rect 34580 11004 34590 11060
rect 35410 11004 35420 11060
rect 35476 11004 35756 11060
rect 35812 11004 35822 11060
rect 38612 11004 43988 11060
rect 15508 10948 15518 11004
rect 15574 10948 15622 11004
rect 15678 10948 15726 11004
rect 15782 10948 15792 11004
rect 22978 10892 22988 10948
rect 23044 10892 23324 10948
rect 23380 10892 23390 10948
rect 26338 10892 26348 10948
rect 26404 10892 27244 10948
rect 27300 10892 27310 10948
rect 1026 10780 1036 10836
rect 1092 10780 2044 10836
rect 2100 10780 2110 10836
rect 7858 10780 7868 10836
rect 7924 10780 8204 10836
rect 8260 10780 15932 10836
rect 15988 10780 15998 10836
rect 16370 10780 16380 10836
rect 16436 10780 20636 10836
rect 20692 10780 20702 10836
rect 23426 10780 23436 10836
rect 23492 10780 25340 10836
rect 25396 10780 26124 10836
rect 26180 10780 27132 10836
rect 27188 10780 27198 10836
rect 29148 10724 29204 11004
rect 29815 10948 29825 11004
rect 29881 10948 29929 11004
rect 29985 10948 30033 11004
rect 30089 10948 30099 11004
rect 38612 10948 38668 11004
rect 30258 10892 30268 10948
rect 30324 10892 38668 10948
rect 43932 10836 43988 11004
rect 44122 10948 44132 11004
rect 44188 10948 44236 11004
rect 44292 10948 44340 11004
rect 44396 10948 44406 11004
rect 58429 10948 58439 11004
rect 58495 10948 58543 11004
rect 58599 10948 58647 11004
rect 58703 10948 58713 11004
rect 29362 10780 29372 10836
rect 29428 10780 31276 10836
rect 31332 10780 32172 10836
rect 32228 10780 32238 10836
rect 32508 10780 39564 10836
rect 39620 10780 41804 10836
rect 41860 10780 41870 10836
rect 43932 10780 53900 10836
rect 53956 10780 53966 10836
rect 1698 10668 1708 10724
rect 1764 10668 3388 10724
rect 3444 10668 3454 10724
rect 7634 10668 7644 10724
rect 7700 10668 8316 10724
rect 8372 10668 19740 10724
rect 19796 10668 19806 10724
rect 22754 10668 22764 10724
rect 22820 10668 23100 10724
rect 23156 10668 23166 10724
rect 27010 10668 27020 10724
rect 27076 10668 27356 10724
rect 27412 10668 27422 10724
rect 29148 10668 31500 10724
rect 31556 10668 31566 10724
rect 32508 10612 32564 10780
rect 33954 10668 33964 10724
rect 34020 10668 36316 10724
rect 36372 10668 37212 10724
rect 37268 10668 38556 10724
rect 38612 10668 38622 10724
rect 39330 10668 39340 10724
rect 39396 10668 41692 10724
rect 41748 10668 41758 10724
rect 8642 10556 8652 10612
rect 8708 10556 8718 10612
rect 8978 10556 8988 10612
rect 9044 10556 13580 10612
rect 13636 10556 13646 10612
rect 19282 10556 19292 10612
rect 19348 10556 23772 10612
rect 23828 10556 23838 10612
rect 28130 10556 28140 10612
rect 28196 10556 29708 10612
rect 29764 10556 29774 10612
rect 29932 10556 32564 10612
rect 33394 10556 33404 10612
rect 33460 10556 34300 10612
rect 34356 10556 34524 10612
rect 34580 10556 34590 10612
rect 38882 10556 38892 10612
rect 38948 10556 40908 10612
rect 40964 10556 40974 10612
rect 43586 10556 43596 10612
rect 43652 10556 44716 10612
rect 44772 10556 44782 10612
rect 8652 10500 8708 10556
rect 29932 10500 29988 10556
rect 8652 10444 9996 10500
rect 10052 10444 10668 10500
rect 10724 10444 11004 10500
rect 11060 10444 11070 10500
rect 15250 10444 15260 10500
rect 15316 10444 19180 10500
rect 19236 10444 21980 10500
rect 22036 10444 22316 10500
rect 22372 10444 22382 10500
rect 22866 10444 22876 10500
rect 22932 10444 29988 10500
rect 33730 10444 33740 10500
rect 33796 10444 34636 10500
rect 34692 10444 35756 10500
rect 35812 10444 35822 10500
rect 41122 10444 41132 10500
rect 41188 10444 41244 10500
rect 41300 10444 41310 10500
rect 41458 10444 41468 10500
rect 41524 10444 41562 10500
rect 0 10304 800 10416
rect 14466 10332 14476 10388
rect 14532 10332 19628 10388
rect 19684 10332 22988 10388
rect 23044 10332 23054 10388
rect 23202 10332 23212 10388
rect 23268 10332 30268 10388
rect 30324 10332 30334 10388
rect 34066 10332 34076 10388
rect 34132 10332 35084 10388
rect 35140 10332 35868 10388
rect 35924 10332 35934 10388
rect 36092 10332 42252 10388
rect 42308 10332 42318 10388
rect 36092 10276 36148 10332
rect 2146 10220 2156 10276
rect 2212 10220 5852 10276
rect 5908 10220 5918 10276
rect 12796 10220 16380 10276
rect 16436 10220 16446 10276
rect 16818 10220 16828 10276
rect 16884 10220 17388 10276
rect 17444 10220 17454 10276
rect 17826 10220 17836 10276
rect 17892 10220 20748 10276
rect 20804 10220 21644 10276
rect 21700 10220 21710 10276
rect 28466 10220 28476 10276
rect 28532 10220 29820 10276
rect 29876 10220 29886 10276
rect 32050 10220 32060 10276
rect 32116 10220 33180 10276
rect 33236 10220 33246 10276
rect 33506 10220 33516 10276
rect 33572 10220 36148 10276
rect 42802 10220 42812 10276
rect 42868 10220 43036 10276
rect 43092 10220 43102 10276
rect 8355 10164 8365 10220
rect 8421 10164 8469 10220
rect 8525 10164 8573 10220
rect 8629 10164 8639 10220
rect 12796 10164 12852 10220
rect 22662 10164 22672 10220
rect 22728 10164 22776 10220
rect 22832 10164 22880 10220
rect 22936 10164 22946 10220
rect 36969 10164 36979 10220
rect 37035 10164 37083 10220
rect 37139 10164 37187 10220
rect 37243 10164 37253 10220
rect 51276 10164 51286 10220
rect 51342 10164 51390 10220
rect 51446 10164 51494 10220
rect 51550 10164 51560 10220
rect 2482 10108 2492 10164
rect 2548 10108 2558 10164
rect 12562 10108 12572 10164
rect 12628 10108 12852 10164
rect 14354 10108 14364 10164
rect 14420 10108 18172 10164
rect 18228 10108 18238 10164
rect 20514 10108 20524 10164
rect 20580 10108 22596 10164
rect 2492 10052 2548 10108
rect 22540 10052 22596 10108
rect 23100 10108 27356 10164
rect 27412 10108 27422 10164
rect 28354 10108 28364 10164
rect 28420 10108 28644 10164
rect 31154 10108 31164 10164
rect 31220 10108 35420 10164
rect 35476 10108 35486 10164
rect 38658 10108 38668 10164
rect 38724 10108 44716 10164
rect 44772 10108 45332 10164
rect 53890 10108 53900 10164
rect 53956 10108 54908 10164
rect 54964 10108 54974 10164
rect 23100 10052 23156 10108
rect 1810 9996 1820 10052
rect 1876 9996 3052 10052
rect 3108 9996 3118 10052
rect 8754 9996 8764 10052
rect 8820 9996 11004 10052
rect 11060 9996 11070 10052
rect 22540 9996 23156 10052
rect 23650 9996 23660 10052
rect 23716 9996 25228 10052
rect 25284 9996 26124 10052
rect 26180 9996 26908 10052
rect 4274 9884 4284 9940
rect 4340 9884 9772 9940
rect 9828 9884 9838 9940
rect 10434 9884 10444 9940
rect 10500 9884 12796 9940
rect 12852 9884 13916 9940
rect 13972 9884 13982 9940
rect 24322 9884 24332 9940
rect 24388 9884 26012 9940
rect 26068 9884 26078 9940
rect 9772 9828 9828 9884
rect 26852 9828 26908 9996
rect 28588 9940 28644 10108
rect 34290 9996 34300 10052
rect 34356 9996 34860 10052
rect 34916 9996 34926 10052
rect 35298 9996 35308 10052
rect 35364 9996 35756 10052
rect 35812 9996 35822 10052
rect 39442 9996 39452 10052
rect 39508 9996 42812 10052
rect 42868 9996 43036 10052
rect 43092 9996 43102 10052
rect 44258 9996 44268 10052
rect 44324 9996 45052 10052
rect 45108 9996 45118 10052
rect 28588 9884 31724 9940
rect 31780 9884 32508 9940
rect 32564 9884 42140 9940
rect 42196 9884 42206 9940
rect 42700 9884 43596 9940
rect 43652 9884 43662 9940
rect 42700 9828 42756 9884
rect 44268 9828 44324 9996
rect 45276 9828 45332 10108
rect 45910 9996 45948 10052
rect 46004 9996 46014 10052
rect 46610 9996 46620 10052
rect 46676 9996 46956 10052
rect 47012 9996 47022 10052
rect 50642 9996 50652 10052
rect 50708 9996 55916 10052
rect 55972 9996 56700 10052
rect 56756 9996 56766 10052
rect 9772 9772 10220 9828
rect 10276 9772 10668 9828
rect 10724 9772 10734 9828
rect 16370 9772 16380 9828
rect 16436 9772 22988 9828
rect 23044 9772 23660 9828
rect 23716 9772 23726 9828
rect 26852 9772 27020 9828
rect 27076 9772 27086 9828
rect 33618 9772 33628 9828
rect 33684 9772 35308 9828
rect 35364 9772 35374 9828
rect 41794 9772 41804 9828
rect 41860 9772 42756 9828
rect 43474 9772 43484 9828
rect 43540 9772 43932 9828
rect 43988 9772 44324 9828
rect 45266 9772 45276 9828
rect 45332 9772 45342 9828
rect 45938 9772 45948 9828
rect 46004 9772 46620 9828
rect 46676 9772 46686 9828
rect 48514 9772 48524 9828
rect 48580 9772 49756 9828
rect 49812 9772 49822 9828
rect 51650 9772 51660 9828
rect 51716 9772 53116 9828
rect 53172 9772 53182 9828
rect 54450 9772 54460 9828
rect 54516 9772 55132 9828
rect 55188 9772 55198 9828
rect 2370 9660 2380 9716
rect 2436 9660 2940 9716
rect 2996 9660 3006 9716
rect 4610 9660 4620 9716
rect 4676 9660 5292 9716
rect 5348 9660 9436 9716
rect 9492 9660 9502 9716
rect 10546 9660 10556 9716
rect 10612 9660 11060 9716
rect 15026 9660 15036 9716
rect 15092 9660 21532 9716
rect 21588 9660 22876 9716
rect 22932 9660 22942 9716
rect 26450 9660 26460 9716
rect 26516 9660 31388 9716
rect 31444 9660 31454 9716
rect 39890 9660 39900 9716
rect 39956 9660 40684 9716
rect 40740 9660 40750 9716
rect 41682 9660 41692 9716
rect 41748 9660 43708 9716
rect 43764 9660 43774 9716
rect 45378 9660 45388 9716
rect 45444 9660 45612 9716
rect 45668 9660 45678 9716
rect 47394 9660 47404 9716
rect 47460 9660 48972 9716
rect 49028 9660 49038 9716
rect 51874 9660 51884 9716
rect 51940 9660 52556 9716
rect 52612 9660 52622 9716
rect 11004 9604 11060 9660
rect 5170 9548 5180 9604
rect 5236 9548 6188 9604
rect 6244 9548 9548 9604
rect 9604 9548 9614 9604
rect 9762 9548 9772 9604
rect 9828 9548 10668 9604
rect 10724 9548 10734 9604
rect 10994 9548 11004 9604
rect 11060 9548 11070 9604
rect 12002 9548 12012 9604
rect 12068 9548 14252 9604
rect 14308 9548 14318 9604
rect 19730 9548 19740 9604
rect 19796 9548 20188 9604
rect 20244 9548 20254 9604
rect 23314 9548 23324 9604
rect 23380 9548 26852 9604
rect 26908 9548 26918 9604
rect 27010 9548 27020 9604
rect 27076 9548 27916 9604
rect 27972 9548 29372 9604
rect 29428 9548 29438 9604
rect 30930 9548 30940 9604
rect 30996 9548 39676 9604
rect 39732 9548 39742 9604
rect 41458 9548 41468 9604
rect 41524 9548 42476 9604
rect 42532 9548 42542 9604
rect 42690 9548 42700 9604
rect 42756 9548 43148 9604
rect 43204 9548 43214 9604
rect 46946 9548 46956 9604
rect 47012 9548 48188 9604
rect 48244 9548 48254 9604
rect 17154 9436 17164 9492
rect 17220 9436 22260 9492
rect 25890 9436 25900 9492
rect 25956 9436 27804 9492
rect 27860 9436 27870 9492
rect 31042 9436 31052 9492
rect 31108 9436 33180 9492
rect 33236 9436 33516 9492
rect 33572 9436 33582 9492
rect 42242 9436 42252 9492
rect 42308 9436 43932 9492
rect 43988 9436 43998 9492
rect 15508 9380 15518 9436
rect 15574 9380 15622 9436
rect 15678 9380 15726 9436
rect 15782 9380 15792 9436
rect 22204 9380 22260 9436
rect 29815 9380 29825 9436
rect 29881 9380 29929 9436
rect 29985 9380 30033 9436
rect 30089 9380 30099 9436
rect 44122 9380 44132 9436
rect 44188 9380 44236 9436
rect 44292 9380 44340 9436
rect 44396 9380 44406 9436
rect 58429 9380 58439 9436
rect 58495 9380 58543 9436
rect 58599 9380 58647 9436
rect 58703 9380 58713 9436
rect 2706 9324 2716 9380
rect 2772 9324 4844 9380
rect 4900 9324 4910 9380
rect 6738 9324 6748 9380
rect 6804 9324 8204 9380
rect 8260 9324 9660 9380
rect 9716 9324 9726 9380
rect 19058 9324 19068 9380
rect 19124 9324 20860 9380
rect 20916 9324 20926 9380
rect 22204 9324 26908 9380
rect 26964 9324 28868 9380
rect 0 9184 800 9296
rect 28812 9268 28868 9324
rect 30268 9324 38332 9380
rect 38388 9324 39004 9380
rect 39060 9324 39070 9380
rect 40338 9324 40348 9380
rect 40404 9324 43988 9380
rect 50194 9324 50204 9380
rect 50260 9324 50988 9380
rect 51044 9324 52332 9380
rect 52388 9324 52398 9380
rect 2146 9212 2156 9268
rect 2212 9212 5068 9268
rect 5124 9212 5134 9268
rect 6290 9212 6300 9268
rect 6356 9212 6972 9268
rect 7028 9212 7038 9268
rect 10210 9212 10220 9268
rect 10276 9212 10286 9268
rect 19618 9212 19628 9268
rect 19684 9212 27132 9268
rect 27188 9212 28028 9268
rect 28084 9212 28094 9268
rect 28802 9212 28812 9268
rect 28868 9212 30044 9268
rect 30100 9212 30110 9268
rect 1810 9100 1820 9156
rect 1876 9100 2716 9156
rect 2772 9100 2782 9156
rect 3042 9100 3052 9156
rect 3108 9100 8988 9156
rect 9044 9100 9054 9156
rect 4610 8988 4620 9044
rect 4676 8988 5404 9044
rect 5460 8988 5470 9044
rect 5842 8988 5852 9044
rect 5908 8988 7644 9044
rect 7700 8988 7710 9044
rect 9650 8876 9660 8932
rect 9716 8876 9996 8932
rect 10052 8876 10062 8932
rect 10220 8820 10276 9212
rect 30268 9156 30324 9324
rect 31714 9212 31724 9268
rect 31780 9212 32844 9268
rect 32900 9212 32910 9268
rect 35186 9212 35196 9268
rect 35252 9212 40908 9268
rect 40964 9212 42028 9268
rect 42084 9212 42094 9268
rect 16818 9100 16828 9156
rect 16884 9100 18060 9156
rect 18116 9100 18126 9156
rect 20402 9100 20412 9156
rect 20468 9100 23100 9156
rect 23156 9100 23166 9156
rect 24546 9100 24556 9156
rect 24612 9100 26684 9156
rect 26740 9100 26750 9156
rect 27794 9100 27804 9156
rect 27860 9100 29932 9156
rect 29988 9100 30324 9156
rect 32162 9100 32172 9156
rect 32228 9100 39452 9156
rect 39508 9100 39518 9156
rect 40002 9100 40012 9156
rect 40068 9100 42588 9156
rect 42644 9100 42654 9156
rect 43932 9044 43988 9324
rect 46022 9212 46060 9268
rect 46116 9212 46126 9268
rect 49746 9100 49756 9156
rect 49812 9100 50988 9156
rect 51044 9100 51054 9156
rect 52882 9100 52892 9156
rect 52948 9100 53788 9156
rect 53844 9100 53854 9156
rect 13122 8988 13132 9044
rect 13188 8988 13916 9044
rect 13972 8988 14700 9044
rect 14756 8988 14766 9044
rect 24098 8988 24108 9044
rect 24164 8988 26124 9044
rect 26180 8988 26190 9044
rect 26898 8988 26908 9044
rect 26964 8988 30492 9044
rect 30548 8988 35644 9044
rect 35700 8988 35710 9044
rect 41206 8988 41244 9044
rect 41300 8988 43036 9044
rect 43092 8988 43102 9044
rect 43922 8988 43932 9044
rect 43988 8988 43998 9044
rect 45490 8988 45500 9044
rect 45556 8988 47404 9044
rect 47460 8988 47470 9044
rect 53106 8988 53116 9044
rect 53172 8988 54012 9044
rect 54068 8988 54078 9044
rect 54898 8988 54908 9044
rect 54964 8988 54974 9044
rect 55682 8988 55692 9044
rect 55748 8988 56588 9044
rect 56644 8988 56654 9044
rect 54908 8932 54964 8988
rect 11218 8876 11228 8932
rect 11284 8876 15484 8932
rect 15540 8876 16044 8932
rect 16100 8876 16110 8932
rect 16258 8876 16268 8932
rect 16324 8876 17836 8932
rect 17892 8876 17902 8932
rect 23426 8876 23436 8932
rect 23492 8876 25900 8932
rect 25956 8876 25966 8932
rect 27570 8876 27580 8932
rect 27636 8876 29036 8932
rect 29092 8876 31500 8932
rect 31556 8876 31566 8932
rect 34598 8876 34636 8932
rect 34692 8876 34702 8932
rect 34850 8876 34860 8932
rect 34916 8876 40964 8932
rect 45378 8876 45388 8932
rect 45444 8876 48524 8932
rect 48580 8876 48590 8932
rect 54562 8876 54572 8932
rect 54628 8876 54964 8932
rect 40908 8820 40964 8876
rect 4946 8764 4956 8820
rect 5012 8764 8204 8820
rect 8260 8764 8270 8820
rect 8530 8764 8540 8820
rect 8596 8764 8820 8820
rect 10210 8764 10220 8820
rect 10276 8764 10286 8820
rect 13010 8764 13020 8820
rect 13076 8764 15148 8820
rect 15204 8764 15214 8820
rect 15372 8764 18172 8820
rect 18228 8764 18238 8820
rect 21634 8764 21644 8820
rect 21700 8764 23996 8820
rect 24052 8764 25788 8820
rect 25844 8764 25854 8820
rect 26786 8764 26796 8820
rect 26852 8764 35980 8820
rect 36036 8764 38668 8820
rect 38724 8764 38734 8820
rect 40908 8764 41804 8820
rect 41860 8764 41870 8820
rect 42998 8764 43036 8820
rect 43092 8764 43102 8820
rect 46274 8764 46284 8820
rect 46340 8764 47068 8820
rect 47124 8764 47134 8820
rect 49970 8764 49980 8820
rect 50036 8764 50316 8820
rect 50372 8764 50382 8820
rect 55906 8764 55916 8820
rect 55972 8764 57484 8820
rect 57540 8764 57550 8820
rect 8355 8596 8365 8652
rect 8421 8596 8469 8652
rect 8525 8596 8573 8652
rect 8629 8596 8639 8652
rect 8764 8372 8820 8764
rect 15372 8708 15428 8764
rect 14242 8652 14252 8708
rect 14308 8652 15428 8708
rect 15484 8652 18620 8708
rect 18676 8652 18686 8708
rect 25666 8652 25676 8708
rect 25732 8652 26348 8708
rect 26404 8652 26414 8708
rect 27794 8652 27804 8708
rect 27860 8652 28252 8708
rect 28308 8652 28318 8708
rect 40226 8652 40236 8708
rect 40292 8652 40796 8708
rect 40852 8652 40862 8708
rect 43250 8652 43260 8708
rect 43316 8652 45388 8708
rect 45444 8652 45454 8708
rect 15484 8596 15540 8652
rect 22662 8596 22672 8652
rect 22728 8596 22776 8652
rect 22832 8596 22880 8652
rect 22936 8596 22946 8652
rect 36969 8596 36979 8652
rect 37035 8596 37083 8652
rect 37139 8596 37187 8652
rect 37243 8596 37253 8652
rect 51276 8596 51286 8652
rect 51342 8596 51390 8652
rect 51446 8596 51494 8652
rect 51550 8596 51560 8652
rect 13794 8540 13804 8596
rect 13860 8540 15540 8596
rect 26852 8540 27692 8596
rect 27748 8540 28476 8596
rect 28532 8540 30268 8596
rect 30324 8540 30334 8596
rect 30706 8540 30716 8596
rect 30772 8540 31276 8596
rect 31332 8540 33740 8596
rect 33796 8540 33806 8596
rect 52098 8540 52108 8596
rect 52164 8540 52892 8596
rect 52948 8540 52958 8596
rect 12450 8428 12460 8484
rect 12516 8428 15148 8484
rect 15092 8372 15148 8428
rect 15260 8428 17500 8484
rect 17556 8428 19740 8484
rect 19796 8428 20412 8484
rect 20468 8428 20478 8484
rect 23314 8428 23324 8484
rect 23380 8428 24108 8484
rect 24164 8428 24174 8484
rect 15260 8372 15316 8428
rect 26852 8372 26908 8540
rect 27794 8428 27804 8484
rect 27860 8428 28140 8484
rect 28196 8428 31052 8484
rect 31108 8428 31118 8484
rect 38770 8428 38780 8484
rect 38836 8428 39900 8484
rect 39956 8428 39966 8484
rect 44034 8428 44044 8484
rect 44100 8428 44604 8484
rect 44660 8428 55356 8484
rect 55412 8428 55422 8484
rect 8764 8316 13356 8372
rect 13412 8316 13692 8372
rect 13748 8316 14924 8372
rect 14980 8316 14990 8372
rect 15092 8316 15316 8372
rect 16818 8316 16828 8372
rect 16884 8316 17724 8372
rect 17780 8316 18396 8372
rect 18452 8316 18462 8372
rect 18620 8316 23100 8372
rect 23156 8316 25228 8372
rect 25284 8316 25294 8372
rect 25554 8316 25564 8372
rect 25620 8316 26908 8372
rect 33394 8316 33404 8372
rect 33460 8316 34300 8372
rect 34356 8316 34366 8372
rect 34738 8316 34748 8372
rect 34804 8316 35420 8372
rect 35476 8316 35486 8372
rect 35970 8316 35980 8372
rect 36036 8316 37772 8372
rect 37828 8316 38892 8372
rect 38948 8316 38958 8372
rect 45602 8316 45612 8372
rect 45668 8316 46396 8372
rect 46452 8316 47292 8372
rect 47348 8316 47358 8372
rect 52994 8316 53004 8372
rect 53060 8316 54348 8372
rect 54404 8316 54414 8372
rect 54674 8316 54684 8372
rect 54740 8316 55468 8372
rect 55524 8316 55534 8372
rect 56242 8316 56252 8372
rect 56308 8316 56924 8372
rect 56980 8316 56990 8372
rect 18620 8260 18676 8316
rect 11890 8204 11900 8260
rect 11956 8204 13580 8260
rect 13636 8204 15708 8260
rect 15764 8204 17164 8260
rect 17220 8204 17230 8260
rect 17490 8204 17500 8260
rect 17556 8204 18676 8260
rect 22754 8204 22764 8260
rect 22820 8204 25900 8260
rect 25956 8204 25966 8260
rect 27234 8204 27244 8260
rect 27300 8204 29596 8260
rect 29652 8204 29662 8260
rect 30370 8204 30380 8260
rect 30436 8204 33180 8260
rect 33236 8204 33246 8260
rect 33842 8204 33852 8260
rect 33908 8204 36092 8260
rect 36148 8204 37212 8260
rect 37268 8204 37278 8260
rect 46050 8204 46060 8260
rect 46116 8204 47068 8260
rect 47124 8204 47572 8260
rect 51426 8204 51436 8260
rect 51492 8204 54572 8260
rect 54628 8204 54638 8260
rect 55794 8204 55804 8260
rect 55860 8204 56476 8260
rect 56532 8204 57260 8260
rect 57316 8204 57326 8260
rect 0 8064 800 8176
rect 47516 8148 47572 8204
rect 12674 8092 12684 8148
rect 12740 8092 15260 8148
rect 15316 8092 15326 8148
rect 15586 8092 15596 8148
rect 15652 8092 15662 8148
rect 15922 8092 15932 8148
rect 15988 8092 19292 8148
rect 19348 8092 19358 8148
rect 23090 8092 23100 8148
rect 23156 8092 23772 8148
rect 23828 8092 23838 8148
rect 26114 8092 26124 8148
rect 26180 8092 32060 8148
rect 32116 8092 32732 8148
rect 32788 8092 34188 8148
rect 34244 8092 34254 8148
rect 36866 8092 36876 8148
rect 36932 8092 38556 8148
rect 38612 8092 38622 8148
rect 43922 8092 43932 8148
rect 43988 8092 46172 8148
rect 46228 8092 46238 8148
rect 47506 8092 47516 8148
rect 47572 8092 47582 8148
rect 48066 8092 48076 8148
rect 48132 8092 48748 8148
rect 48804 8092 48814 8148
rect 15596 8036 15652 8092
rect 2818 7980 2828 8036
rect 2884 7980 5740 8036
rect 5796 7980 5806 8036
rect 8754 7980 8764 8036
rect 8820 7980 10780 8036
rect 10836 7980 10846 8036
rect 12786 7980 12796 8036
rect 12852 7980 14028 8036
rect 14084 7980 14094 8036
rect 14466 7980 14476 8036
rect 14532 7980 15652 8036
rect 21746 7980 21756 8036
rect 21812 7980 21822 8036
rect 27122 7980 27132 8036
rect 27188 7980 30940 8036
rect 30996 7980 31612 8036
rect 31668 7980 31678 8036
rect 33618 7980 33628 8036
rect 33684 7980 35868 8036
rect 35924 7980 35934 8036
rect 41570 7980 41580 8036
rect 41636 7980 42364 8036
rect 42420 7980 42430 8036
rect 43698 7980 43708 8036
rect 43764 7980 44716 8036
rect 44772 7980 44782 8036
rect 44930 7980 44940 8036
rect 44996 7980 46620 8036
rect 46676 7980 46686 8036
rect 53330 7980 53340 8036
rect 53396 7980 54908 8036
rect 54964 7980 54974 8036
rect 21756 7924 21812 7980
rect 2258 7868 2268 7924
rect 2324 7868 3276 7924
rect 3332 7868 3836 7924
rect 3892 7868 3902 7924
rect 13346 7868 13356 7924
rect 13412 7868 14364 7924
rect 14420 7868 14430 7924
rect 15932 7868 20860 7924
rect 20916 7868 20926 7924
rect 21756 7868 27692 7924
rect 27748 7868 27758 7924
rect 38658 7868 38668 7924
rect 38724 7868 40236 7924
rect 40292 7868 40302 7924
rect 44818 7868 44828 7924
rect 44884 7868 46060 7924
rect 46116 7868 48748 7924
rect 48804 7868 48814 7924
rect 15508 7812 15518 7868
rect 15574 7812 15622 7868
rect 15678 7812 15726 7868
rect 15782 7812 15792 7868
rect 15932 7700 15988 7868
rect 29815 7812 29825 7868
rect 29881 7812 29929 7868
rect 29985 7812 30033 7868
rect 30089 7812 30099 7868
rect 44122 7812 44132 7868
rect 44188 7812 44236 7868
rect 44292 7812 44340 7868
rect 44396 7812 44406 7868
rect 58429 7812 58439 7868
rect 58495 7812 58543 7868
rect 58599 7812 58647 7868
rect 58703 7812 58713 7868
rect 17826 7756 17836 7812
rect 17892 7756 26572 7812
rect 26628 7756 26908 7812
rect 34486 7756 34524 7812
rect 34580 7756 34590 7812
rect 36418 7756 36428 7812
rect 36484 7756 37772 7812
rect 37828 7756 37838 7812
rect 26852 7700 26908 7756
rect 2258 7644 2268 7700
rect 2324 7644 3500 7700
rect 3556 7644 3566 7700
rect 5618 7644 5628 7700
rect 5684 7644 6636 7700
rect 6692 7644 7196 7700
rect 7252 7644 7262 7700
rect 15026 7644 15036 7700
rect 15092 7644 15988 7700
rect 16482 7644 16492 7700
rect 16548 7644 20188 7700
rect 20244 7644 20254 7700
rect 20850 7644 20860 7700
rect 20916 7644 23100 7700
rect 23156 7644 23166 7700
rect 26852 7644 27020 7700
rect 27076 7644 27086 7700
rect 28018 7644 28028 7700
rect 28084 7644 28700 7700
rect 28756 7644 28766 7700
rect 30156 7644 33516 7700
rect 33572 7644 33582 7700
rect 35410 7644 35420 7700
rect 35476 7644 39452 7700
rect 39508 7644 39518 7700
rect 42578 7644 42588 7700
rect 42644 7644 44828 7700
rect 44884 7644 44894 7700
rect 50372 7644 52444 7700
rect 52500 7644 52510 7700
rect 55010 7644 55020 7700
rect 55076 7644 57148 7700
rect 57204 7644 57214 7700
rect 30156 7588 30212 7644
rect 33516 7588 33572 7644
rect 14018 7532 14028 7588
rect 14084 7532 15372 7588
rect 15428 7532 15438 7588
rect 15922 7532 15932 7588
rect 15988 7532 15998 7588
rect 19170 7532 19180 7588
rect 19236 7532 21700 7588
rect 23874 7532 23884 7588
rect 23940 7532 30212 7588
rect 30370 7532 30380 7588
rect 30436 7532 30940 7588
rect 30996 7532 31006 7588
rect 33516 7532 36876 7588
rect 36932 7532 36942 7588
rect 46946 7532 46956 7588
rect 47012 7532 47628 7588
rect 47684 7532 47694 7588
rect 49522 7532 49532 7588
rect 49588 7532 50316 7588
rect 50372 7532 50428 7644
rect 51762 7532 51772 7588
rect 51828 7532 54124 7588
rect 54180 7532 54190 7588
rect 5954 7420 5964 7476
rect 6020 7420 7196 7476
rect 7252 7420 7262 7476
rect 15932 7364 15988 7532
rect 21644 7476 21700 7532
rect 18834 7420 18844 7476
rect 18900 7420 20076 7476
rect 20132 7420 20142 7476
rect 21634 7420 21644 7476
rect 21700 7420 22988 7476
rect 23044 7420 23054 7476
rect 31378 7420 31388 7476
rect 31444 7420 32284 7476
rect 32340 7420 33740 7476
rect 33796 7420 33806 7476
rect 38210 7420 38220 7476
rect 38276 7420 40908 7476
rect 40964 7420 40974 7476
rect 43474 7420 43484 7476
rect 43540 7420 44604 7476
rect 44660 7420 44670 7476
rect 45714 7420 45724 7476
rect 45780 7420 46396 7476
rect 46452 7420 48076 7476
rect 48132 7420 48142 7476
rect 49186 7420 49196 7476
rect 49252 7420 50540 7476
rect 50596 7420 50606 7476
rect 4722 7308 4732 7364
rect 4788 7308 5516 7364
rect 5572 7308 5582 7364
rect 6738 7308 6748 7364
rect 6804 7308 7308 7364
rect 7364 7308 7374 7364
rect 8642 7308 8652 7364
rect 8708 7308 15988 7364
rect 19842 7308 19852 7364
rect 19908 7308 20860 7364
rect 20916 7308 20926 7364
rect 29586 7308 29596 7364
rect 29652 7308 31052 7364
rect 31108 7308 31118 7364
rect 33842 7308 33852 7364
rect 33908 7308 38668 7364
rect 43362 7308 43372 7364
rect 43428 7308 46508 7364
rect 46564 7308 46574 7364
rect 46722 7308 46732 7364
rect 46788 7308 51548 7364
rect 51604 7308 55244 7364
rect 55300 7308 57036 7364
rect 57092 7308 57102 7364
rect 5394 7196 5404 7252
rect 5460 7196 6860 7252
rect 6916 7196 7756 7252
rect 7812 7196 7822 7252
rect 8306 7196 8316 7252
rect 8372 7196 15148 7252
rect 15698 7196 15708 7252
rect 15764 7196 18732 7252
rect 18788 7196 18798 7252
rect 20178 7196 20188 7252
rect 20244 7196 25564 7252
rect 25620 7196 26236 7252
rect 26292 7196 26302 7252
rect 32722 7196 32732 7252
rect 32788 7196 37436 7252
rect 37492 7196 37502 7252
rect 0 6944 800 7056
rect 8355 7028 8365 7084
rect 8421 7028 8469 7084
rect 8525 7028 8573 7084
rect 8629 7028 8639 7084
rect 15092 6916 15148 7196
rect 38612 7140 38668 7308
rect 46508 7252 46564 7308
rect 46508 7196 48188 7252
rect 48244 7196 48254 7252
rect 50372 7196 51828 7252
rect 50372 7140 50428 7196
rect 51772 7140 51828 7196
rect 15250 7084 15260 7140
rect 15316 7084 19964 7140
rect 20020 7084 20030 7140
rect 31602 7084 31612 7140
rect 31668 7084 33180 7140
rect 33236 7084 34972 7140
rect 35028 7084 35038 7140
rect 38612 7084 50428 7140
rect 51762 7084 51772 7140
rect 51828 7084 51838 7140
rect 22662 7028 22672 7084
rect 22728 7028 22776 7084
rect 22832 7028 22880 7084
rect 22936 7028 22946 7084
rect 36969 7028 36979 7084
rect 37035 7028 37083 7084
rect 37139 7028 37187 7084
rect 37243 7028 37253 7084
rect 51276 7028 51286 7084
rect 51342 7028 51390 7084
rect 51446 7028 51494 7084
rect 51550 7028 51560 7084
rect 15362 6972 15372 7028
rect 15428 6972 21308 7028
rect 21364 6972 21868 7028
rect 21924 6972 21934 7028
rect 26674 6972 26684 7028
rect 26740 6972 30044 7028
rect 30100 6972 30110 7028
rect 34290 6972 34300 7028
rect 34356 6972 34748 7028
rect 34804 6972 34814 7028
rect 44370 6972 44380 7028
rect 44436 6972 45724 7028
rect 45780 6972 46844 7028
rect 46900 6972 46910 7028
rect 51874 6972 51884 7028
rect 51940 6972 53452 7028
rect 53508 6972 53518 7028
rect 3602 6860 3612 6916
rect 3668 6860 13468 6916
rect 13524 6860 13534 6916
rect 15092 6860 17500 6916
rect 17556 6860 17566 6916
rect 21074 6860 21084 6916
rect 21140 6860 22764 6916
rect 22820 6860 22830 6916
rect 29138 6860 29148 6916
rect 29204 6860 38780 6916
rect 38836 6860 38846 6916
rect 42018 6860 42028 6916
rect 42084 6860 56812 6916
rect 56868 6860 56878 6916
rect 12786 6748 12796 6804
rect 12852 6748 14700 6804
rect 14756 6748 15148 6804
rect 15204 6748 15214 6804
rect 15474 6748 15484 6804
rect 15540 6748 16828 6804
rect 16884 6748 16894 6804
rect 32610 6748 32620 6804
rect 32676 6748 35084 6804
rect 35140 6748 35980 6804
rect 36036 6748 36540 6804
rect 36596 6748 36606 6804
rect 42466 6748 42476 6804
rect 42532 6748 44156 6804
rect 44212 6748 44222 6804
rect 45910 6748 45948 6804
rect 46004 6748 46014 6804
rect 53218 6748 53228 6804
rect 53284 6748 54012 6804
rect 54068 6748 54078 6804
rect 4946 6636 4956 6692
rect 5012 6636 5740 6692
rect 5796 6636 5806 6692
rect 10770 6636 10780 6692
rect 10836 6636 12124 6692
rect 12180 6636 12190 6692
rect 16370 6636 16380 6692
rect 16436 6636 17836 6692
rect 17892 6636 17902 6692
rect 20514 6636 20524 6692
rect 20580 6636 25788 6692
rect 25844 6636 25854 6692
rect 27346 6636 27356 6692
rect 27412 6636 29820 6692
rect 29876 6636 32508 6692
rect 32564 6636 32956 6692
rect 33012 6636 33022 6692
rect 33282 6636 33292 6692
rect 33348 6636 33628 6692
rect 33684 6636 33694 6692
rect 34290 6636 34300 6692
rect 34356 6636 34860 6692
rect 34916 6636 35756 6692
rect 35812 6636 35822 6692
rect 42130 6636 42140 6692
rect 42196 6636 43260 6692
rect 43316 6636 44044 6692
rect 44100 6636 44110 6692
rect 46274 6636 46284 6692
rect 46340 6636 47740 6692
rect 47796 6636 47806 6692
rect 50418 6636 50428 6692
rect 50484 6636 53004 6692
rect 53060 6636 54124 6692
rect 54180 6636 54190 6692
rect 6178 6524 6188 6580
rect 6244 6524 8988 6580
rect 9044 6524 11228 6580
rect 11284 6524 11294 6580
rect 17490 6524 17500 6580
rect 17556 6524 23548 6580
rect 23604 6524 26124 6580
rect 26180 6524 26190 6580
rect 26852 6524 29148 6580
rect 29204 6524 29214 6580
rect 30818 6524 30828 6580
rect 30884 6524 31724 6580
rect 31780 6524 32844 6580
rect 32900 6524 32910 6580
rect 41682 6524 41692 6580
rect 41748 6524 42364 6580
rect 42420 6524 42430 6580
rect 48850 6524 48860 6580
rect 48916 6524 50316 6580
rect 50372 6524 50876 6580
rect 50932 6524 51324 6580
rect 51380 6524 51390 6580
rect 53442 6524 53452 6580
rect 53508 6524 53676 6580
rect 53732 6524 54796 6580
rect 54852 6524 54862 6580
rect 20626 6412 20636 6468
rect 20692 6412 22428 6468
rect 22484 6412 22494 6468
rect 26852 6356 26908 6524
rect 27570 6412 27580 6468
rect 27636 6412 29708 6468
rect 29764 6412 29774 6468
rect 31154 6412 31164 6468
rect 31220 6412 31444 6468
rect 38098 6412 38108 6468
rect 38164 6412 40796 6468
rect 40852 6412 40862 6468
rect 56130 6412 56140 6468
rect 56196 6412 57820 6468
rect 57876 6412 57886 6468
rect 31388 6356 31444 6412
rect 10770 6300 10780 6356
rect 10836 6300 14924 6356
rect 14980 6300 15148 6356
rect 16706 6300 16716 6356
rect 16772 6300 25228 6356
rect 25284 6300 25294 6356
rect 26674 6300 26684 6356
rect 26740 6300 26908 6356
rect 31378 6300 31388 6356
rect 31444 6300 31454 6356
rect 57026 6300 57036 6356
rect 57092 6300 58044 6356
rect 58100 6300 58110 6356
rect 15092 6132 15148 6300
rect 15508 6244 15518 6300
rect 15574 6244 15622 6300
rect 15678 6244 15726 6300
rect 15782 6244 15792 6300
rect 29815 6244 29825 6300
rect 29881 6244 29929 6300
rect 29985 6244 30033 6300
rect 30089 6244 30099 6300
rect 44122 6244 44132 6300
rect 44188 6244 44236 6300
rect 44292 6244 44340 6300
rect 44396 6244 44406 6300
rect 58429 6244 58439 6300
rect 58495 6244 58543 6300
rect 58599 6244 58647 6300
rect 58703 6244 58713 6300
rect 1922 6076 1932 6132
rect 1988 6076 3388 6132
rect 3938 6076 3948 6132
rect 4004 6076 5292 6132
rect 5348 6076 5964 6132
rect 6020 6076 6524 6132
rect 6580 6076 6590 6132
rect 7858 6076 7868 6132
rect 7924 6076 8988 6132
rect 9044 6076 9660 6132
rect 9716 6076 9726 6132
rect 11106 6076 11116 6132
rect 11172 6076 14476 6132
rect 14532 6076 14542 6132
rect 14802 6076 14812 6132
rect 14868 6076 14878 6132
rect 15092 6076 15820 6132
rect 15876 6076 15886 6132
rect 17042 6076 17052 6132
rect 17108 6076 20412 6132
rect 20468 6076 20478 6132
rect 22642 6076 22652 6132
rect 22708 6076 23436 6132
rect 23492 6076 23502 6132
rect 24658 6076 24668 6132
rect 24724 6076 26292 6132
rect 28690 6076 28700 6132
rect 28756 6076 29708 6132
rect 29764 6076 29774 6132
rect 34738 6076 34748 6132
rect 34804 6076 35644 6132
rect 35700 6076 41300 6132
rect 3332 6020 3388 6076
rect 3332 5964 6748 6020
rect 6804 5964 8652 6020
rect 8708 5964 8718 6020
rect 10434 5964 10444 6020
rect 10500 5964 11228 6020
rect 11284 5964 11294 6020
rect 11890 5964 11900 6020
rect 11956 5964 12124 6020
rect 12180 5964 12190 6020
rect 12338 5964 12348 6020
rect 12404 5964 12908 6020
rect 12964 5964 12974 6020
rect 0 5824 800 5936
rect 14812 5908 14868 6076
rect 26236 5908 26292 6076
rect 41244 6020 41300 6076
rect 26450 5964 26460 6020
rect 26516 5964 27804 6020
rect 27860 5964 30380 6020
rect 30436 5964 30446 6020
rect 30594 5964 30604 6020
rect 30660 5964 31836 6020
rect 31892 5964 31902 6020
rect 33954 5964 33964 6020
rect 34020 5964 34524 6020
rect 34580 5964 34590 6020
rect 37314 5964 37324 6020
rect 37380 5964 38668 6020
rect 38724 5964 38734 6020
rect 41234 5964 41244 6020
rect 41300 5964 41310 6020
rect 3602 5852 3612 5908
rect 3668 5852 6300 5908
rect 6356 5852 11116 5908
rect 11172 5852 11182 5908
rect 12562 5852 12572 5908
rect 12628 5852 13356 5908
rect 13412 5852 13422 5908
rect 14812 5852 16212 5908
rect 16706 5852 16716 5908
rect 16772 5852 24780 5908
rect 24836 5852 26012 5908
rect 26068 5852 26078 5908
rect 26236 5852 27468 5908
rect 27524 5852 27534 5908
rect 28914 5852 28924 5908
rect 28980 5852 32956 5908
rect 33012 5852 33022 5908
rect 33842 5852 33852 5908
rect 33908 5852 34300 5908
rect 34356 5852 34366 5908
rect 40226 5852 40236 5908
rect 40292 5852 42476 5908
rect 42532 5852 42542 5908
rect 47170 5852 47180 5908
rect 47236 5852 47628 5908
rect 47684 5852 50428 5908
rect 50484 5852 50494 5908
rect 56018 5852 56028 5908
rect 56084 5852 56588 5908
rect 56644 5852 58156 5908
rect 58212 5852 58222 5908
rect 16156 5796 16212 5852
rect 13122 5740 13132 5796
rect 13188 5740 14028 5796
rect 14084 5740 14094 5796
rect 16146 5740 16156 5796
rect 16212 5740 18284 5796
rect 18340 5740 18350 5796
rect 31042 5740 31052 5796
rect 31108 5740 38556 5796
rect 38612 5740 38622 5796
rect 39106 5740 39116 5796
rect 39172 5740 41020 5796
rect 41076 5740 41692 5796
rect 41748 5740 41758 5796
rect 47842 5740 47852 5796
rect 47908 5740 49756 5796
rect 49812 5740 49822 5796
rect 15922 5628 15932 5684
rect 15988 5628 26236 5684
rect 26292 5628 26302 5684
rect 26852 5628 34076 5684
rect 34132 5628 34300 5684
rect 34356 5628 35196 5684
rect 35252 5628 35262 5684
rect 38322 5628 38332 5684
rect 38388 5628 39676 5684
rect 39732 5628 39742 5684
rect 48178 5628 48188 5684
rect 48244 5628 48972 5684
rect 49028 5628 49038 5684
rect 26852 5572 26908 5628
rect 8866 5516 8876 5572
rect 8932 5516 14700 5572
rect 14756 5516 14766 5572
rect 23314 5516 23324 5572
rect 23380 5516 26908 5572
rect 27458 5516 27468 5572
rect 27524 5516 29708 5572
rect 29764 5516 29774 5572
rect 8355 5460 8365 5516
rect 8421 5460 8469 5516
rect 8525 5460 8573 5516
rect 8629 5460 8639 5516
rect 22662 5460 22672 5516
rect 22728 5460 22776 5516
rect 22832 5460 22880 5516
rect 22936 5460 22946 5516
rect 36969 5460 36979 5516
rect 37035 5460 37083 5516
rect 37139 5460 37187 5516
rect 37243 5460 37253 5516
rect 51276 5460 51286 5516
rect 51342 5460 51390 5516
rect 51446 5460 51494 5516
rect 51550 5460 51560 5516
rect 13122 5404 13132 5460
rect 13188 5404 21140 5460
rect 25218 5404 25228 5460
rect 25284 5404 25788 5460
rect 25844 5404 29260 5460
rect 29316 5404 29326 5460
rect 47954 5404 47964 5460
rect 48020 5404 49252 5460
rect 49746 5404 49756 5460
rect 49812 5404 50988 5460
rect 51044 5404 51054 5460
rect 21084 5348 21140 5404
rect 49196 5348 49252 5404
rect 6626 5292 6636 5348
rect 6692 5292 10108 5348
rect 10164 5292 10174 5348
rect 12898 5292 12908 5348
rect 12964 5292 18060 5348
rect 18116 5292 18126 5348
rect 21084 5292 22764 5348
rect 22820 5292 25676 5348
rect 25732 5292 25742 5348
rect 26338 5292 26348 5348
rect 26404 5292 29596 5348
rect 29652 5292 29662 5348
rect 32386 5292 32396 5348
rect 32452 5292 37100 5348
rect 37156 5292 37166 5348
rect 43484 5292 44268 5348
rect 44324 5292 45388 5348
rect 45444 5292 45454 5348
rect 48962 5292 48972 5348
rect 49028 5292 49038 5348
rect 49196 5292 52108 5348
rect 52164 5292 53116 5348
rect 53172 5292 54684 5348
rect 54740 5292 54750 5348
rect 43484 5236 43540 5292
rect 48972 5236 49028 5292
rect 2034 5180 2044 5236
rect 2100 5180 3948 5236
rect 4004 5180 4014 5236
rect 7858 5180 7868 5236
rect 7924 5180 8988 5236
rect 9044 5180 9054 5236
rect 9202 5180 9212 5236
rect 9268 5180 9772 5236
rect 9828 5180 10444 5236
rect 10500 5180 10510 5236
rect 12450 5180 12460 5236
rect 12516 5180 15036 5236
rect 15092 5180 15102 5236
rect 15260 5180 15596 5236
rect 15652 5180 18508 5236
rect 18564 5180 18574 5236
rect 20290 5180 20300 5236
rect 20356 5180 22540 5236
rect 22596 5180 22606 5236
rect 28578 5180 28588 5236
rect 28644 5180 31612 5236
rect 31668 5180 33068 5236
rect 33124 5180 33134 5236
rect 34514 5180 34524 5236
rect 34580 5180 35756 5236
rect 35812 5180 35822 5236
rect 41794 5180 41804 5236
rect 41860 5180 43484 5236
rect 43540 5180 43550 5236
rect 43698 5180 43708 5236
rect 43764 5180 44828 5236
rect 44884 5180 44894 5236
rect 48972 5180 50764 5236
rect 50820 5180 50830 5236
rect 51660 5180 56252 5236
rect 56308 5180 56924 5236
rect 56980 5180 56990 5236
rect 15260 5124 15316 5180
rect 51660 5124 51716 5180
rect 8194 5068 8204 5124
rect 8260 5068 9548 5124
rect 9604 5068 10780 5124
rect 10836 5068 15316 5124
rect 15810 5068 15820 5124
rect 15876 5068 17388 5124
rect 17444 5068 17454 5124
rect 18610 5068 18620 5124
rect 18676 5068 19292 5124
rect 19348 5068 19358 5124
rect 23090 5068 23100 5124
rect 23156 5068 24332 5124
rect 24388 5068 24398 5124
rect 24994 5068 25004 5124
rect 25060 5068 34972 5124
rect 35028 5068 35038 5124
rect 38770 5068 38780 5124
rect 38836 5068 40348 5124
rect 40404 5068 40414 5124
rect 40674 5068 40684 5124
rect 40740 5068 42364 5124
rect 42420 5068 42430 5124
rect 47170 5068 47180 5124
rect 47236 5068 48076 5124
rect 48132 5068 48142 5124
rect 48738 5068 48748 5124
rect 48804 5068 50204 5124
rect 50260 5068 50270 5124
rect 50372 5068 51436 5124
rect 51492 5068 51502 5124
rect 51650 5068 51660 5124
rect 51716 5068 51726 5124
rect 54002 5068 54012 5124
rect 54068 5068 55692 5124
rect 55748 5068 56588 5124
rect 56644 5068 58044 5124
rect 58100 5068 58110 5124
rect 50372 5012 50428 5068
rect 11004 4956 11340 5012
rect 11396 4956 11406 5012
rect 12786 4956 12796 5012
rect 12852 4956 16828 5012
rect 16884 4956 16894 5012
rect 23202 4956 23212 5012
rect 23268 4956 26572 5012
rect 26628 4956 26638 5012
rect 36082 4956 36092 5012
rect 36148 4956 37548 5012
rect 37604 4956 37614 5012
rect 39890 4956 39900 5012
rect 39956 4956 41020 5012
rect 41076 4956 41086 5012
rect 49298 4956 49308 5012
rect 49364 4956 50428 5012
rect 51202 4956 51212 5012
rect 51268 4956 52220 5012
rect 52276 4956 52286 5012
rect 11004 4900 11060 4956
rect 6402 4844 6412 4900
rect 6468 4844 8092 4900
rect 8148 4844 8158 4900
rect 10994 4844 11004 4900
rect 11060 4844 11070 4900
rect 12674 4844 12684 4900
rect 12740 4844 13580 4900
rect 13636 4844 13646 4900
rect 15138 4844 15148 4900
rect 15204 4844 21084 4900
rect 21140 4844 21150 4900
rect 23986 4844 23996 4900
rect 24052 4844 25116 4900
rect 25172 4844 25452 4900
rect 25508 4844 25518 4900
rect 25666 4844 25676 4900
rect 25732 4844 32396 4900
rect 32452 4844 32462 4900
rect 33618 4844 33628 4900
rect 33684 4844 34524 4900
rect 34580 4844 34590 4900
rect 38546 4844 38556 4900
rect 38612 4844 40236 4900
rect 40292 4844 42700 4900
rect 42756 4844 42766 4900
rect 43708 4844 44716 4900
rect 44772 4844 44782 4900
rect 0 4704 800 4816
rect 43708 4788 43764 4844
rect 11330 4732 11340 4788
rect 11396 4732 13468 4788
rect 13524 4732 13534 4788
rect 17714 4732 17724 4788
rect 17780 4732 28364 4788
rect 28420 4732 28430 4788
rect 29362 4732 29372 4788
rect 29428 4732 29438 4788
rect 39218 4732 39228 4788
rect 39284 4732 43708 4788
rect 43764 4732 43774 4788
rect 15508 4676 15518 4732
rect 15574 4676 15622 4732
rect 15678 4676 15726 4732
rect 15782 4676 15792 4732
rect 29372 4676 29428 4732
rect 29815 4676 29825 4732
rect 29881 4676 29929 4732
rect 29985 4676 30033 4732
rect 30089 4676 30099 4732
rect 44122 4676 44132 4732
rect 44188 4676 44236 4732
rect 44292 4676 44340 4732
rect 44396 4676 44406 4732
rect 58429 4676 58439 4732
rect 58495 4676 58543 4732
rect 58599 4676 58647 4732
rect 58703 4676 58713 4732
rect 11778 4620 11788 4676
rect 11844 4620 15372 4676
rect 15428 4620 15438 4676
rect 15922 4620 15932 4676
rect 15988 4620 18508 4676
rect 18564 4620 19180 4676
rect 19236 4620 19246 4676
rect 22306 4620 22316 4676
rect 22372 4620 25452 4676
rect 25508 4620 25518 4676
rect 25666 4620 25676 4676
rect 25732 4620 29428 4676
rect 37090 4620 37100 4676
rect 37156 4620 38332 4676
rect 38388 4620 40124 4676
rect 40180 4620 40190 4676
rect 41458 4620 41468 4676
rect 41524 4620 42812 4676
rect 42868 4620 43596 4676
rect 43652 4620 43662 4676
rect 8978 4508 8988 4564
rect 9044 4508 18116 4564
rect 18274 4508 18284 4564
rect 18340 4508 21252 4564
rect 22642 4508 22652 4564
rect 22708 4508 24332 4564
rect 24388 4508 24398 4564
rect 24882 4508 24892 4564
rect 24948 4508 28812 4564
rect 28868 4508 28878 4564
rect 30370 4508 30380 4564
rect 30436 4508 32620 4564
rect 32676 4508 34076 4564
rect 34132 4508 34142 4564
rect 34626 4508 34636 4564
rect 34692 4508 56588 4564
rect 56644 4508 56654 4564
rect 10658 4396 10668 4452
rect 10724 4396 12124 4452
rect 12180 4396 12190 4452
rect 12898 4396 12908 4452
rect 12964 4396 12974 4452
rect 13458 4396 13468 4452
rect 13524 4396 14028 4452
rect 14084 4396 14094 4452
rect 15026 4396 15036 4452
rect 15092 4396 16044 4452
rect 16100 4396 16110 4452
rect 11442 4284 11452 4340
rect 11508 4284 11900 4340
rect 11956 4284 11966 4340
rect 12908 4116 12964 4396
rect 18060 4340 18116 4508
rect 21196 4452 21252 4508
rect 19394 4396 19404 4452
rect 19460 4396 20972 4452
rect 21028 4396 21038 4452
rect 21196 4396 25340 4452
rect 25396 4396 25406 4452
rect 25554 4396 25564 4452
rect 25620 4396 27132 4452
rect 27188 4396 27804 4452
rect 27860 4396 27870 4452
rect 30594 4396 30604 4452
rect 30660 4396 33852 4452
rect 33908 4396 33918 4452
rect 37762 4396 37772 4452
rect 37828 4396 38892 4452
rect 38948 4396 38958 4452
rect 43250 4396 43260 4452
rect 43316 4396 46620 4452
rect 46676 4396 47516 4452
rect 47572 4396 47582 4452
rect 51090 4396 51100 4452
rect 51156 4396 51996 4452
rect 52052 4396 52062 4452
rect 15362 4284 15372 4340
rect 15428 4284 17500 4340
rect 17556 4284 17566 4340
rect 18050 4284 18060 4340
rect 18116 4284 18126 4340
rect 19842 4284 19852 4340
rect 19908 4284 20412 4340
rect 20468 4284 20860 4340
rect 20916 4284 20926 4340
rect 21970 4284 21980 4340
rect 22036 4284 29820 4340
rect 29876 4284 29886 4340
rect 33282 4284 33292 4340
rect 33348 4284 34188 4340
rect 34244 4284 34254 4340
rect 39330 4284 39340 4340
rect 39396 4284 40460 4340
rect 40516 4284 40526 4340
rect 41122 4284 41132 4340
rect 41188 4284 41468 4340
rect 41524 4284 42140 4340
rect 42196 4284 42206 4340
rect 13794 4172 13804 4228
rect 13860 4172 16268 4228
rect 16324 4172 16334 4228
rect 16706 4172 16716 4228
rect 16772 4172 20972 4228
rect 21028 4172 22876 4228
rect 22932 4172 22942 4228
rect 26562 4172 26572 4228
rect 26628 4172 27580 4228
rect 27636 4172 27646 4228
rect 27906 4172 27916 4228
rect 27972 4172 29932 4228
rect 29988 4172 29998 4228
rect 32498 4172 32508 4228
rect 32564 4172 40796 4228
rect 40852 4172 42476 4228
rect 42532 4172 43820 4228
rect 43876 4172 43886 4228
rect 45714 4172 45724 4228
rect 45780 4172 47852 4228
rect 47908 4172 47918 4228
rect 8418 4060 8428 4116
rect 8484 4060 11452 4116
rect 11508 4060 11518 4116
rect 12908 4060 19068 4116
rect 19124 4060 19134 4116
rect 27682 4060 27692 4116
rect 27748 4060 28588 4116
rect 28644 4060 28654 4116
rect 29474 4060 29484 4116
rect 29540 4060 37324 4116
rect 37380 4060 37390 4116
rect 28588 4004 28644 4060
rect 10882 3948 10892 4004
rect 10948 3948 10958 4004
rect 11554 3948 11564 4004
rect 11620 3948 13468 4004
rect 13524 3948 13534 4004
rect 15092 3948 15820 4004
rect 15876 3948 15886 4004
rect 17490 3948 17500 4004
rect 17556 3948 22316 4004
rect 22372 3948 22382 4004
rect 28588 3948 34636 4004
rect 34692 3948 34702 4004
rect 8355 3892 8365 3948
rect 8421 3892 8469 3948
rect 8525 3892 8573 3948
rect 8629 3892 8639 3948
rect 10892 3892 10948 3948
rect 15092 3892 15148 3948
rect 22662 3892 22672 3948
rect 22728 3892 22776 3948
rect 22832 3892 22880 3948
rect 22936 3892 22946 3948
rect 36969 3892 36979 3948
rect 37035 3892 37083 3948
rect 37139 3892 37187 3948
rect 37243 3892 37253 3948
rect 51276 3892 51286 3948
rect 51342 3892 51390 3948
rect 51446 3892 51494 3948
rect 51550 3892 51560 3948
rect 10892 3836 15148 3892
rect 7634 3724 7644 3780
rect 7700 3724 10556 3780
rect 10612 3724 12572 3780
rect 12628 3724 12638 3780
rect 16370 3724 16380 3780
rect 16436 3724 21420 3780
rect 21476 3724 21486 3780
rect 28466 3724 28476 3780
rect 28532 3724 29708 3780
rect 29764 3724 29774 3780
rect 29922 3724 29932 3780
rect 29988 3724 34636 3780
rect 34692 3724 34702 3780
rect 44594 3724 44604 3780
rect 44660 3724 45948 3780
rect 46004 3724 46956 3780
rect 47012 3724 47404 3780
rect 47460 3724 47470 3780
rect 0 3584 800 3696
rect 4386 3612 4396 3668
rect 4452 3612 6300 3668
rect 6356 3612 7196 3668
rect 7252 3612 12012 3668
rect 12068 3612 12078 3668
rect 23986 3612 23996 3668
rect 24052 3612 33292 3668
rect 33348 3612 33358 3668
rect 12226 3500 12236 3556
rect 12292 3500 14700 3556
rect 14756 3500 14766 3556
rect 19842 3500 19852 3556
rect 19908 3500 25004 3556
rect 25060 3500 25070 3556
rect 27346 3500 27356 3556
rect 27412 3500 30604 3556
rect 30660 3500 35084 3556
rect 35140 3500 35150 3556
rect 5842 3388 5852 3444
rect 5908 3388 8092 3444
rect 8148 3388 8158 3444
rect 8866 3388 8876 3444
rect 8932 3388 11228 3444
rect 11284 3388 11294 3444
rect 14802 3388 14812 3444
rect 14868 3388 17500 3444
rect 17556 3388 17566 3444
rect 25666 3388 25676 3444
rect 25732 3388 30940 3444
rect 30996 3388 31006 3444
rect 32834 3388 32844 3444
rect 32900 3388 34188 3444
rect 34244 3388 34254 3444
rect 7746 3276 7756 3332
rect 7812 3276 17836 3332
rect 17892 3276 17902 3332
rect 28914 3276 28924 3332
rect 28980 3276 33740 3332
rect 33796 3276 33806 3332
rect 45042 3276 45052 3332
rect 45108 3276 50652 3332
rect 50708 3276 50718 3332
rect 15508 3108 15518 3164
rect 15574 3108 15622 3164
rect 15678 3108 15726 3164
rect 15782 3108 15792 3164
rect 29815 3108 29825 3164
rect 29881 3108 29929 3164
rect 29985 3108 30033 3164
rect 30089 3108 30099 3164
rect 44122 3108 44132 3164
rect 44188 3108 44236 3164
rect 44292 3108 44340 3164
rect 44396 3108 44406 3164
rect 58429 3108 58439 3164
rect 58495 3108 58543 3164
rect 58599 3108 58647 3164
rect 58703 3108 58713 3164
rect 11218 2940 11228 2996
rect 11284 2940 30268 2996
rect 30324 2940 30334 2996
rect 16482 2828 16492 2884
rect 16548 2828 25900 2884
rect 25956 2828 25966 2884
rect 11666 2716 11676 2772
rect 11732 2716 45724 2772
rect 45780 2716 45790 2772
rect 18386 2604 18396 2660
rect 18452 2604 52780 2660
rect 52836 2604 52846 2660
rect 0 2464 800 2576
rect 11106 2492 11116 2548
rect 11172 2492 20748 2548
rect 20804 2492 20814 2548
rect 15250 2380 15260 2436
rect 15316 2380 31276 2436
rect 31332 2380 31342 2436
rect 11106 2268 11116 2324
rect 11172 2268 28924 2324
rect 28980 2268 28990 2324
rect 16594 2156 16604 2212
rect 16660 2156 38444 2212
rect 38500 2156 38510 2212
<< via3 >>
rect 8365 36820 8421 36876
rect 8469 36820 8525 36876
rect 8573 36820 8629 36876
rect 22672 36820 22728 36876
rect 22776 36820 22832 36876
rect 22880 36820 22936 36876
rect 36979 36820 37035 36876
rect 37083 36820 37139 36876
rect 37187 36820 37243 36876
rect 51286 36820 51342 36876
rect 51390 36820 51446 36876
rect 51494 36820 51550 36876
rect 15518 36036 15574 36092
rect 15622 36036 15678 36092
rect 15726 36036 15782 36092
rect 29825 36036 29881 36092
rect 29929 36036 29985 36092
rect 30033 36036 30089 36092
rect 44132 36036 44188 36092
rect 44236 36036 44292 36092
rect 44340 36036 44396 36092
rect 58439 36036 58495 36092
rect 58543 36036 58599 36092
rect 58647 36036 58703 36092
rect 8365 35252 8421 35308
rect 8469 35252 8525 35308
rect 8573 35252 8629 35308
rect 22672 35252 22728 35308
rect 22776 35252 22832 35308
rect 22880 35252 22936 35308
rect 36979 35252 37035 35308
rect 37083 35252 37139 35308
rect 37187 35252 37243 35308
rect 51286 35252 51342 35308
rect 51390 35252 51446 35308
rect 51494 35252 51550 35308
rect 29372 34524 29428 34580
rect 15518 34468 15574 34524
rect 15622 34468 15678 34524
rect 15726 34468 15782 34524
rect 29825 34468 29881 34524
rect 29929 34468 29985 34524
rect 30033 34468 30089 34524
rect 44132 34468 44188 34524
rect 44236 34468 44292 34524
rect 44340 34468 44396 34524
rect 58439 34468 58495 34524
rect 58543 34468 58599 34524
rect 58647 34468 58703 34524
rect 8365 33684 8421 33740
rect 8469 33684 8525 33740
rect 8573 33684 8629 33740
rect 22672 33684 22728 33740
rect 22776 33684 22832 33740
rect 22880 33684 22936 33740
rect 36979 33684 37035 33740
rect 37083 33684 37139 33740
rect 37187 33684 37243 33740
rect 51286 33684 51342 33740
rect 51390 33684 51446 33740
rect 51494 33684 51550 33740
rect 15518 32900 15574 32956
rect 15622 32900 15678 32956
rect 15726 32900 15782 32956
rect 29825 32900 29881 32956
rect 29929 32900 29985 32956
rect 30033 32900 30089 32956
rect 38892 32732 38948 32788
rect 44132 32900 44188 32956
rect 44236 32900 44292 32956
rect 44340 32900 44396 32956
rect 58439 32900 58495 32956
rect 58543 32900 58599 32956
rect 58647 32900 58703 32956
rect 38892 32284 38948 32340
rect 8365 32116 8421 32172
rect 8469 32116 8525 32172
rect 8573 32116 8629 32172
rect 22672 32116 22728 32172
rect 22776 32116 22832 32172
rect 22880 32116 22936 32172
rect 36979 32116 37035 32172
rect 37083 32116 37139 32172
rect 37187 32116 37243 32172
rect 51286 32116 51342 32172
rect 51390 32116 51446 32172
rect 51494 32116 51550 32172
rect 56924 31724 56980 31780
rect 15518 31332 15574 31388
rect 15622 31332 15678 31388
rect 15726 31332 15782 31388
rect 29825 31332 29881 31388
rect 29929 31332 29985 31388
rect 30033 31332 30089 31388
rect 44132 31332 44188 31388
rect 44236 31332 44292 31388
rect 44340 31332 44396 31388
rect 58439 31332 58495 31388
rect 58543 31332 58599 31388
rect 58647 31332 58703 31388
rect 56924 31052 56980 31108
rect 8365 30548 8421 30604
rect 8469 30548 8525 30604
rect 8573 30548 8629 30604
rect 22672 30548 22728 30604
rect 22776 30548 22832 30604
rect 22880 30548 22936 30604
rect 36979 30548 37035 30604
rect 37083 30548 37139 30604
rect 37187 30548 37243 30604
rect 51286 30548 51342 30604
rect 51390 30548 51446 30604
rect 51494 30548 51550 30604
rect 15518 29764 15574 29820
rect 15622 29764 15678 29820
rect 15726 29764 15782 29820
rect 29825 29764 29881 29820
rect 29929 29764 29985 29820
rect 30033 29764 30089 29820
rect 44132 29764 44188 29820
rect 44236 29764 44292 29820
rect 44340 29764 44396 29820
rect 58439 29764 58495 29820
rect 58543 29764 58599 29820
rect 58647 29764 58703 29820
rect 2156 29036 2212 29092
rect 8365 28980 8421 29036
rect 8469 28980 8525 29036
rect 8573 28980 8629 29036
rect 22672 28980 22728 29036
rect 22776 28980 22832 29036
rect 22880 28980 22936 29036
rect 36979 28980 37035 29036
rect 37083 28980 37139 29036
rect 37187 28980 37243 29036
rect 51286 28980 51342 29036
rect 51390 28980 51446 29036
rect 51494 28980 51550 29036
rect 15518 28196 15574 28252
rect 15622 28196 15678 28252
rect 15726 28196 15782 28252
rect 11900 28028 11956 28084
rect 29825 28196 29881 28252
rect 29929 28196 29985 28252
rect 30033 28196 30089 28252
rect 44132 28196 44188 28252
rect 44236 28196 44292 28252
rect 44340 28196 44396 28252
rect 58439 28196 58495 28252
rect 58543 28196 58599 28252
rect 58647 28196 58703 28252
rect 34748 27580 34804 27636
rect 8365 27412 8421 27468
rect 8469 27412 8525 27468
rect 8573 27412 8629 27468
rect 22672 27412 22728 27468
rect 22776 27412 22832 27468
rect 22880 27412 22936 27468
rect 36979 27412 37035 27468
rect 37083 27412 37139 27468
rect 37187 27412 37243 27468
rect 51286 27412 51342 27468
rect 51390 27412 51446 27468
rect 51494 27412 51550 27468
rect 15518 26628 15574 26684
rect 15622 26628 15678 26684
rect 15726 26628 15782 26684
rect 29825 26628 29881 26684
rect 29929 26628 29985 26684
rect 30033 26628 30089 26684
rect 44132 26628 44188 26684
rect 44236 26628 44292 26684
rect 44340 26628 44396 26684
rect 58439 26628 58495 26684
rect 58543 26628 58599 26684
rect 58647 26628 58703 26684
rect 12012 26460 12068 26516
rect 44492 26348 44548 26404
rect 37996 26236 38052 26292
rect 37884 25900 37940 25956
rect 38220 25900 38276 25956
rect 8365 25844 8421 25900
rect 8469 25844 8525 25900
rect 8573 25844 8629 25900
rect 22672 25844 22728 25900
rect 22776 25844 22832 25900
rect 22880 25844 22936 25900
rect 36979 25844 37035 25900
rect 37083 25844 37139 25900
rect 37187 25844 37243 25900
rect 51286 25844 51342 25900
rect 51390 25844 51446 25900
rect 51494 25844 51550 25900
rect 23100 25788 23156 25844
rect 38332 25788 38388 25844
rect 38108 25676 38164 25732
rect 2044 25452 2100 25508
rect 12012 25452 12068 25508
rect 37548 25340 37604 25396
rect 38332 25340 38388 25396
rect 23100 25228 23156 25284
rect 15518 25060 15574 25116
rect 15622 25060 15678 25116
rect 15726 25060 15782 25116
rect 29825 25060 29881 25116
rect 29929 25060 29985 25116
rect 30033 25060 30089 25116
rect 29372 25004 29428 25060
rect 44132 25060 44188 25116
rect 44236 25060 44292 25116
rect 44340 25060 44396 25116
rect 58439 25060 58495 25116
rect 58543 25060 58599 25116
rect 58647 25060 58703 25116
rect 37884 24780 37940 24836
rect 3388 24556 3444 24612
rect 44492 24668 44548 24724
rect 37548 24556 37604 24612
rect 38108 24556 38164 24612
rect 56924 24444 56980 24500
rect 38220 24332 38276 24388
rect 44716 24332 44772 24388
rect 8365 24276 8421 24332
rect 8469 24276 8525 24332
rect 8573 24276 8629 24332
rect 22672 24276 22728 24332
rect 22776 24276 22832 24332
rect 22880 24276 22936 24332
rect 36979 24276 37035 24332
rect 37083 24276 37139 24332
rect 37187 24276 37243 24332
rect 51286 24276 51342 24332
rect 51390 24276 51446 24332
rect 51494 24276 51550 24332
rect 11900 23772 11956 23828
rect 12012 23660 12068 23716
rect 37548 23660 37604 23716
rect 37996 23660 38052 23716
rect 50540 23660 50596 23716
rect 15518 23492 15574 23548
rect 15622 23492 15678 23548
rect 15726 23492 15782 23548
rect 29825 23492 29881 23548
rect 29929 23492 29985 23548
rect 30033 23492 30089 23548
rect 44132 23492 44188 23548
rect 44236 23492 44292 23548
rect 44340 23492 44396 23548
rect 58439 23492 58495 23548
rect 58543 23492 58599 23548
rect 58647 23492 58703 23548
rect 44716 23436 44772 23492
rect 45276 23436 45332 23492
rect 9212 23212 9268 23268
rect 14028 23212 14084 23268
rect 33180 23100 33236 23156
rect 45276 23100 45332 23156
rect 13804 22876 13860 22932
rect 32060 22876 32116 22932
rect 8365 22708 8421 22764
rect 8469 22708 8525 22764
rect 8573 22708 8629 22764
rect 22672 22708 22728 22764
rect 22776 22708 22832 22764
rect 22880 22708 22936 22764
rect 36979 22708 37035 22764
rect 37083 22708 37139 22764
rect 37187 22708 37243 22764
rect 51286 22708 51342 22764
rect 51390 22708 51446 22764
rect 51494 22708 51550 22764
rect 37996 22652 38052 22708
rect 7196 22428 7252 22484
rect 3724 22204 3780 22260
rect 46060 22204 46116 22260
rect 14140 22092 14196 22148
rect 31948 22092 32004 22148
rect 2828 21980 2884 22036
rect 14028 21980 14084 22036
rect 4284 21868 4340 21924
rect 15518 21924 15574 21980
rect 15622 21924 15678 21980
rect 15726 21924 15782 21980
rect 29825 21924 29881 21980
rect 29929 21924 29985 21980
rect 30033 21924 30089 21980
rect 44132 21924 44188 21980
rect 44236 21924 44292 21980
rect 44340 21924 44396 21980
rect 33516 21756 33572 21812
rect 58439 21924 58495 21980
rect 58543 21924 58599 21980
rect 58647 21924 58703 21980
rect 3388 21532 3444 21588
rect 47068 21532 47124 21588
rect 48300 21532 48356 21588
rect 32060 21420 32116 21476
rect 33180 21196 33236 21252
rect 8365 21140 8421 21196
rect 8469 21140 8525 21196
rect 8573 21140 8629 21196
rect 22672 21140 22728 21196
rect 22776 21140 22832 21196
rect 22880 21140 22936 21196
rect 31948 21084 32004 21140
rect 33516 21084 33572 21140
rect 36979 21140 37035 21196
rect 37083 21140 37139 21196
rect 37187 21140 37243 21196
rect 51286 21140 51342 21196
rect 51390 21140 51446 21196
rect 51494 21140 51550 21196
rect 37996 21084 38052 21140
rect 49084 20860 49140 20916
rect 32172 20636 32228 20692
rect 15518 20356 15574 20412
rect 15622 20356 15678 20412
rect 15726 20356 15782 20412
rect 29825 20356 29881 20412
rect 29929 20356 29985 20412
rect 30033 20356 30089 20412
rect 44132 20356 44188 20412
rect 44236 20356 44292 20412
rect 44340 20356 44396 20412
rect 58439 20356 58495 20412
rect 58543 20356 58599 20412
rect 58647 20356 58703 20412
rect 8988 20188 9044 20244
rect 28140 20076 28196 20132
rect 46060 19852 46116 19908
rect 50540 19628 50596 19684
rect 8365 19572 8421 19628
rect 8469 19572 8525 19628
rect 8573 19572 8629 19628
rect 22672 19572 22728 19628
rect 22776 19572 22832 19628
rect 22880 19572 22936 19628
rect 36979 19572 37035 19628
rect 37083 19572 37139 19628
rect 37187 19572 37243 19628
rect 51286 19572 51342 19628
rect 51390 19572 51446 19628
rect 51494 19572 51550 19628
rect 9212 19292 9268 19348
rect 35644 19068 35700 19124
rect 3500 18844 3556 18900
rect 36428 18844 36484 18900
rect 15518 18788 15574 18844
rect 15622 18788 15678 18844
rect 15726 18788 15782 18844
rect 29825 18788 29881 18844
rect 29929 18788 29985 18844
rect 30033 18788 30089 18844
rect 49084 18844 49140 18900
rect 44132 18788 44188 18844
rect 44236 18788 44292 18844
rect 44340 18788 44396 18844
rect 58439 18788 58495 18844
rect 58543 18788 58599 18844
rect 58647 18788 58703 18844
rect 13580 18620 13636 18676
rect 36764 18620 36820 18676
rect 12348 18284 12404 18340
rect 42924 18284 42980 18340
rect 8365 18004 8421 18060
rect 8469 18004 8525 18060
rect 8573 18004 8629 18060
rect 22672 18004 22728 18060
rect 22776 18004 22832 18060
rect 22880 18004 22936 18060
rect 36979 18004 37035 18060
rect 37083 18004 37139 18060
rect 37187 18004 37243 18060
rect 51286 18004 51342 18060
rect 51390 18004 51446 18060
rect 51494 18004 51550 18060
rect 45164 17948 45220 18004
rect 47068 17948 47124 18004
rect 47516 17948 47572 18004
rect 7196 17724 7252 17780
rect 13580 17500 13636 17556
rect 35644 17500 35700 17556
rect 2828 17276 2884 17332
rect 16044 17276 16100 17332
rect 15518 17220 15574 17276
rect 15622 17220 15678 17276
rect 15726 17220 15782 17276
rect 29825 17220 29881 17276
rect 29929 17220 29985 17276
rect 30033 17220 30089 17276
rect 44132 17220 44188 17276
rect 44236 17220 44292 17276
rect 44340 17220 44396 17276
rect 58439 17220 58495 17276
rect 58543 17220 58599 17276
rect 58647 17220 58703 17276
rect 26908 17164 26964 17220
rect 42812 16828 42868 16884
rect 36428 16716 36484 16772
rect 36764 16716 36820 16772
rect 48748 16604 48804 16660
rect 49196 16604 49252 16660
rect 8365 16436 8421 16492
rect 8469 16436 8525 16492
rect 8573 16436 8629 16492
rect 22672 16436 22728 16492
rect 22776 16436 22832 16492
rect 22880 16436 22936 16492
rect 36979 16436 37035 16492
rect 37083 16436 37139 16492
rect 37187 16436 37243 16492
rect 51286 16436 51342 16492
rect 51390 16436 51446 16492
rect 51494 16436 51550 16492
rect 34748 16380 34804 16436
rect 3500 16156 3556 16212
rect 13580 16156 13636 16212
rect 23324 16044 23380 16100
rect 8988 15820 9044 15876
rect 47516 15820 47572 15876
rect 15518 15652 15574 15708
rect 15622 15652 15678 15708
rect 15726 15652 15782 15708
rect 28140 15596 28196 15652
rect 29825 15652 29881 15708
rect 29929 15652 29985 15708
rect 30033 15652 30089 15708
rect 44132 15652 44188 15708
rect 44236 15652 44292 15708
rect 44340 15652 44396 15708
rect 58439 15652 58495 15708
rect 58543 15652 58599 15708
rect 58647 15652 58703 15708
rect 45164 15596 45220 15652
rect 16044 15484 16100 15540
rect 34748 15372 34804 15428
rect 23100 15148 23156 15204
rect 8988 14924 9044 14980
rect 8365 14868 8421 14924
rect 8469 14868 8525 14924
rect 8573 14868 8629 14924
rect 22672 14868 22728 14924
rect 22776 14868 22832 14924
rect 22880 14868 22936 14924
rect 36979 14868 37035 14924
rect 37083 14868 37139 14924
rect 37187 14868 37243 14924
rect 51286 14868 51342 14924
rect 51390 14868 51446 14924
rect 51494 14868 51550 14924
rect 23100 14812 23156 14868
rect 26908 14700 26964 14756
rect 4284 14588 4340 14644
rect 14140 14364 14196 14420
rect 42812 14140 42868 14196
rect 48300 14140 48356 14196
rect 15518 14084 15574 14140
rect 15622 14084 15678 14140
rect 15726 14084 15782 14140
rect 29825 14084 29881 14140
rect 29929 14084 29985 14140
rect 30033 14084 30089 14140
rect 44132 14084 44188 14140
rect 44236 14084 44292 14140
rect 44340 14084 44396 14140
rect 58439 14084 58495 14140
rect 58543 14084 58599 14140
rect 58647 14084 58703 14140
rect 32172 14028 32228 14084
rect 2044 13916 2100 13972
rect 3500 13916 3556 13972
rect 42924 13804 42980 13860
rect 12348 13356 12404 13412
rect 23324 13356 23380 13412
rect 8365 13300 8421 13356
rect 8469 13300 8525 13356
rect 8573 13300 8629 13356
rect 22672 13300 22728 13356
rect 22776 13300 22832 13356
rect 22880 13300 22936 13356
rect 36979 13300 37035 13356
rect 37083 13300 37139 13356
rect 37187 13300 37243 13356
rect 51286 13300 51342 13356
rect 51390 13300 51446 13356
rect 51494 13300 51550 13356
rect 23436 13244 23492 13300
rect 23436 13020 23492 13076
rect 46060 12908 46116 12964
rect 3724 12796 3780 12852
rect 15518 12516 15574 12572
rect 15622 12516 15678 12572
rect 15726 12516 15782 12572
rect 29825 12516 29881 12572
rect 29929 12516 29985 12572
rect 30033 12516 30089 12572
rect 44132 12516 44188 12572
rect 44236 12516 44292 12572
rect 44340 12516 44396 12572
rect 58439 12516 58495 12572
rect 58543 12516 58599 12572
rect 58647 12516 58703 12572
rect 13804 12348 13860 12404
rect 46060 11788 46116 11844
rect 8365 11732 8421 11788
rect 8469 11732 8525 11788
rect 8573 11732 8629 11788
rect 22672 11732 22728 11788
rect 22776 11732 22832 11788
rect 22880 11732 22936 11788
rect 36979 11732 37035 11788
rect 37083 11732 37139 11788
rect 37187 11732 37243 11788
rect 51286 11732 51342 11788
rect 51390 11732 51446 11788
rect 51494 11732 51550 11788
rect 34300 11676 34356 11732
rect 26684 11452 26740 11508
rect 27020 11452 27076 11508
rect 34300 11116 34356 11172
rect 35308 11116 35364 11172
rect 15518 10948 15574 11004
rect 15622 10948 15678 11004
rect 15726 10948 15782 11004
rect 29825 10948 29881 11004
rect 29929 10948 29985 11004
rect 30033 10948 30089 11004
rect 30268 10892 30324 10948
rect 44132 10948 44188 11004
rect 44236 10948 44292 11004
rect 44340 10948 44396 11004
rect 58439 10948 58495 11004
rect 58543 10948 58599 11004
rect 58647 10948 58703 11004
rect 23100 10668 23156 10724
rect 34524 10556 34580 10612
rect 34636 10444 34692 10500
rect 41244 10444 41300 10500
rect 41468 10444 41524 10500
rect 30268 10332 30324 10388
rect 43036 10220 43092 10276
rect 8365 10164 8421 10220
rect 8469 10164 8525 10220
rect 8573 10164 8629 10220
rect 22672 10164 22728 10220
rect 22776 10164 22832 10220
rect 22880 10164 22936 10220
rect 36979 10164 37035 10220
rect 37083 10164 37139 10220
rect 37187 10164 37243 10220
rect 51286 10164 51342 10220
rect 51390 10164 51446 10220
rect 51494 10164 51550 10220
rect 35308 9996 35364 10052
rect 45948 9996 46004 10052
rect 26852 9548 26908 9604
rect 15518 9380 15574 9436
rect 15622 9380 15678 9436
rect 15726 9380 15782 9436
rect 29825 9380 29881 9436
rect 29929 9380 29985 9436
rect 30033 9380 30089 9436
rect 44132 9380 44188 9436
rect 44236 9380 44292 9436
rect 44340 9380 44396 9436
rect 58439 9380 58495 9436
rect 58543 9380 58599 9436
rect 58647 9380 58703 9436
rect 46060 9212 46116 9268
rect 26908 8988 26964 9044
rect 41244 8988 41300 9044
rect 34636 8876 34692 8932
rect 43036 8764 43092 8820
rect 8365 8596 8421 8652
rect 8469 8596 8525 8652
rect 8573 8596 8629 8652
rect 22672 8596 22728 8652
rect 22776 8596 22832 8652
rect 22880 8596 22936 8652
rect 36979 8596 37035 8652
rect 37083 8596 37139 8652
rect 37187 8596 37243 8652
rect 51286 8596 51342 8652
rect 51390 8596 51446 8652
rect 51494 8596 51550 8652
rect 23100 8316 23156 8372
rect 46060 7868 46116 7924
rect 15518 7812 15574 7868
rect 15622 7812 15678 7868
rect 15726 7812 15782 7868
rect 29825 7812 29881 7868
rect 29929 7812 29985 7868
rect 30033 7812 30089 7868
rect 44132 7812 44188 7868
rect 44236 7812 44292 7868
rect 44340 7812 44396 7868
rect 58439 7812 58495 7868
rect 58543 7812 58599 7868
rect 58647 7812 58703 7868
rect 34524 7756 34580 7812
rect 8365 7028 8421 7084
rect 8469 7028 8525 7084
rect 8573 7028 8629 7084
rect 22672 7028 22728 7084
rect 22776 7028 22832 7084
rect 22880 7028 22936 7084
rect 36979 7028 37035 7084
rect 37083 7028 37139 7084
rect 37187 7028 37243 7084
rect 51286 7028 51342 7084
rect 51390 7028 51446 7084
rect 51494 7028 51550 7084
rect 45948 6748 46004 6804
rect 15518 6244 15574 6300
rect 15622 6244 15678 6300
rect 15726 6244 15782 6300
rect 29825 6244 29881 6300
rect 29929 6244 29985 6300
rect 30033 6244 30089 6300
rect 44132 6244 44188 6300
rect 44236 6244 44292 6300
rect 44340 6244 44396 6300
rect 58439 6244 58495 6300
rect 58543 6244 58599 6300
rect 58647 6244 58703 6300
rect 34300 5852 34356 5908
rect 8365 5460 8421 5516
rect 8469 5460 8525 5516
rect 8573 5460 8629 5516
rect 22672 5460 22728 5516
rect 22776 5460 22832 5516
rect 22880 5460 22936 5516
rect 36979 5460 37035 5516
rect 37083 5460 37139 5516
rect 37187 5460 37243 5516
rect 51286 5460 51342 5516
rect 51390 5460 51446 5516
rect 51494 5460 51550 5516
rect 25676 4844 25732 4900
rect 15518 4676 15574 4732
rect 15622 4676 15678 4732
rect 15726 4676 15782 4732
rect 29825 4676 29881 4732
rect 29929 4676 29985 4732
rect 30033 4676 30089 4732
rect 44132 4676 44188 4732
rect 44236 4676 44292 4732
rect 44340 4676 44396 4732
rect 58439 4676 58495 4732
rect 58543 4676 58599 4732
rect 58647 4676 58703 4732
rect 15372 4620 15428 4676
rect 25340 4396 25396 4452
rect 15372 4284 15428 4340
rect 41468 4284 41524 4340
rect 8365 3892 8421 3948
rect 8469 3892 8525 3948
rect 8573 3892 8629 3948
rect 22672 3892 22728 3948
rect 22776 3892 22832 3948
rect 22880 3892 22936 3948
rect 36979 3892 37035 3948
rect 37083 3892 37139 3948
rect 37187 3892 37243 3948
rect 51286 3892 51342 3948
rect 51390 3892 51446 3948
rect 51494 3892 51550 3948
rect 15518 3108 15574 3164
rect 15622 3108 15678 3164
rect 15726 3108 15782 3164
rect 29825 3108 29881 3164
rect 29929 3108 29985 3164
rect 30033 3108 30089 3164
rect 44132 3108 44188 3164
rect 44236 3108 44292 3164
rect 44340 3108 44396 3164
rect 58439 3108 58495 3164
rect 58543 3108 58599 3164
rect 58647 3108 58703 3164
<< metal4 >>
rect 8337 36876 8657 36908
rect 8337 36820 8365 36876
rect 8421 36820 8469 36876
rect 8525 36820 8573 36876
rect 8629 36820 8657 36876
rect 8337 35308 8657 36820
rect 8337 35252 8365 35308
rect 8421 35252 8469 35308
rect 8525 35252 8573 35308
rect 8629 35252 8657 35308
rect 8337 33740 8657 35252
rect 8337 33684 8365 33740
rect 8421 33684 8469 33740
rect 8525 33684 8573 33740
rect 8629 33684 8657 33740
rect 8337 32172 8657 33684
rect 8337 32116 8365 32172
rect 8421 32116 8469 32172
rect 8525 32116 8573 32172
rect 8629 32116 8657 32172
rect 8337 30604 8657 32116
rect 8337 30548 8365 30604
rect 8421 30548 8469 30604
rect 8525 30548 8573 30604
rect 8629 30548 8657 30604
rect 2156 29092 2212 29102
rect 2156 26908 2212 29036
rect 2044 26852 2212 26908
rect 8337 29036 8657 30548
rect 8337 28980 8365 29036
rect 8421 28980 8469 29036
rect 8525 28980 8573 29036
rect 8629 28980 8657 29036
rect 8337 27468 8657 28980
rect 15490 36092 15810 36908
rect 15490 36036 15518 36092
rect 15574 36036 15622 36092
rect 15678 36036 15726 36092
rect 15782 36036 15810 36092
rect 15490 34524 15810 36036
rect 15490 34468 15518 34524
rect 15574 34468 15622 34524
rect 15678 34468 15726 34524
rect 15782 34468 15810 34524
rect 15490 32956 15810 34468
rect 15490 32900 15518 32956
rect 15574 32900 15622 32956
rect 15678 32900 15726 32956
rect 15782 32900 15810 32956
rect 15490 31388 15810 32900
rect 15490 31332 15518 31388
rect 15574 31332 15622 31388
rect 15678 31332 15726 31388
rect 15782 31332 15810 31388
rect 15490 29820 15810 31332
rect 15490 29764 15518 29820
rect 15574 29764 15622 29820
rect 15678 29764 15726 29820
rect 15782 29764 15810 29820
rect 15490 28252 15810 29764
rect 15490 28196 15518 28252
rect 15574 28196 15622 28252
rect 15678 28196 15726 28252
rect 15782 28196 15810 28252
rect 8337 27412 8365 27468
rect 8421 27412 8469 27468
rect 8525 27412 8573 27468
rect 8629 27412 8657 27468
rect 2044 25508 2100 26852
rect 2044 13972 2100 25452
rect 8337 25900 8657 27412
rect 8337 25844 8365 25900
rect 8421 25844 8469 25900
rect 8525 25844 8573 25900
rect 8629 25844 8657 25900
rect 3388 24612 3444 24622
rect 2828 22036 2884 22046
rect 2828 17332 2884 21980
rect 3388 21588 3444 24556
rect 8337 24332 8657 25844
rect 8337 24276 8365 24332
rect 8421 24276 8469 24332
rect 8525 24276 8573 24332
rect 8629 24276 8657 24332
rect 8337 22764 8657 24276
rect 11900 28084 11956 28094
rect 11900 23828 11956 28028
rect 15490 26684 15810 28196
rect 15490 26628 15518 26684
rect 15574 26628 15622 26684
rect 15678 26628 15726 26684
rect 15782 26628 15810 26684
rect 11900 23762 11956 23772
rect 12012 26516 12068 26526
rect 12012 25508 12068 26460
rect 12012 23716 12068 25452
rect 12012 23650 12068 23660
rect 15490 25116 15810 26628
rect 15490 25060 15518 25116
rect 15574 25060 15622 25116
rect 15678 25060 15726 25116
rect 15782 25060 15810 25116
rect 15490 23548 15810 25060
rect 15490 23492 15518 23548
rect 15574 23492 15622 23548
rect 15678 23492 15726 23548
rect 15782 23492 15810 23548
rect 8337 22708 8365 22764
rect 8421 22708 8469 22764
rect 8525 22708 8573 22764
rect 8629 22708 8657 22764
rect 7196 22484 7252 22494
rect 3388 21522 3444 21532
rect 3724 22260 3780 22270
rect 2828 17266 2884 17276
rect 3500 18900 3556 18910
rect 2044 13906 2100 13916
rect 3500 16212 3556 18844
rect 3500 13972 3556 16156
rect 3500 13906 3556 13916
rect 3724 12852 3780 22204
rect 4284 21924 4340 21934
rect 4284 14644 4340 21868
rect 7196 17780 7252 22428
rect 7196 17714 7252 17724
rect 8337 21196 8657 22708
rect 8337 21140 8365 21196
rect 8421 21140 8469 21196
rect 8525 21140 8573 21196
rect 8629 21140 8657 21196
rect 8337 19628 8657 21140
rect 9212 23268 9268 23278
rect 8337 19572 8365 19628
rect 8421 19572 8469 19628
rect 8525 19572 8573 19628
rect 8629 19572 8657 19628
rect 8337 18060 8657 19572
rect 8337 18004 8365 18060
rect 8421 18004 8469 18060
rect 8525 18004 8573 18060
rect 8629 18004 8657 18060
rect 4284 14578 4340 14588
rect 8337 16492 8657 18004
rect 8337 16436 8365 16492
rect 8421 16436 8469 16492
rect 8525 16436 8573 16492
rect 8629 16436 8657 16492
rect 8337 14924 8657 16436
rect 8337 14868 8365 14924
rect 8421 14868 8469 14924
rect 8525 14868 8573 14924
rect 8629 14868 8657 14924
rect 8988 20244 9044 20254
rect 8988 15876 9044 20188
rect 9212 19348 9268 23212
rect 14028 23268 14084 23278
rect 9212 19282 9268 19292
rect 13804 22932 13860 22942
rect 13580 18676 13636 18686
rect 8988 14980 9044 15820
rect 8988 14914 9044 14924
rect 12348 18340 12404 18350
rect 3724 12786 3780 12796
rect 8337 13356 8657 14868
rect 8337 13300 8365 13356
rect 8421 13300 8469 13356
rect 8525 13300 8573 13356
rect 8629 13300 8657 13356
rect 12348 13412 12404 18284
rect 13580 17556 13636 18620
rect 13580 16212 13636 17500
rect 13580 16146 13636 16156
rect 12348 13346 12404 13356
rect 8337 11788 8657 13300
rect 13804 12404 13860 22876
rect 14028 22036 14084 23212
rect 14028 21970 14084 21980
rect 14140 22148 14196 22158
rect 14140 14420 14196 22092
rect 14140 14354 14196 14364
rect 15490 21980 15810 23492
rect 15490 21924 15518 21980
rect 15574 21924 15622 21980
rect 15678 21924 15726 21980
rect 15782 21924 15810 21980
rect 15490 20412 15810 21924
rect 15490 20356 15518 20412
rect 15574 20356 15622 20412
rect 15678 20356 15726 20412
rect 15782 20356 15810 20412
rect 15490 18844 15810 20356
rect 15490 18788 15518 18844
rect 15574 18788 15622 18844
rect 15678 18788 15726 18844
rect 15782 18788 15810 18844
rect 15490 17276 15810 18788
rect 22644 36876 22964 36908
rect 22644 36820 22672 36876
rect 22728 36820 22776 36876
rect 22832 36820 22880 36876
rect 22936 36820 22964 36876
rect 22644 35308 22964 36820
rect 22644 35252 22672 35308
rect 22728 35252 22776 35308
rect 22832 35252 22880 35308
rect 22936 35252 22964 35308
rect 22644 33740 22964 35252
rect 29797 36092 30117 36908
rect 29797 36036 29825 36092
rect 29881 36036 29929 36092
rect 29985 36036 30033 36092
rect 30089 36036 30117 36092
rect 22644 33684 22672 33740
rect 22728 33684 22776 33740
rect 22832 33684 22880 33740
rect 22936 33684 22964 33740
rect 22644 32172 22964 33684
rect 22644 32116 22672 32172
rect 22728 32116 22776 32172
rect 22832 32116 22880 32172
rect 22936 32116 22964 32172
rect 22644 30604 22964 32116
rect 22644 30548 22672 30604
rect 22728 30548 22776 30604
rect 22832 30548 22880 30604
rect 22936 30548 22964 30604
rect 22644 29036 22964 30548
rect 22644 28980 22672 29036
rect 22728 28980 22776 29036
rect 22832 28980 22880 29036
rect 22936 28980 22964 29036
rect 22644 27468 22964 28980
rect 22644 27412 22672 27468
rect 22728 27412 22776 27468
rect 22832 27412 22880 27468
rect 22936 27412 22964 27468
rect 22644 25900 22964 27412
rect 22644 25844 22672 25900
rect 22728 25844 22776 25900
rect 22832 25844 22880 25900
rect 22936 25844 22964 25900
rect 29372 34580 29428 34590
rect 22644 24332 22964 25844
rect 23100 25844 23156 25854
rect 23100 25284 23156 25788
rect 23100 25218 23156 25228
rect 29372 25060 29428 34524
rect 29372 24994 29428 25004
rect 29797 34524 30117 36036
rect 29797 34468 29825 34524
rect 29881 34468 29929 34524
rect 29985 34468 30033 34524
rect 30089 34468 30117 34524
rect 29797 32956 30117 34468
rect 29797 32900 29825 32956
rect 29881 32900 29929 32956
rect 29985 32900 30033 32956
rect 30089 32900 30117 32956
rect 29797 31388 30117 32900
rect 29797 31332 29825 31388
rect 29881 31332 29929 31388
rect 29985 31332 30033 31388
rect 30089 31332 30117 31388
rect 29797 29820 30117 31332
rect 29797 29764 29825 29820
rect 29881 29764 29929 29820
rect 29985 29764 30033 29820
rect 30089 29764 30117 29820
rect 29797 28252 30117 29764
rect 29797 28196 29825 28252
rect 29881 28196 29929 28252
rect 29985 28196 30033 28252
rect 30089 28196 30117 28252
rect 29797 26684 30117 28196
rect 36951 36876 37271 36908
rect 36951 36820 36979 36876
rect 37035 36820 37083 36876
rect 37139 36820 37187 36876
rect 37243 36820 37271 36876
rect 36951 35308 37271 36820
rect 36951 35252 36979 35308
rect 37035 35252 37083 35308
rect 37139 35252 37187 35308
rect 37243 35252 37271 35308
rect 36951 33740 37271 35252
rect 36951 33684 36979 33740
rect 37035 33684 37083 33740
rect 37139 33684 37187 33740
rect 37243 33684 37271 33740
rect 36951 32172 37271 33684
rect 44104 36092 44424 36908
rect 44104 36036 44132 36092
rect 44188 36036 44236 36092
rect 44292 36036 44340 36092
rect 44396 36036 44424 36092
rect 44104 34524 44424 36036
rect 44104 34468 44132 34524
rect 44188 34468 44236 34524
rect 44292 34468 44340 34524
rect 44396 34468 44424 34524
rect 44104 32956 44424 34468
rect 44104 32900 44132 32956
rect 44188 32900 44236 32956
rect 44292 32900 44340 32956
rect 44396 32900 44424 32956
rect 38892 32788 38948 32798
rect 38892 32340 38948 32732
rect 38892 32274 38948 32284
rect 36951 32116 36979 32172
rect 37035 32116 37083 32172
rect 37139 32116 37187 32172
rect 37243 32116 37271 32172
rect 36951 30604 37271 32116
rect 36951 30548 36979 30604
rect 37035 30548 37083 30604
rect 37139 30548 37187 30604
rect 37243 30548 37271 30604
rect 36951 29036 37271 30548
rect 36951 28980 36979 29036
rect 37035 28980 37083 29036
rect 37139 28980 37187 29036
rect 37243 28980 37271 29036
rect 29797 26628 29825 26684
rect 29881 26628 29929 26684
rect 29985 26628 30033 26684
rect 30089 26628 30117 26684
rect 29797 25116 30117 26628
rect 29797 25060 29825 25116
rect 29881 25060 29929 25116
rect 29985 25060 30033 25116
rect 30089 25060 30117 25116
rect 22644 24276 22672 24332
rect 22728 24276 22776 24332
rect 22832 24276 22880 24332
rect 22936 24276 22964 24332
rect 22644 22764 22964 24276
rect 22644 22708 22672 22764
rect 22728 22708 22776 22764
rect 22832 22708 22880 22764
rect 22936 22708 22964 22764
rect 22644 21196 22964 22708
rect 22644 21140 22672 21196
rect 22728 21140 22776 21196
rect 22832 21140 22880 21196
rect 22936 21140 22964 21196
rect 22644 19628 22964 21140
rect 29797 23548 30117 25060
rect 29797 23492 29825 23548
rect 29881 23492 29929 23548
rect 29985 23492 30033 23548
rect 30089 23492 30117 23548
rect 29797 21980 30117 23492
rect 34748 27636 34804 27646
rect 33180 23156 33236 23166
rect 32060 22932 32116 22942
rect 29797 21924 29825 21980
rect 29881 21924 29929 21980
rect 29985 21924 30033 21980
rect 30089 21924 30117 21980
rect 29797 20412 30117 21924
rect 31948 22148 32004 22158
rect 31948 21140 32004 22092
rect 32060 21476 32116 22876
rect 32060 21410 32116 21420
rect 33180 21252 33236 23100
rect 33180 21186 33236 21196
rect 33516 21812 33572 21822
rect 31948 21074 32004 21084
rect 33516 21140 33572 21756
rect 33516 21074 33572 21084
rect 29797 20356 29825 20412
rect 29881 20356 29929 20412
rect 29985 20356 30033 20412
rect 30089 20356 30117 20412
rect 22644 19572 22672 19628
rect 22728 19572 22776 19628
rect 22832 19572 22880 19628
rect 22936 19572 22964 19628
rect 22644 18060 22964 19572
rect 22644 18004 22672 18060
rect 22728 18004 22776 18060
rect 22832 18004 22880 18060
rect 22936 18004 22964 18060
rect 15490 17220 15518 17276
rect 15574 17220 15622 17276
rect 15678 17220 15726 17276
rect 15782 17220 15810 17276
rect 15490 15708 15810 17220
rect 15490 15652 15518 15708
rect 15574 15652 15622 15708
rect 15678 15652 15726 15708
rect 15782 15652 15810 15708
rect 13804 12338 13860 12348
rect 15490 14140 15810 15652
rect 16044 17332 16100 17342
rect 16044 15540 16100 17276
rect 16044 15474 16100 15484
rect 22644 16492 22964 18004
rect 28140 20132 28196 20142
rect 22644 16436 22672 16492
rect 22728 16436 22776 16492
rect 22832 16436 22880 16492
rect 22936 16436 22964 16492
rect 15490 14084 15518 14140
rect 15574 14084 15622 14140
rect 15678 14084 15726 14140
rect 15782 14084 15810 14140
rect 15490 12572 15810 14084
rect 15490 12516 15518 12572
rect 15574 12516 15622 12572
rect 15678 12516 15726 12572
rect 15782 12516 15810 12572
rect 8337 11732 8365 11788
rect 8421 11732 8469 11788
rect 8525 11732 8573 11788
rect 8629 11732 8657 11788
rect 8337 10220 8657 11732
rect 8337 10164 8365 10220
rect 8421 10164 8469 10220
rect 8525 10164 8573 10220
rect 8629 10164 8657 10220
rect 8337 8652 8657 10164
rect 8337 8596 8365 8652
rect 8421 8596 8469 8652
rect 8525 8596 8573 8652
rect 8629 8596 8657 8652
rect 8337 7084 8657 8596
rect 8337 7028 8365 7084
rect 8421 7028 8469 7084
rect 8525 7028 8573 7084
rect 8629 7028 8657 7084
rect 8337 5516 8657 7028
rect 8337 5460 8365 5516
rect 8421 5460 8469 5516
rect 8525 5460 8573 5516
rect 8629 5460 8657 5516
rect 8337 3948 8657 5460
rect 15490 11004 15810 12516
rect 15490 10948 15518 11004
rect 15574 10948 15622 11004
rect 15678 10948 15726 11004
rect 15782 10948 15810 11004
rect 15490 9436 15810 10948
rect 15490 9380 15518 9436
rect 15574 9380 15622 9436
rect 15678 9380 15726 9436
rect 15782 9380 15810 9436
rect 15490 7868 15810 9380
rect 15490 7812 15518 7868
rect 15574 7812 15622 7868
rect 15678 7812 15726 7868
rect 15782 7812 15810 7868
rect 15490 6300 15810 7812
rect 15490 6244 15518 6300
rect 15574 6244 15622 6300
rect 15678 6244 15726 6300
rect 15782 6244 15810 6300
rect 15490 4732 15810 6244
rect 15372 4676 15428 4686
rect 15372 4340 15428 4620
rect 15372 4274 15428 4284
rect 15490 4676 15518 4732
rect 15574 4676 15622 4732
rect 15678 4676 15726 4732
rect 15782 4676 15810 4732
rect 8337 3892 8365 3948
rect 8421 3892 8469 3948
rect 8525 3892 8573 3948
rect 8629 3892 8657 3948
rect 8337 3076 8657 3892
rect 15490 3164 15810 4676
rect 15490 3108 15518 3164
rect 15574 3108 15622 3164
rect 15678 3108 15726 3164
rect 15782 3108 15810 3164
rect 15490 3076 15810 3108
rect 22644 14924 22964 16436
rect 26908 17220 26964 17230
rect 23324 16100 23380 16110
rect 22644 14868 22672 14924
rect 22728 14868 22776 14924
rect 22832 14868 22880 14924
rect 22936 14868 22964 14924
rect 22644 13356 22964 14868
rect 23100 15204 23156 15214
rect 23100 14868 23156 15148
rect 23100 14802 23156 14812
rect 22644 13300 22672 13356
rect 22728 13300 22776 13356
rect 22832 13300 22880 13356
rect 22936 13300 22964 13356
rect 23324 13412 23380 16044
rect 26908 14756 26964 17164
rect 28140 15652 28196 20076
rect 28140 15586 28196 15596
rect 29797 18844 30117 20356
rect 29797 18788 29825 18844
rect 29881 18788 29929 18844
rect 29985 18788 30033 18844
rect 30089 18788 30117 18844
rect 29797 17276 30117 18788
rect 29797 17220 29825 17276
rect 29881 17220 29929 17276
rect 29985 17220 30033 17276
rect 30089 17220 30117 17276
rect 29797 15708 30117 17220
rect 29797 15652 29825 15708
rect 29881 15652 29929 15708
rect 29985 15652 30033 15708
rect 30089 15652 30117 15708
rect 26908 14690 26964 14700
rect 23324 13346 23380 13356
rect 29797 14140 30117 15652
rect 29797 14084 29825 14140
rect 29881 14084 29929 14140
rect 29985 14084 30033 14140
rect 30089 14084 30117 14140
rect 22644 11788 22964 13300
rect 23436 13300 23492 13310
rect 23436 13076 23492 13244
rect 23436 13010 23492 13020
rect 22644 11732 22672 11788
rect 22728 11732 22776 11788
rect 22832 11732 22880 11788
rect 22936 11732 22964 11788
rect 22644 10220 22964 11732
rect 29797 12572 30117 14084
rect 32172 20692 32228 20702
rect 32172 14084 32228 20636
rect 34748 16436 34804 27580
rect 36951 27468 37271 28980
rect 36951 27412 36979 27468
rect 37035 27412 37083 27468
rect 37139 27412 37187 27468
rect 37243 27412 37271 27468
rect 36951 25900 37271 27412
rect 44104 31388 44424 32900
rect 44104 31332 44132 31388
rect 44188 31332 44236 31388
rect 44292 31332 44340 31388
rect 44396 31332 44424 31388
rect 44104 29820 44424 31332
rect 44104 29764 44132 29820
rect 44188 29764 44236 29820
rect 44292 29764 44340 29820
rect 44396 29764 44424 29820
rect 44104 28252 44424 29764
rect 44104 28196 44132 28252
rect 44188 28196 44236 28252
rect 44292 28196 44340 28252
rect 44396 28196 44424 28252
rect 44104 26684 44424 28196
rect 44104 26628 44132 26684
rect 44188 26628 44236 26684
rect 44292 26628 44340 26684
rect 44396 26628 44424 26684
rect 37996 26292 38052 26302
rect 36951 25844 36979 25900
rect 37035 25844 37083 25900
rect 37139 25844 37187 25900
rect 37243 25844 37271 25900
rect 36951 24332 37271 25844
rect 37884 25956 37940 25966
rect 36951 24276 36979 24332
rect 37035 24276 37083 24332
rect 37139 24276 37187 24332
rect 37243 24276 37271 24332
rect 36951 22764 37271 24276
rect 37548 25396 37604 25406
rect 37548 24612 37604 25340
rect 37884 24836 37940 25900
rect 37884 24770 37940 24780
rect 37548 23716 37604 24556
rect 37548 23650 37604 23660
rect 37996 23716 38052 26236
rect 38220 25956 38276 25966
rect 38108 25732 38164 25742
rect 38108 24612 38164 25676
rect 38108 24546 38164 24556
rect 38220 24388 38276 25900
rect 38332 25844 38388 25854
rect 38332 25396 38388 25788
rect 38332 25330 38388 25340
rect 38220 24322 38276 24332
rect 44104 25116 44424 26628
rect 51258 36876 51578 36908
rect 51258 36820 51286 36876
rect 51342 36820 51390 36876
rect 51446 36820 51494 36876
rect 51550 36820 51578 36876
rect 51258 35308 51578 36820
rect 51258 35252 51286 35308
rect 51342 35252 51390 35308
rect 51446 35252 51494 35308
rect 51550 35252 51578 35308
rect 51258 33740 51578 35252
rect 51258 33684 51286 33740
rect 51342 33684 51390 33740
rect 51446 33684 51494 33740
rect 51550 33684 51578 33740
rect 51258 32172 51578 33684
rect 51258 32116 51286 32172
rect 51342 32116 51390 32172
rect 51446 32116 51494 32172
rect 51550 32116 51578 32172
rect 51258 30604 51578 32116
rect 58411 36092 58731 36908
rect 58411 36036 58439 36092
rect 58495 36036 58543 36092
rect 58599 36036 58647 36092
rect 58703 36036 58731 36092
rect 58411 34524 58731 36036
rect 58411 34468 58439 34524
rect 58495 34468 58543 34524
rect 58599 34468 58647 34524
rect 58703 34468 58731 34524
rect 58411 32956 58731 34468
rect 58411 32900 58439 32956
rect 58495 32900 58543 32956
rect 58599 32900 58647 32956
rect 58703 32900 58731 32956
rect 51258 30548 51286 30604
rect 51342 30548 51390 30604
rect 51446 30548 51494 30604
rect 51550 30548 51578 30604
rect 51258 29036 51578 30548
rect 51258 28980 51286 29036
rect 51342 28980 51390 29036
rect 51446 28980 51494 29036
rect 51550 28980 51578 29036
rect 51258 27468 51578 28980
rect 51258 27412 51286 27468
rect 51342 27412 51390 27468
rect 51446 27412 51494 27468
rect 51550 27412 51578 27468
rect 44104 25060 44132 25116
rect 44188 25060 44236 25116
rect 44292 25060 44340 25116
rect 44396 25060 44424 25116
rect 37996 23650 38052 23660
rect 36951 22708 36979 22764
rect 37035 22708 37083 22764
rect 37139 22708 37187 22764
rect 37243 22708 37271 22764
rect 44104 23548 44424 25060
rect 44492 26404 44548 26414
rect 44492 24724 44548 26348
rect 44492 24658 44548 24668
rect 51258 25900 51578 27412
rect 51258 25844 51286 25900
rect 51342 25844 51390 25900
rect 51446 25844 51494 25900
rect 51550 25844 51578 25900
rect 44104 23492 44132 23548
rect 44188 23492 44236 23548
rect 44292 23492 44340 23548
rect 44396 23492 44424 23548
rect 36951 21196 37271 22708
rect 36951 21140 36979 21196
rect 37035 21140 37083 21196
rect 37139 21140 37187 21196
rect 37243 21140 37271 21196
rect 36951 19628 37271 21140
rect 37996 22708 38052 22718
rect 37996 21140 38052 22652
rect 37996 21074 38052 21084
rect 44104 21980 44424 23492
rect 44716 24388 44772 24398
rect 44716 23492 44772 24332
rect 51258 24332 51578 25844
rect 56924 31780 56980 31790
rect 56924 31108 56980 31724
rect 56924 24500 56980 31052
rect 56924 24434 56980 24444
rect 58411 31388 58731 32900
rect 58411 31332 58439 31388
rect 58495 31332 58543 31388
rect 58599 31332 58647 31388
rect 58703 31332 58731 31388
rect 58411 29820 58731 31332
rect 58411 29764 58439 29820
rect 58495 29764 58543 29820
rect 58599 29764 58647 29820
rect 58703 29764 58731 29820
rect 58411 28252 58731 29764
rect 58411 28196 58439 28252
rect 58495 28196 58543 28252
rect 58599 28196 58647 28252
rect 58703 28196 58731 28252
rect 58411 26684 58731 28196
rect 58411 26628 58439 26684
rect 58495 26628 58543 26684
rect 58599 26628 58647 26684
rect 58703 26628 58731 26684
rect 58411 25116 58731 26628
rect 58411 25060 58439 25116
rect 58495 25060 58543 25116
rect 58599 25060 58647 25116
rect 58703 25060 58731 25116
rect 51258 24276 51286 24332
rect 51342 24276 51390 24332
rect 51446 24276 51494 24332
rect 51550 24276 51578 24332
rect 50540 23716 50596 23726
rect 44716 23426 44772 23436
rect 45276 23492 45332 23502
rect 45276 23156 45332 23436
rect 45276 23090 45332 23100
rect 44104 21924 44132 21980
rect 44188 21924 44236 21980
rect 44292 21924 44340 21980
rect 44396 21924 44424 21980
rect 36951 19572 36979 19628
rect 37035 19572 37083 19628
rect 37139 19572 37187 19628
rect 37243 19572 37271 19628
rect 35644 19124 35700 19134
rect 35644 17556 35700 19068
rect 35644 17490 35700 17500
rect 36428 18900 36484 18910
rect 36428 16772 36484 18844
rect 36428 16706 36484 16716
rect 36764 18676 36820 18686
rect 36764 16772 36820 18620
rect 36764 16706 36820 16716
rect 36951 18060 37271 19572
rect 44104 20412 44424 21924
rect 44104 20356 44132 20412
rect 44188 20356 44236 20412
rect 44292 20356 44340 20412
rect 44396 20356 44424 20412
rect 44104 18844 44424 20356
rect 46060 22260 46116 22270
rect 46060 19908 46116 22204
rect 46060 19842 46116 19852
rect 47068 21588 47124 21598
rect 44104 18788 44132 18844
rect 44188 18788 44236 18844
rect 44292 18788 44340 18844
rect 44396 18788 44424 18844
rect 36951 18004 36979 18060
rect 37035 18004 37083 18060
rect 37139 18004 37187 18060
rect 37243 18004 37271 18060
rect 34748 15428 34804 16380
rect 34748 15362 34804 15372
rect 36951 16492 37271 18004
rect 42924 18340 42980 18350
rect 36951 16436 36979 16492
rect 37035 16436 37083 16492
rect 37139 16436 37187 16492
rect 37243 16436 37271 16492
rect 32172 14018 32228 14028
rect 36951 14924 37271 16436
rect 36951 14868 36979 14924
rect 37035 14868 37083 14924
rect 37139 14868 37187 14924
rect 37243 14868 37271 14924
rect 29797 12516 29825 12572
rect 29881 12516 29929 12572
rect 29985 12516 30033 12572
rect 30089 12516 30117 12572
rect 26684 11508 26740 11518
rect 27020 11508 27076 11518
rect 26740 11452 27020 11458
rect 26684 11402 27076 11452
rect 29797 11004 30117 12516
rect 36951 13356 37271 14868
rect 42812 16884 42868 16894
rect 42812 14196 42868 16828
rect 42812 14130 42868 14140
rect 42924 13860 42980 18284
rect 42924 13794 42980 13804
rect 44104 17276 44424 18788
rect 44104 17220 44132 17276
rect 44188 17220 44236 17276
rect 44292 17220 44340 17276
rect 44396 17220 44424 17276
rect 44104 15708 44424 17220
rect 44104 15652 44132 15708
rect 44188 15652 44236 15708
rect 44292 15652 44340 15708
rect 44396 15652 44424 15708
rect 44104 14140 44424 15652
rect 45164 18004 45220 18014
rect 45164 15652 45220 17948
rect 47068 18004 47124 21532
rect 48300 21588 48356 21598
rect 47068 17938 47124 17948
rect 47516 18004 47572 18014
rect 47516 15876 47572 17948
rect 47516 15810 47572 15820
rect 45164 15586 45220 15596
rect 44104 14084 44132 14140
rect 44188 14084 44236 14140
rect 44292 14084 44340 14140
rect 44396 14084 44424 14140
rect 48300 14196 48356 21532
rect 49084 20916 49140 20926
rect 49084 18900 49140 20860
rect 50540 19684 50596 23660
rect 50540 19618 50596 19628
rect 51258 22764 51578 24276
rect 51258 22708 51286 22764
rect 51342 22708 51390 22764
rect 51446 22708 51494 22764
rect 51550 22708 51578 22764
rect 51258 21196 51578 22708
rect 51258 21140 51286 21196
rect 51342 21140 51390 21196
rect 51446 21140 51494 21196
rect 51550 21140 51578 21196
rect 51258 19628 51578 21140
rect 49084 18834 49140 18844
rect 51258 19572 51286 19628
rect 51342 19572 51390 19628
rect 51446 19572 51494 19628
rect 51550 19572 51578 19628
rect 51258 18060 51578 19572
rect 51258 18004 51286 18060
rect 51342 18004 51390 18060
rect 51446 18004 51494 18060
rect 51550 18004 51578 18060
rect 48748 16660 49252 16678
rect 48804 16622 49196 16660
rect 48748 16594 48804 16604
rect 49196 16594 49252 16604
rect 48300 14130 48356 14140
rect 51258 16492 51578 18004
rect 51258 16436 51286 16492
rect 51342 16436 51390 16492
rect 51446 16436 51494 16492
rect 51550 16436 51578 16492
rect 51258 14924 51578 16436
rect 51258 14868 51286 14924
rect 51342 14868 51390 14924
rect 51446 14868 51494 14924
rect 51550 14868 51578 14924
rect 36951 13300 36979 13356
rect 37035 13300 37083 13356
rect 37139 13300 37187 13356
rect 37243 13300 37271 13356
rect 36951 11788 37271 13300
rect 29797 10948 29825 11004
rect 29881 10948 29929 11004
rect 29985 10948 30033 11004
rect 30089 10948 30117 11004
rect 34300 11732 34356 11742
rect 34300 11172 34356 11676
rect 36951 11732 36979 11788
rect 37035 11732 37083 11788
rect 37139 11732 37187 11788
rect 37243 11732 37271 11788
rect 22644 10164 22672 10220
rect 22728 10164 22776 10220
rect 22832 10164 22880 10220
rect 22936 10164 22964 10220
rect 22644 8652 22964 10164
rect 22644 8596 22672 8652
rect 22728 8596 22776 8652
rect 22832 8596 22880 8652
rect 22936 8596 22964 8652
rect 22644 7084 22964 8596
rect 23100 10724 23156 10734
rect 23100 8372 23156 10668
rect 26852 9604 26908 9614
rect 26852 9478 26908 9548
rect 26852 9422 26964 9478
rect 26908 9044 26964 9422
rect 26908 8978 26964 8988
rect 29797 9436 30117 10948
rect 30268 10948 30324 10958
rect 30268 10388 30324 10892
rect 30268 10322 30324 10332
rect 29797 9380 29825 9436
rect 29881 9380 29929 9436
rect 29985 9380 30033 9436
rect 30089 9380 30117 9436
rect 23100 8306 23156 8316
rect 22644 7028 22672 7084
rect 22728 7028 22776 7084
rect 22832 7028 22880 7084
rect 22936 7028 22964 7084
rect 22644 5516 22964 7028
rect 22644 5460 22672 5516
rect 22728 5460 22776 5516
rect 22832 5460 22880 5516
rect 22936 5460 22964 5516
rect 22644 3948 22964 5460
rect 29797 7868 30117 9380
rect 29797 7812 29825 7868
rect 29881 7812 29929 7868
rect 29985 7812 30033 7868
rect 30089 7812 30117 7868
rect 29797 6300 30117 7812
rect 29797 6244 29825 6300
rect 29881 6244 29929 6300
rect 29985 6244 30033 6300
rect 30089 6244 30117 6300
rect 25676 4900 25732 4910
rect 25676 4798 25732 4844
rect 25340 4742 25732 4798
rect 25340 4452 25396 4742
rect 25340 4386 25396 4396
rect 29797 4732 30117 6244
rect 34300 5908 34356 11116
rect 35308 11172 35364 11182
rect 34524 10612 34580 10622
rect 34524 7812 34580 10556
rect 34636 10500 34692 10510
rect 34636 8932 34692 10444
rect 35308 10052 35364 11116
rect 35308 9986 35364 9996
rect 36951 10220 37271 11732
rect 44104 12572 44424 14084
rect 51258 13356 51578 14868
rect 51258 13300 51286 13356
rect 51342 13300 51390 13356
rect 51446 13300 51494 13356
rect 51550 13300 51578 13356
rect 44104 12516 44132 12572
rect 44188 12516 44236 12572
rect 44292 12516 44340 12572
rect 44396 12516 44424 12572
rect 44104 11004 44424 12516
rect 46060 12964 46116 12974
rect 46060 11844 46116 12908
rect 46060 11778 46116 11788
rect 51258 11788 51578 13300
rect 44104 10948 44132 11004
rect 44188 10948 44236 11004
rect 44292 10948 44340 11004
rect 44396 10948 44424 11004
rect 36951 10164 36979 10220
rect 37035 10164 37083 10220
rect 37139 10164 37187 10220
rect 37243 10164 37271 10220
rect 34636 8866 34692 8876
rect 34524 7746 34580 7756
rect 36951 8652 37271 10164
rect 41244 10500 41300 10510
rect 41244 9044 41300 10444
rect 41244 8978 41300 8988
rect 41468 10500 41524 10510
rect 36951 8596 36979 8652
rect 37035 8596 37083 8652
rect 37139 8596 37187 8652
rect 37243 8596 37271 8652
rect 34300 5842 34356 5852
rect 36951 7084 37271 8596
rect 36951 7028 36979 7084
rect 37035 7028 37083 7084
rect 37139 7028 37187 7084
rect 37243 7028 37271 7084
rect 29797 4676 29825 4732
rect 29881 4676 29929 4732
rect 29985 4676 30033 4732
rect 30089 4676 30117 4732
rect 22644 3892 22672 3948
rect 22728 3892 22776 3948
rect 22832 3892 22880 3948
rect 22936 3892 22964 3948
rect 22644 3076 22964 3892
rect 29797 3164 30117 4676
rect 29797 3108 29825 3164
rect 29881 3108 29929 3164
rect 29985 3108 30033 3164
rect 30089 3108 30117 3164
rect 29797 3076 30117 3108
rect 36951 5516 37271 7028
rect 36951 5460 36979 5516
rect 37035 5460 37083 5516
rect 37139 5460 37187 5516
rect 37243 5460 37271 5516
rect 36951 3948 37271 5460
rect 41468 4340 41524 10444
rect 43036 10276 43092 10286
rect 43036 8820 43092 10220
rect 43036 8754 43092 8764
rect 44104 9436 44424 10948
rect 51258 11732 51286 11788
rect 51342 11732 51390 11788
rect 51446 11732 51494 11788
rect 51550 11732 51578 11788
rect 51258 10220 51578 11732
rect 51258 10164 51286 10220
rect 51342 10164 51390 10220
rect 51446 10164 51494 10220
rect 51550 10164 51578 10220
rect 44104 9380 44132 9436
rect 44188 9380 44236 9436
rect 44292 9380 44340 9436
rect 44396 9380 44424 9436
rect 41468 4274 41524 4284
rect 44104 7868 44424 9380
rect 44104 7812 44132 7868
rect 44188 7812 44236 7868
rect 44292 7812 44340 7868
rect 44396 7812 44424 7868
rect 44104 6300 44424 7812
rect 45948 10052 46004 10062
rect 45948 6804 46004 9996
rect 46060 9268 46116 9278
rect 46060 7924 46116 9212
rect 46060 7858 46116 7868
rect 51258 8652 51578 10164
rect 51258 8596 51286 8652
rect 51342 8596 51390 8652
rect 51446 8596 51494 8652
rect 51550 8596 51578 8652
rect 45948 6738 46004 6748
rect 51258 7084 51578 8596
rect 51258 7028 51286 7084
rect 51342 7028 51390 7084
rect 51446 7028 51494 7084
rect 51550 7028 51578 7084
rect 44104 6244 44132 6300
rect 44188 6244 44236 6300
rect 44292 6244 44340 6300
rect 44396 6244 44424 6300
rect 44104 4732 44424 6244
rect 44104 4676 44132 4732
rect 44188 4676 44236 4732
rect 44292 4676 44340 4732
rect 44396 4676 44424 4732
rect 36951 3892 36979 3948
rect 37035 3892 37083 3948
rect 37139 3892 37187 3948
rect 37243 3892 37271 3948
rect 36951 3076 37271 3892
rect 44104 3164 44424 4676
rect 44104 3108 44132 3164
rect 44188 3108 44236 3164
rect 44292 3108 44340 3164
rect 44396 3108 44424 3164
rect 44104 3076 44424 3108
rect 51258 5516 51578 7028
rect 51258 5460 51286 5516
rect 51342 5460 51390 5516
rect 51446 5460 51494 5516
rect 51550 5460 51578 5516
rect 51258 3948 51578 5460
rect 51258 3892 51286 3948
rect 51342 3892 51390 3948
rect 51446 3892 51494 3948
rect 51550 3892 51578 3948
rect 51258 3076 51578 3892
rect 58411 23548 58731 25060
rect 58411 23492 58439 23548
rect 58495 23492 58543 23548
rect 58599 23492 58647 23548
rect 58703 23492 58731 23548
rect 58411 21980 58731 23492
rect 58411 21924 58439 21980
rect 58495 21924 58543 21980
rect 58599 21924 58647 21980
rect 58703 21924 58731 21980
rect 58411 20412 58731 21924
rect 58411 20356 58439 20412
rect 58495 20356 58543 20412
rect 58599 20356 58647 20412
rect 58703 20356 58731 20412
rect 58411 18844 58731 20356
rect 58411 18788 58439 18844
rect 58495 18788 58543 18844
rect 58599 18788 58647 18844
rect 58703 18788 58731 18844
rect 58411 17276 58731 18788
rect 58411 17220 58439 17276
rect 58495 17220 58543 17276
rect 58599 17220 58647 17276
rect 58703 17220 58731 17276
rect 58411 15708 58731 17220
rect 58411 15652 58439 15708
rect 58495 15652 58543 15708
rect 58599 15652 58647 15708
rect 58703 15652 58731 15708
rect 58411 14140 58731 15652
rect 58411 14084 58439 14140
rect 58495 14084 58543 14140
rect 58599 14084 58647 14140
rect 58703 14084 58731 14140
rect 58411 12572 58731 14084
rect 58411 12516 58439 12572
rect 58495 12516 58543 12572
rect 58599 12516 58647 12572
rect 58703 12516 58731 12572
rect 58411 11004 58731 12516
rect 58411 10948 58439 11004
rect 58495 10948 58543 11004
rect 58599 10948 58647 11004
rect 58703 10948 58731 11004
rect 58411 9436 58731 10948
rect 58411 9380 58439 9436
rect 58495 9380 58543 9436
rect 58599 9380 58647 9436
rect 58703 9380 58731 9436
rect 58411 7868 58731 9380
rect 58411 7812 58439 7868
rect 58495 7812 58543 7868
rect 58599 7812 58647 7868
rect 58703 7812 58731 7868
rect 58411 6300 58731 7812
rect 58411 6244 58439 6300
rect 58495 6244 58543 6300
rect 58599 6244 58647 6300
rect 58703 6244 58731 6300
rect 58411 4732 58731 6244
rect 58411 4676 58439 4732
rect 58495 4676 58543 4732
rect 58599 4676 58647 4732
rect 58703 4676 58731 4732
rect 58411 3164 58731 4676
rect 58411 3108 58439 3164
rect 58495 3108 58543 3164
rect 58599 3108 58647 3164
rect 58703 3108 58731 3164
rect 58411 3076 58731 3108
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1357_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15680 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1358_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1359_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29008 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1360_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1361_
timestamp 1698431365
transform 1 0 30800 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1362_
timestamp 1698431365
transform -1 0 33936 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1363_
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1364_
timestamp 1698431365
transform 1 0 39536 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1365_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6944 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1366_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46704 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1367_
timestamp 1698431365
transform -1 0 8848 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1368_
timestamp 1698431365
transform -1 0 47488 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1369_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8736 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1370_
timestamp 1698431365
transform -1 0 7840 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1371_
timestamp 1698431365
transform 1 0 42336 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1372_
timestamp 1698431365
transform -1 0 9184 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1373_
timestamp 1698431365
transform -1 0 48720 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1374_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42448 0 -1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1375_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22064 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1376_
timestamp 1698431365
transform -1 0 8960 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1377_
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1378_
timestamp 1698431365
transform -1 0 12096 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1379_
timestamp 1698431365
transform 1 0 35616 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1380_
timestamp 1698431365
transform -1 0 8400 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1381_
timestamp 1698431365
transform -1 0 5936 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1382_
timestamp 1698431365
transform -1 0 41664 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1383_
timestamp 1698431365
transform -1 0 8400 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1384_
timestamp 1698431365
transform 1 0 37408 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1385_
timestamp 1698431365
transform -1 0 42336 0 1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1386_
timestamp 1698431365
transform -1 0 20944 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1387_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1388_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20608 0 -1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1389_
timestamp 1698431365
transform -1 0 19712 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1390_
timestamp 1698431365
transform -1 0 5824 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1391_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  _1392_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5264 0 -1 9408
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1393_
timestamp 1698431365
transform -1 0 8512 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1394_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8512 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1395_
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1396_
timestamp 1698431365
transform -1 0 5936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or4_4  _1397_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45472 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or4_4  _1398_
timestamp 1698431365
transform -1 0 40544 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1399_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10528 0 1 14112
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1400_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8400 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1401_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7728 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1402_
timestamp 1698431365
transform -1 0 6944 0 -1 14112
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1403_
timestamp 1698431365
transform -1 0 6048 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1404_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7504 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1405_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7504 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1406_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6048 0 1 9408
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1407_
timestamp 1698431365
transform 1 0 15792 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1408_
timestamp 1698431365
transform 1 0 7504 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1409_
timestamp 1698431365
transform -1 0 20048 0 -1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1410_
timestamp 1698431365
transform 1 0 14560 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1411_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10976 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1412_
timestamp 1698431365
transform -1 0 15008 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1413_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10976 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1414_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1415_
timestamp 1698431365
transform 1 0 22176 0 1 3136
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1416_
timestamp 1698431365
transform 1 0 33152 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1417_
timestamp 1698431365
transform 1 0 34272 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1418_
timestamp 1698431365
transform -1 0 25760 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1419_
timestamp 1698431365
transform 1 0 15008 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1420_
timestamp 1698431365
transform 1 0 21504 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1421_
timestamp 1698431365
transform -1 0 35728 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1422_
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1423_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41664 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1424_
timestamp 1698431365
transform -1 0 48384 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1425_
timestamp 1698431365
transform 1 0 27328 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1426_
timestamp 1698431365
transform 1 0 31248 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1427_
timestamp 1698431365
transform 1 0 41888 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1428_
timestamp 1698431365
transform -1 0 44352 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1429_
timestamp 1698431365
transform 1 0 12432 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1430_
timestamp 1698431365
transform -1 0 30128 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1431_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22176 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1432_
timestamp 1698431365
transform 1 0 22176 0 -1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1433_
timestamp 1698431365
transform 1 0 16240 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1434_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1435_
timestamp 1698431365
transform -1 0 16128 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1436_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18256 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _1437_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20048 0 -1 7840
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1438_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27328 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1439_
timestamp 1698431365
transform 1 0 32928 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1440_
timestamp 1698431365
transform -1 0 32704 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1441_
timestamp 1698431365
transform -1 0 43008 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1442_
timestamp 1698431365
transform -1 0 44240 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1443_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41552 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1444_
timestamp 1698431365
transform 1 0 45808 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1445_
timestamp 1698431365
transform 1 0 43456 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1446_
timestamp 1698431365
transform 1 0 41328 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1447_
timestamp 1698431365
transform 1 0 46256 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1448_
timestamp 1698431365
transform 1 0 44128 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1449_
timestamp 1698431365
transform 1 0 47376 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1450_
timestamp 1698431365
transform 1 0 49280 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1451_
timestamp 1698431365
transform -1 0 48384 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1452_
timestamp 1698431365
transform -1 0 46480 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1453_
timestamp 1698431365
transform -1 0 32704 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1454_
timestamp 1698431365
transform 1 0 46368 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1455_
timestamp 1698431365
transform 1 0 47488 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1456_
timestamp 1698431365
transform -1 0 49280 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1457_
timestamp 1698431365
transform -1 0 46032 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1458_
timestamp 1698431365
transform -1 0 44464 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1459_
timestamp 1698431365
transform 1 0 48608 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1460_
timestamp 1698431365
transform 1 0 48832 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1461_
timestamp 1698431365
transform -1 0 47600 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1462_
timestamp 1698431365
transform -1 0 45584 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1463_
timestamp 1698431365
transform -1 0 44464 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1464_
timestamp 1698431365
transform -1 0 47152 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1465_
timestamp 1698431365
transform -1 0 46480 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1466_
timestamp 1698431365
transform -1 0 45584 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1467_
timestamp 1698431365
transform 1 0 45136 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1468_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46032 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1469_
timestamp 1698431365
transform 1 0 46480 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1470_
timestamp 1698431365
transform 1 0 47152 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1471_
timestamp 1698431365
transform -1 0 44912 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1472_
timestamp 1698431365
transform 1 0 44800 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1473_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46032 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1474_
timestamp 1698431365
transform -1 0 47488 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1475_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45024 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1476_
timestamp 1698431365
transform 1 0 47824 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1477_
timestamp 1698431365
transform 1 0 47600 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1478_
timestamp 1698431365
transform 1 0 23744 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1479_
timestamp 1698431365
transform 1 0 34048 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1480_
timestamp 1698431365
transform 1 0 34160 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1481_
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1482_
timestamp 1698431365
transform -1 0 45136 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1483_
timestamp 1698431365
transform -1 0 41888 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1484_
timestamp 1698431365
transform 1 0 42224 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1485_
timestamp 1698431365
transform -1 0 34384 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1486_
timestamp 1698431365
transform -1 0 15792 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1487_
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1488_
timestamp 1698431365
transform 1 0 17696 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1489_
timestamp 1698431365
transform 1 0 15680 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1490_
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1491_
timestamp 1698431365
transform 1 0 25536 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1492_
timestamp 1698431365
transform 1 0 25872 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1493_
timestamp 1698431365
transform 1 0 25536 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1494_
timestamp 1698431365
transform 1 0 29680 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1495_
timestamp 1698431365
transform -1 0 31136 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1496_
timestamp 1698431365
transform -1 0 33712 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1497_
timestamp 1698431365
transform 1 0 30128 0 -1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1498_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1499_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46368 0 1 4704
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1500_
timestamp 1698431365
transform 1 0 46032 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1501_
timestamp 1698431365
transform 1 0 45920 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1502_
timestamp 1698431365
transform 1 0 46704 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1503_
timestamp 1698431365
transform -1 0 41552 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1504_
timestamp 1698431365
transform -1 0 50960 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1505_
timestamp 1698431365
transform 1 0 48608 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1506_
timestamp 1698431365
transform 1 0 47936 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1507_
timestamp 1698431365
transform -1 0 50064 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1508_
timestamp 1698431365
transform -1 0 50624 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1509_
timestamp 1698431365
transform 1 0 31584 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1510_
timestamp 1698431365
transform 1 0 33488 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1511_
timestamp 1698431365
transform 1 0 46592 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1512_
timestamp 1698431365
transform 1 0 46816 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1513_
timestamp 1698431365
transform 1 0 47712 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1514_
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1515_
timestamp 1698431365
transform 1 0 49056 0 -1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1516_
timestamp 1698431365
transform 1 0 50848 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1517_
timestamp 1698431365
transform -1 0 52192 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1518_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 49168 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1519_
timestamp 1698431365
transform 1 0 47376 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1520_
timestamp 1698431365
transform -1 0 42560 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1521_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42560 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1522_
timestamp 1698431365
transform 1 0 45136 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1523_
timestamp 1698431365
transform 1 0 43008 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1524_
timestamp 1698431365
transform 1 0 43568 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1525_
timestamp 1698431365
transform 1 0 44912 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1526_
timestamp 1698431365
transform 1 0 45472 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1527_
timestamp 1698431365
transform -1 0 46592 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1528_
timestamp 1698431365
transform 1 0 46592 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1529_
timestamp 1698431365
transform -1 0 46704 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1530_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46032 0 1 9408
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1531_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 49392 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1532_
timestamp 1698431365
transform -1 0 50288 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1533_
timestamp 1698431365
transform -1 0 48384 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1534_
timestamp 1698431365
transform 1 0 31920 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1535_
timestamp 1698431365
transform -1 0 34832 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1536_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33600 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1537_
timestamp 1698431365
transform 1 0 33824 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1538_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35392 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1539_
timestamp 1698431365
transform 1 0 30352 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1540_
timestamp 1698431365
transform 1 0 16688 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1541_
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1542_
timestamp 1698431365
transform 1 0 31136 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1543_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31472 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1544_
timestamp 1698431365
transform 1 0 28336 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1545_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32368 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1546_
timestamp 1698431365
transform -1 0 32704 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1547_
timestamp 1698431365
transform -1 0 30128 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1548_
timestamp 1698431365
transform -1 0 33488 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1549_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1550_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1551_
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1552_
timestamp 1698431365
transform -1 0 15680 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1553_
timestamp 1698431365
transform 1 0 14336 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1554_
timestamp 1698431365
transform -1 0 12432 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1555_
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1556_
timestamp 1698431365
transform -1 0 24416 0 -1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1557_
timestamp 1698431365
transform 1 0 18032 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1558_
timestamp 1698431365
transform -1 0 16128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1559_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1560_
timestamp 1698431365
transform -1 0 24752 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1561_
timestamp 1698431365
transform -1 0 8848 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1562_
timestamp 1698431365
transform 1 0 13328 0 -1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1563_
timestamp 1698431365
transform 1 0 21392 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1564_
timestamp 1698431365
transform 1 0 23744 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1565_
timestamp 1698431365
transform 1 0 28112 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1566_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28000 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1567_
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1568_
timestamp 1698431365
transform -1 0 44016 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1569_
timestamp 1698431365
transform 1 0 40656 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1570_
timestamp 1698431365
transform 1 0 41328 0 1 3136
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _1571_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43680 0 -1 4704
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1572_
timestamp 1698431365
transform 1 0 49280 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1573_
timestamp 1698431365
transform 1 0 49392 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1574_
timestamp 1698431365
transform 1 0 49840 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1575_
timestamp 1698431365
transform 1 0 49168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1576_
timestamp 1698431365
transform 1 0 50960 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1577_
timestamp 1698431365
transform 1 0 50736 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1578_
timestamp 1698431365
transform 1 0 48272 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1579_
timestamp 1698431365
transform 1 0 49168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1580_
timestamp 1698431365
transform 1 0 48832 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1581_
timestamp 1698431365
transform 1 0 42896 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1582_
timestamp 1698431365
transform 1 0 23520 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1583_
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1584_
timestamp 1698431365
transform -1 0 40096 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1585_
timestamp 1698431365
transform 1 0 40992 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1586_
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1587_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41552 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1588_
timestamp 1698431365
transform 1 0 43008 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1589_
timestamp 1698431365
transform 1 0 51184 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1590_
timestamp 1698431365
transform 1 0 52640 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1591_
timestamp 1698431365
transform 1 0 51184 0 -1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1592_
timestamp 1698431365
transform 1 0 51408 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1593_
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1594_
timestamp 1698431365
transform -1 0 53648 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1595_
timestamp 1698431365
transform -1 0 50848 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1596_
timestamp 1698431365
transform -1 0 50064 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1597_
timestamp 1698431365
transform -1 0 20944 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1598_
timestamp 1698431365
transform 1 0 53648 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1599_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 49168 0 1 9408
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1600_
timestamp 1698431365
transform 1 0 35392 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1601_
timestamp 1698431365
transform -1 0 35168 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1602_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 50064 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1603_
timestamp 1698431365
transform 1 0 44016 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1604_
timestamp 1698431365
transform 1 0 43344 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1605_
timestamp 1698431365
transform 1 0 44688 0 1 3136
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1606_
timestamp 1698431365
transform 1 0 37408 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1607_
timestamp 1698431365
transform 1 0 39984 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1608_
timestamp 1698431365
transform -1 0 38976 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1609_
timestamp 1698431365
transform 1 0 38080 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1610_
timestamp 1698431365
transform -1 0 36624 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1611_
timestamp 1698431365
transform 1 0 33824 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1612_
timestamp 1698431365
transform 1 0 32144 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1613_
timestamp 1698431365
transform 1 0 34832 0 -1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1614_
timestamp 1698431365
transform -1 0 27664 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1615_
timestamp 1698431365
transform 1 0 29232 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1616_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27216 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1617_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1618_
timestamp 1698431365
transform 1 0 28000 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1619_
timestamp 1698431365
transform 1 0 32368 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1620_
timestamp 1698431365
transform -1 0 36288 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1621_
timestamp 1698431365
transform -1 0 8624 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1622_
timestamp 1698431365
transform 1 0 14448 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1623_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26656 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1624_
timestamp 1698431365
transform 1 0 20720 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1625_
timestamp 1698431365
transform -1 0 23632 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1626_
timestamp 1698431365
transform 1 0 21952 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1627_
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1628_
timestamp 1698431365
transform 1 0 25424 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1629_
timestamp 1698431365
transform -1 0 20496 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1630_
timestamp 1698431365
transform -1 0 24640 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1631_
timestamp 1698431365
transform -1 0 27104 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1632_
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1633_
timestamp 1698431365
transform 1 0 37856 0 1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1634_
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1635_
timestamp 1698431365
transform 1 0 43680 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1636_
timestamp 1698431365
transform 1 0 50624 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1637_
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1638_
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1639_
timestamp 1698431365
transform 1 0 42000 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1640_
timestamp 1698431365
transform 1 0 42784 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1641_
timestamp 1698431365
transform 1 0 43456 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1642_
timestamp 1698431365
transform 1 0 47376 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1643_
timestamp 1698431365
transform 1 0 48608 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1644_
timestamp 1698431365
transform 1 0 46032 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1645_
timestamp 1698431365
transform 1 0 22960 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1646_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21840 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1647_
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1648_
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1649_
timestamp 1698431365
transform 1 0 45472 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1650_
timestamp 1698431365
transform 1 0 52416 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1651_
timestamp 1698431365
transform 1 0 53872 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1652_
timestamp 1698431365
transform -1 0 57904 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1653_
timestamp 1698431365
transform 1 0 50624 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1654_
timestamp 1698431365
transform 1 0 50288 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1655_
timestamp 1698431365
transform 1 0 49728 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1656_
timestamp 1698431365
transform 1 0 54768 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1657_
timestamp 1698431365
transform -1 0 57904 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1658_
timestamp 1698431365
transform -1 0 57568 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1659_
timestamp 1698431365
transform -1 0 55552 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1660_
timestamp 1698431365
transform 1 0 54096 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1661_
timestamp 1698431365
transform 1 0 54656 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1662_
timestamp 1698431365
transform 1 0 54208 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1663_
timestamp 1698431365
transform 1 0 54880 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1664_
timestamp 1698431365
transform -1 0 55776 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1665_
timestamp 1698431365
transform -1 0 56224 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1666_
timestamp 1698431365
transform -1 0 22512 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1667_
timestamp 1698431365
transform -1 0 20272 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1668_
timestamp 1698431365
transform -1 0 14336 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1669_
timestamp 1698431365
transform -1 0 23072 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1670_
timestamp 1698431365
transform 1 0 17696 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1671_
timestamp 1698431365
transform 1 0 19824 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1672_
timestamp 1698431365
transform -1 0 28560 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1673_
timestamp 1698431365
transform 1 0 30352 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1674_
timestamp 1698431365
transform 1 0 55104 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1675_
timestamp 1698431365
transform 1 0 54768 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1676_
timestamp 1698431365
transform 1 0 55216 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1677_
timestamp 1698431365
transform -1 0 57904 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1678_
timestamp 1698431365
transform 1 0 50960 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1679_
timestamp 1698431365
transform 1 0 50848 0 1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1680_
timestamp 1698431365
transform -1 0 56224 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1681_
timestamp 1698431365
transform 1 0 54544 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1682_
timestamp 1698431365
transform 1 0 55104 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1683_
timestamp 1698431365
transform 1 0 54656 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1684_
timestamp 1698431365
transform -1 0 56112 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1685_
timestamp 1698431365
transform 1 0 55328 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1686_
timestamp 1698431365
transform 1 0 45920 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1687_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1688_
timestamp 1698431365
transform -1 0 43904 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1689_
timestamp 1698431365
transform 1 0 40880 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1690_
timestamp 1698431365
transform -1 0 38528 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1691_
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1692_
timestamp 1698431365
transform 1 0 40880 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1693_
timestamp 1698431365
transform 1 0 34720 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1694_
timestamp 1698431365
transform 1 0 35616 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1695_
timestamp 1698431365
transform 1 0 35168 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1696_
timestamp 1698431365
transform -1 0 33488 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1697_
timestamp 1698431365
transform 1 0 39088 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1698_
timestamp 1698431365
transform 1 0 39536 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1699_
timestamp 1698431365
transform -1 0 38976 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1700_
timestamp 1698431365
transform 1 0 40544 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1701_
timestamp 1698431365
transform -1 0 40432 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1702_
timestamp 1698431365
transform 1 0 35616 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1703_
timestamp 1698431365
transform 1 0 31808 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1704_
timestamp 1698431365
transform 1 0 22288 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1705_
timestamp 1698431365
transform 1 0 22848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1706_
timestamp 1698431365
transform -1 0 33376 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1707_
timestamp 1698431365
transform 1 0 30912 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1708_
timestamp 1698431365
transform -1 0 35616 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1709_
timestamp 1698431365
transform 1 0 34496 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1710_
timestamp 1698431365
transform 1 0 35616 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1711_
timestamp 1698431365
transform -1 0 39088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1712_
timestamp 1698431365
transform -1 0 38192 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1713_
timestamp 1698431365
transform 1 0 25872 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1714_
timestamp 1698431365
transform 1 0 27664 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1715_
timestamp 1698431365
transform 1 0 24976 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1716_
timestamp 1698431365
transform 1 0 29344 0 -1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1717_
timestamp 1698431365
transform 1 0 31808 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1718_
timestamp 1698431365
transform 1 0 32256 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1719_
timestamp 1698431365
transform 1 0 32816 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1720_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1721_
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1722_
timestamp 1698431365
transform 1 0 44576 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1723_
timestamp 1698431365
transform 1 0 41552 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1724_
timestamp 1698431365
transform 1 0 54320 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1725_
timestamp 1698431365
transform 1 0 55552 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1726_
timestamp 1698431365
transform 1 0 56560 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1727_
timestamp 1698431365
transform 1 0 57568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1728_
timestamp 1698431365
transform 1 0 54544 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1729_
timestamp 1698431365
transform -1 0 54544 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1730_
timestamp 1698431365
transform 1 0 45360 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1731_
timestamp 1698431365
transform -1 0 45360 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1732_
timestamp 1698431365
transform -1 0 45584 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1733_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45696 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1734_
timestamp 1698431365
transform 1 0 45696 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1735_
timestamp 1698431365
transform -1 0 45360 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1736_
timestamp 1698431365
transform -1 0 40320 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1737_
timestamp 1698431365
transform 1 0 45584 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1738_
timestamp 1698431365
transform 1 0 45472 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1739_
timestamp 1698431365
transform 1 0 49952 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1740_
timestamp 1698431365
transform 1 0 47600 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1741_
timestamp 1698431365
transform 1 0 50288 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1742_
timestamp 1698431365
transform 1 0 48832 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1743_
timestamp 1698431365
transform 1 0 49616 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1744_
timestamp 1698431365
transform -1 0 51744 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1745_
timestamp 1698431365
transform -1 0 53088 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1746_
timestamp 1698431365
transform 1 0 50288 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1747_
timestamp 1698431365
transform 1 0 50848 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1748_
timestamp 1698431365
transform 1 0 52976 0 -1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1749_
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1750_
timestamp 1698431365
transform 1 0 55776 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1751_
timestamp 1698431365
transform 1 0 55776 0 1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _1752_
timestamp 1698431365
transform -1 0 58352 0 1 12544
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1753_
timestamp 1698431365
transform -1 0 19824 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1754_
timestamp 1698431365
transform -1 0 19152 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1755_
timestamp 1698431365
transform -1 0 12656 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1756_
timestamp 1698431365
transform 1 0 19712 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1757_
timestamp 1698431365
transform -1 0 20608 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1758_
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1759_
timestamp 1698431365
transform 1 0 57120 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1760_
timestamp 1698431365
transform -1 0 58128 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1761_
timestamp 1698431365
transform -1 0 54320 0 -1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1762_
timestamp 1698431365
transform -1 0 58352 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1763_
timestamp 1698431365
transform -1 0 57568 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1764_
timestamp 1698431365
transform -1 0 56224 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1765_
timestamp 1698431365
transform -1 0 57904 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1766_
timestamp 1698431365
transform 1 0 55664 0 1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1767_
timestamp 1698431365
transform -1 0 57904 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1768_
timestamp 1698431365
transform 1 0 55552 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1769_
timestamp 1698431365
transform 1 0 54880 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1770_
timestamp 1698431365
transform 1 0 53872 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1771_
timestamp 1698431365
transform 1 0 53200 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1772_
timestamp 1698431365
transform 1 0 52976 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1773_
timestamp 1698431365
transform 1 0 46816 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1774_
timestamp 1698431365
transform 1 0 43792 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1775_
timestamp 1698431365
transform 1 0 44352 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1776_
timestamp 1698431365
transform -1 0 44800 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1777_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1778_
timestamp 1698431365
transform -1 0 38304 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1779_
timestamp 1698431365
transform 1 0 38976 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1780_
timestamp 1698431365
transform 1 0 38080 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1781_
timestamp 1698431365
transform -1 0 38416 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1782_
timestamp 1698431365
transform 1 0 42448 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1783_
timestamp 1698431365
transform 1 0 38080 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1784_
timestamp 1698431365
transform 1 0 39200 0 1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1785_
timestamp 1698431365
transform 1 0 44240 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1786_
timestamp 1698431365
transform 1 0 53760 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1787_
timestamp 1698431365
transform -1 0 54768 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1788_
timestamp 1698431365
transform -1 0 52752 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1789_
timestamp 1698431365
transform -1 0 52752 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1790_
timestamp 1698431365
transform 1 0 41440 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1791_
timestamp 1698431365
transform -1 0 44576 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1792_
timestamp 1698431365
transform 1 0 41216 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _1793_
timestamp 1698431365
transform 1 0 42560 0 -1 20384
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1794_
timestamp 1698431365
transform 1 0 43568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1795_
timestamp 1698431365
transform 1 0 38416 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1796_
timestamp 1698431365
transform 1 0 39648 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1797_
timestamp 1698431365
transform 1 0 39088 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1798_
timestamp 1698431365
transform -1 0 41440 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1799_
timestamp 1698431365
transform 1 0 39648 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1800_
timestamp 1698431365
transform -1 0 34496 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1801_
timestamp 1698431365
transform 1 0 33488 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1802_
timestamp 1698431365
transform 1 0 34048 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1803_
timestamp 1698431365
transform -1 0 35168 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1804_
timestamp 1698431365
transform 1 0 35168 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1805_
timestamp 1698431365
transform 1 0 36176 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1806_
timestamp 1698431365
transform -1 0 37408 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1807_
timestamp 1698431365
transform -1 0 36624 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1808_
timestamp 1698431365
transform 1 0 21168 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1809_
timestamp 1698431365
transform -1 0 31808 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1810_
timestamp 1698431365
transform 1 0 32816 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1811_
timestamp 1698431365
transform -1 0 33600 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1812_
timestamp 1698431365
transform -1 0 34160 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1813_
timestamp 1698431365
transform 1 0 31920 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1814_
timestamp 1698431365
transform 1 0 26768 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1815_
timestamp 1698431365
transform 1 0 29344 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1816_
timestamp 1698431365
transform -1 0 32256 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1817_
timestamp 1698431365
transform 1 0 29120 0 1 9408
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1818_
timestamp 1698431365
transform -1 0 31360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1819_
timestamp 1698431365
transform 1 0 26880 0 1 9408
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1820_
timestamp 1698431365
transform 1 0 26768 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1821_
timestamp 1698431365
transform -1 0 31808 0 -1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1822_
timestamp 1698431365
transform 1 0 34496 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1823_
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1824_
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1825_
timestamp 1698431365
transform 1 0 42112 0 -1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1826_
timestamp 1698431365
transform -1 0 45808 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1827_
timestamp 1698431365
transform -1 0 45248 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1828_
timestamp 1698431365
transform 1 0 44576 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1829_
timestamp 1698431365
transform 1 0 45472 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1830_
timestamp 1698431365
transform 1 0 50848 0 -1 34496
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1831_
timestamp 1698431365
transform 1 0 53760 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1832_
timestamp 1698431365
transform -1 0 58016 0 1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1833_
timestamp 1698431365
transform -1 0 57792 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1834_
timestamp 1698431365
transform 1 0 19152 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1835_
timestamp 1698431365
transform -1 0 20160 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1836_
timestamp 1698431365
transform -1 0 10416 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1837_
timestamp 1698431365
transform -1 0 21728 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1838_
timestamp 1698431365
transform 1 0 20160 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1839_
timestamp 1698431365
transform -1 0 34272 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1840_
timestamp 1698431365
transform 1 0 56336 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1841_
timestamp 1698431365
transform 1 0 55664 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1842_
timestamp 1698431365
transform -1 0 58352 0 1 32928
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1843_
timestamp 1698431365
transform 1 0 53536 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1844_
timestamp 1698431365
transform -1 0 57008 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1845_
timestamp 1698431365
transform 1 0 54432 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1846_
timestamp 1698431365
transform 1 0 50288 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1847_
timestamp 1698431365
transform -1 0 51520 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1848_
timestamp 1698431365
transform -1 0 50848 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1849_
timestamp 1698431365
transform 1 0 51184 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1850_
timestamp 1698431365
transform -1 0 54320 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1851_
timestamp 1698431365
transform 1 0 52864 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1852_
timestamp 1698431365
transform -1 0 40544 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1853_
timestamp 1698431365
transform -1 0 44240 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1854_
timestamp 1698431365
transform -1 0 44464 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1855_
timestamp 1698431365
transform -1 0 41664 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1856_
timestamp 1698431365
transform -1 0 14560 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1857_
timestamp 1698431365
transform -1 0 31024 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1858_
timestamp 1698431365
transform 1 0 34048 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1859_
timestamp 1698431365
transform -1 0 38080 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1860_
timestamp 1698431365
transform -1 0 38080 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1861_
timestamp 1698431365
transform 1 0 35168 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1862_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1863_
timestamp 1698431365
transform 1 0 39424 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1864_
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1865_
timestamp 1698431365
transform 1 0 46032 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1866_
timestamp 1698431365
transform -1 0 44576 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1867_
timestamp 1698431365
transform 1 0 42672 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1868_
timestamp 1698431365
transform -1 0 44464 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1869_
timestamp 1698431365
transform 1 0 43456 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1870_
timestamp 1698431365
transform -1 0 41328 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform -1 0 40544 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1872_
timestamp 1698431365
transform -1 0 40320 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1873_
timestamp 1698431365
transform -1 0 42224 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1874_
timestamp 1698431365
transform -1 0 44688 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1875_
timestamp 1698431365
transform -1 0 41776 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1876_
timestamp 1698431365
transform -1 0 44464 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1877_
timestamp 1698431365
transform 1 0 39648 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1878_
timestamp 1698431365
transform 1 0 40992 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1879_
timestamp 1698431365
transform -1 0 42336 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1880_
timestamp 1698431365
transform 1 0 34048 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1881_
timestamp 1698431365
transform -1 0 35280 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1882_
timestamp 1698431365
transform -1 0 36512 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1883_
timestamp 1698431365
transform -1 0 35728 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1884_
timestamp 1698431365
transform 1 0 35840 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1885_
timestamp 1698431365
transform -1 0 38080 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1886_
timestamp 1698431365
transform -1 0 37744 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1887_
timestamp 1698431365
transform -1 0 31360 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1888_
timestamp 1698431365
transform -1 0 26768 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1889_
timestamp 1698431365
transform -1 0 28672 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1890_
timestamp 1698431365
transform 1 0 26320 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1891_
timestamp 1698431365
transform -1 0 30464 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1892_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18928 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1893_
timestamp 1698431365
transform 1 0 30128 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1894_
timestamp 1698431365
transform -1 0 25760 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1895_
timestamp 1698431365
transform -1 0 30464 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1896_
timestamp 1698431365
transform -1 0 30352 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1897_
timestamp 1698431365
transform 1 0 29120 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1898_
timestamp 1698431365
transform 1 0 30128 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1899_
timestamp 1698431365
transform -1 0 32704 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1900_
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1901_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1902_
timestamp 1698431365
transform -1 0 34160 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1903_
timestamp 1698431365
transform -1 0 33488 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1904_
timestamp 1698431365
transform -1 0 35168 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1905_
timestamp 1698431365
transform -1 0 32704 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1906_
timestamp 1698431365
transform 1 0 30800 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1907_
timestamp 1698431365
transform 1 0 33600 0 -1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1908_
timestamp 1698431365
transform 1 0 36176 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1909_
timestamp 1698431365
transform -1 0 37408 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1910_
timestamp 1698431365
transform -1 0 37296 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1911_
timestamp 1698431365
transform -1 0 36512 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1912_
timestamp 1698431365
transform 1 0 35840 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1913_
timestamp 1698431365
transform 1 0 38304 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1914_
timestamp 1698431365
transform 1 0 40992 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1915_
timestamp 1698431365
transform 1 0 46480 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1916_
timestamp 1698431365
transform 1 0 50064 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1917_
timestamp 1698431365
transform -1 0 53424 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1918_
timestamp 1698431365
transform -1 0 51184 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1919_
timestamp 1698431365
transform -1 0 20832 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1920_
timestamp 1698431365
transform -1 0 8400 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1921_
timestamp 1698431365
transform 1 0 48720 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1922_
timestamp 1698431365
transform 1 0 51408 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1923_
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1924_
timestamp 1698431365
transform 1 0 21840 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1925_
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1926_
timestamp 1698431365
transform 1 0 51632 0 -1 36064
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1927_
timestamp 1698431365
transform 1 0 46592 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1928_
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1929_
timestamp 1698431365
transform -1 0 50288 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1930_
timestamp 1698431365
transform -1 0 49728 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1931_
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1932_
timestamp 1698431365
transform -1 0 42224 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1933_
timestamp 1698431365
transform -1 0 41664 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1934_
timestamp 1698431365
transform 1 0 40208 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1935_
timestamp 1698431365
transform 1 0 40880 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1936_
timestamp 1698431365
transform -1 0 45248 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1937_
timestamp 1698431365
transform 1 0 43568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1938_
timestamp 1698431365
transform -1 0 39424 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1939_
timestamp 1698431365
transform -1 0 36848 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1940_
timestamp 1698431365
transform 1 0 38528 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1941_
timestamp 1698431365
transform -1 0 35056 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1942_
timestamp 1698431365
transform 1 0 33712 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1943_
timestamp 1698431365
transform 1 0 33600 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1944_
timestamp 1698431365
transform 1 0 30688 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1945_
timestamp 1698431365
transform 1 0 32256 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1946_
timestamp 1698431365
transform -1 0 34832 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1947_
timestamp 1698431365
transform -1 0 37520 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1948_
timestamp 1698431365
transform 1 0 22624 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1949_
timestamp 1698431365
transform -1 0 34048 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1950_
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1951_
timestamp 1698431365
transform 1 0 35280 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1952_
timestamp 1698431365
transform -1 0 38304 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1953_
timestamp 1698431365
transform -1 0 38528 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1954_
timestamp 1698431365
transform -1 0 35840 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1955_
timestamp 1698431365
transform -1 0 37744 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1956_
timestamp 1698431365
transform -1 0 37520 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1957_
timestamp 1698431365
transform -1 0 36624 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1958_
timestamp 1698431365
transform -1 0 36624 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1959_
timestamp 1698431365
transform 1 0 35504 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1960_
timestamp 1698431365
transform 1 0 36624 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1961_
timestamp 1698431365
transform -1 0 39872 0 1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1962_
timestamp 1698431365
transform -1 0 33376 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1963_
timestamp 1698431365
transform -1 0 32704 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1964_
timestamp 1698431365
transform -1 0 34832 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1965_
timestamp 1698431365
transform -1 0 33936 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1966_
timestamp 1698431365
transform -1 0 33600 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1967_
timestamp 1698431365
transform -1 0 34608 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1968_
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1969_
timestamp 1698431365
transform 1 0 29568 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1970_
timestamp 1698431365
transform 1 0 30800 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1971_
timestamp 1698431365
transform -1 0 31808 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1972_
timestamp 1698431365
transform 1 0 27776 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1973_
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1974_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1975_
timestamp 1698431365
transform -1 0 23856 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1976_
timestamp 1698431365
transform -1 0 24752 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1977_
timestamp 1698431365
transform -1 0 27216 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1978_
timestamp 1698431365
transform 1 0 23744 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1979_
timestamp 1698431365
transform 1 0 25760 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1980_
timestamp 1698431365
transform -1 0 28112 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1981_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1982_
timestamp 1698431365
transform 1 0 30352 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1983_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1984_
timestamp 1698431365
transform -1 0 32816 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1985_
timestamp 1698431365
transform -1 0 30240 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1986_
timestamp 1698431365
transform -1 0 30800 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1987_
timestamp 1698431365
transform -1 0 30464 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1988_
timestamp 1698431365
transform 1 0 26880 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1989_
timestamp 1698431365
transform 1 0 27440 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1990_
timestamp 1698431365
transform 1 0 27440 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1991_
timestamp 1698431365
transform -1 0 29792 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1992_
timestamp 1698431365
transform 1 0 13328 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1993_
timestamp 1698431365
transform -1 0 22288 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1994_
timestamp 1698431365
transform 1 0 14000 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1995_
timestamp 1698431365
transform -1 0 25760 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1996_
timestamp 1698431365
transform 1 0 22064 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1997_
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1998_
timestamp 1698431365
transform 1 0 27216 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _1999_
timestamp 1698431365
transform 1 0 35840 0 -1 31360
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2000_
timestamp 1698431365
transform 1 0 37184 0 -1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2001_
timestamp 1698431365
transform -1 0 42112 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2002_
timestamp 1698431365
transform -1 0 36512 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2003_
timestamp 1698431365
transform -1 0 25872 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2004_
timestamp 1698431365
transform 1 0 21392 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2005_
timestamp 1698431365
transform -1 0 23072 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2006_
timestamp 1698431365
transform -1 0 21952 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2007_
timestamp 1698431365
transform 1 0 23408 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2008_
timestamp 1698431365
transform 1 0 25872 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2009_
timestamp 1698431365
transform -1 0 26096 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2010_
timestamp 1698431365
transform -1 0 37520 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2011_
timestamp 1698431365
transform -1 0 37072 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2012_
timestamp 1698431365
transform 1 0 33600 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2013_
timestamp 1698431365
transform -1 0 40208 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2014_
timestamp 1698431365
transform -1 0 38080 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2015_
timestamp 1698431365
transform -1 0 40320 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2016_
timestamp 1698431365
transform -1 0 35728 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2017_
timestamp 1698431365
transform 1 0 26320 0 1 28224
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2018_
timestamp 1698431365
transform 1 0 27440 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2019_
timestamp 1698431365
transform 1 0 31248 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2020_
timestamp 1698431365
transform 1 0 31136 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2021_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2022_
timestamp 1698431365
transform -1 0 32928 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2023_
timestamp 1698431365
transform -1 0 39648 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2024_
timestamp 1698431365
transform -1 0 38528 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2025_
timestamp 1698431365
transform -1 0 26096 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2026_
timestamp 1698431365
transform 1 0 24752 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2027_
timestamp 1698431365
transform -1 0 24752 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2028_
timestamp 1698431365
transform -1 0 33600 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2029_
timestamp 1698431365
transform -1 0 25984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2030_
timestamp 1698431365
transform 1 0 29792 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2031_
timestamp 1698431365
transform -1 0 28784 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2032_
timestamp 1698431365
transform -1 0 31696 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2033_
timestamp 1698431365
transform -1 0 30800 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2034_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2035_
timestamp 1698431365
transform 1 0 30464 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2036_
timestamp 1698431365
transform 1 0 29008 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2037_
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2038_
timestamp 1698431365
transform -1 0 28560 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2039_
timestamp 1698431365
transform 1 0 25872 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2040_
timestamp 1698431365
transform 1 0 27104 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2041_
timestamp 1698431365
transform -1 0 23744 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2042_
timestamp 1698431365
transform 1 0 22736 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2043_
timestamp 1698431365
transform -1 0 22512 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2044_
timestamp 1698431365
transform -1 0 21952 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2045_
timestamp 1698431365
transform 1 0 28336 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2046_
timestamp 1698431365
transform 1 0 25088 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2047_
timestamp 1698431365
transform -1 0 32256 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2048_
timestamp 1698431365
transform -1 0 25872 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2049_
timestamp 1698431365
transform -1 0 25648 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2050_
timestamp 1698431365
transform -1 0 26544 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2051_
timestamp 1698431365
transform -1 0 23856 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2052_
timestamp 1698431365
transform -1 0 22512 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2053_
timestamp 1698431365
transform 1 0 21504 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _2054_
timestamp 1698431365
transform -1 0 23296 0 1 18816
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2055_
timestamp 1698431365
transform -1 0 21056 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2056_
timestamp 1698431365
transform -1 0 22624 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2057_
timestamp 1698431365
transform -1 0 20496 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2058_
timestamp 1698431365
transform 1 0 18144 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2059_
timestamp 1698431365
transform 1 0 17360 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2060_
timestamp 1698431365
transform 1 0 24304 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2061_
timestamp 1698431365
transform 1 0 33152 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2062_
timestamp 1698431365
transform 1 0 34160 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2063_
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2064_
timestamp 1698431365
transform 1 0 32928 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2065_
timestamp 1698431365
transform -1 0 35056 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2066_
timestamp 1698431365
transform -1 0 27216 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2067_
timestamp 1698431365
transform 1 0 25984 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2068_
timestamp 1698431365
transform 1 0 31584 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2069_
timestamp 1698431365
transform -1 0 35168 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2070_
timestamp 1698431365
transform -1 0 32704 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2071_
timestamp 1698431365
transform -1 0 26544 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2072_
timestamp 1698431365
transform -1 0 23072 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2073_
timestamp 1698431365
transform -1 0 3248 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2074_
timestamp 1698431365
transform -1 0 23856 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2075_
timestamp 1698431365
transform -1 0 35056 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2076_
timestamp 1698431365
transform 1 0 32592 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2077_
timestamp 1698431365
transform -1 0 23632 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2078_
timestamp 1698431365
transform 1 0 31024 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2079_
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2080_
timestamp 1698431365
transform 1 0 30128 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2081_
timestamp 1698431365
transform -1 0 24192 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2082_
timestamp 1698431365
transform 1 0 22624 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2083_
timestamp 1698431365
transform -1 0 22512 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2084_
timestamp 1698431365
transform 1 0 20384 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2085_
timestamp 1698431365
transform 1 0 20944 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2086_
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2087_
timestamp 1698431365
transform 1 0 21504 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2088_
timestamp 1698431365
transform -1 0 23520 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2089_
timestamp 1698431365
transform -1 0 26656 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2090_
timestamp 1698431365
transform 1 0 24080 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2091_
timestamp 1698431365
transform -1 0 24864 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2092_
timestamp 1698431365
transform -1 0 26992 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2093_
timestamp 1698431365
transform -1 0 26432 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2094_
timestamp 1698431365
transform -1 0 24864 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2095_
timestamp 1698431365
transform 1 0 22512 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2096_
timestamp 1698431365
transform -1 0 21168 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2097_
timestamp 1698431365
transform 1 0 20384 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2098_
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2099_
timestamp 1698431365
transform -1 0 26656 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2100_
timestamp 1698431365
transform 1 0 24640 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2101_
timestamp 1698431365
transform 1 0 21504 0 1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2102_
timestamp 1698431365
transform -1 0 24080 0 -1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2103_
timestamp 1698431365
transform 1 0 18592 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2104_
timestamp 1698431365
transform 1 0 18256 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2105_
timestamp 1698431365
transform -1 0 20384 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2106_
timestamp 1698431365
transform 1 0 19152 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2107_
timestamp 1698431365
transform -1 0 27888 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2108_
timestamp 1698431365
transform 1 0 25424 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2109_
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2110_
timestamp 1698431365
transform -1 0 21728 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2111_
timestamp 1698431365
transform 1 0 21056 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2112_
timestamp 1698431365
transform 1 0 31808 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2113_
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2114_
timestamp 1698431365
transform 1 0 23744 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2115_
timestamp 1698431365
transform -1 0 24752 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2116_
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2117_
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2118_
timestamp 1698431365
transform 1 0 21840 0 -1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2119_
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2120_
timestamp 1698431365
transform 1 0 21056 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2121_
timestamp 1698431365
transform -1 0 25424 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2122_
timestamp 1698431365
transform 1 0 23856 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2123_
timestamp 1698431365
transform 1 0 22288 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2124_
timestamp 1698431365
transform -1 0 7504 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2125_
timestamp 1698431365
transform -1 0 17024 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2126_
timestamp 1698431365
transform -1 0 16800 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2127_
timestamp 1698431365
transform 1 0 7840 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2128_
timestamp 1698431365
transform -1 0 8960 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2129_
timestamp 1698431365
transform -1 0 5152 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2130_
timestamp 1698431365
transform 1 0 3920 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2131_
timestamp 1698431365
transform -1 0 7616 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2132_
timestamp 1698431365
transform -1 0 5152 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2133_
timestamp 1698431365
transform -1 0 6160 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7952 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2135_
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2136_
timestamp 1698431365
transform 1 0 6160 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2137_
timestamp 1698431365
transform 1 0 8736 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2138_
timestamp 1698431365
transform 1 0 5936 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2139_
timestamp 1698431365
transform -1 0 8512 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2140_
timestamp 1698431365
transform 1 0 6832 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2141_
timestamp 1698431365
transform -1 0 8064 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2142_
timestamp 1698431365
transform -1 0 3024 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2143_
timestamp 1698431365
transform -1 0 4144 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2144_
timestamp 1698431365
transform -1 0 7056 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2145_
timestamp 1698431365
transform -1 0 7504 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2146_
timestamp 1698431365
transform 1 0 5264 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2147_
timestamp 1698431365
transform 1 0 2576 0 -1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2148_
timestamp 1698431365
transform 1 0 4480 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2149_
timestamp 1698431365
transform -1 0 9408 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2150_
timestamp 1698431365
transform -1 0 6496 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2151_
timestamp 1698431365
transform -1 0 5264 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2152_
timestamp 1698431365
transform 1 0 5600 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2153_
timestamp 1698431365
transform -1 0 8512 0 1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2154_
timestamp 1698431365
transform 1 0 7952 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2155_
timestamp 1698431365
transform -1 0 14000 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2156_
timestamp 1698431365
transform 1 0 9408 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2157_
timestamp 1698431365
transform 1 0 9744 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2158_
timestamp 1698431365
transform -1 0 10976 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2159_
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2160_
timestamp 1698431365
transform -1 0 31472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2161_
timestamp 1698431365
transform -1 0 11760 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2162_
timestamp 1698431365
transform 1 0 11760 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2163_
timestamp 1698431365
transform 1 0 13104 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2164_
timestamp 1698431365
transform -1 0 15904 0 1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2165_
timestamp 1698431365
transform 1 0 12432 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2166_
timestamp 1698431365
transform 1 0 12880 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2167_
timestamp 1698431365
transform 1 0 12656 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2168_
timestamp 1698431365
transform 1 0 12096 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2169_
timestamp 1698431365
transform -1 0 14224 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2170_
timestamp 1698431365
transform -1 0 14672 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2171_
timestamp 1698431365
transform -1 0 3696 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2172_
timestamp 1698431365
transform -1 0 13104 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2173_
timestamp 1698431365
transform -1 0 14560 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2174_
timestamp 1698431365
transform -1 0 15792 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2175_
timestamp 1698431365
transform 1 0 12544 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2176_
timestamp 1698431365
transform 1 0 13440 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2177_
timestamp 1698431365
transform 1 0 16352 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2178_
timestamp 1698431365
transform -1 0 9520 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2179_
timestamp 1698431365
transform -1 0 8176 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2180_
timestamp 1698431365
transform -1 0 2912 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2181_
timestamp 1698431365
transform -1 0 48160 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2182_
timestamp 1698431365
transform 1 0 46592 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2183_
timestamp 1698431365
transform 1 0 50176 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2184_
timestamp 1698431365
transform 1 0 47824 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2185_
timestamp 1698431365
transform 1 0 18816 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2186_
timestamp 1698431365
transform 1 0 47152 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2187_
timestamp 1698431365
transform 1 0 48720 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2188_
timestamp 1698431365
transform 1 0 48496 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2189_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 50176 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2190_
timestamp 1698431365
transform -1 0 46256 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2191_
timestamp 1698431365
transform -1 0 48048 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2192_
timestamp 1698431365
transform 1 0 49280 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2193_
timestamp 1698431365
transform 1 0 46032 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2194_
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2195_
timestamp 1698431365
transform 1 0 47488 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2196_
timestamp 1698431365
transform 1 0 50624 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2197_
timestamp 1698431365
transform 1 0 49952 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2198_
timestamp 1698431365
transform 1 0 50176 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2199_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40544 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2200_
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2201_
timestamp 1698431365
transform 1 0 50736 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2202_
timestamp 1698431365
transform -1 0 48384 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2203_
timestamp 1698431365
transform 1 0 50064 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2204_
timestamp 1698431365
transform -1 0 34944 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2205_
timestamp 1698431365
transform 1 0 47712 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2206_
timestamp 1698431365
transform 1 0 51296 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2207_
timestamp 1698431365
transform 1 0 51296 0 -1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2208_
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2209_
timestamp 1698431365
transform -1 0 53984 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2210_
timestamp 1698431365
transform -1 0 51408 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2211_
timestamp 1698431365
transform 1 0 49952 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2212_
timestamp 1698431365
transform -1 0 46480 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2213_
timestamp 1698431365
transform 1 0 47152 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2214_
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2215_
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2216_
timestamp 1698431365
transform 1 0 46256 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2217_
timestamp 1698431365
transform 1 0 45136 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2218_
timestamp 1698431365
transform 1 0 48384 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2219_
timestamp 1698431365
transform -1 0 52416 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2220_
timestamp 1698431365
transform 1 0 51408 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2221_
timestamp 1698431365
transform 1 0 53872 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2222_
timestamp 1698431365
transform -1 0 54992 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2223_
timestamp 1698431365
transform -1 0 54544 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2224_
timestamp 1698431365
transform 1 0 53872 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2225_
timestamp 1698431365
transform 1 0 53088 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2226_
timestamp 1698431365
transform -1 0 55328 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2227_
timestamp 1698431365
transform 1 0 36288 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2228_
timestamp 1698431365
transform 1 0 46256 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2229_
timestamp 1698431365
transform 1 0 45584 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2230_
timestamp 1698431365
transform 1 0 53424 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2231_
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2232_
timestamp 1698431365
transform 1 0 51408 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2233_
timestamp 1698431365
transform -1 0 53312 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2234_
timestamp 1698431365
transform 1 0 50176 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2235_
timestamp 1698431365
transform 1 0 34944 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2236_
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2237_
timestamp 1698431365
transform -1 0 49952 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2238_
timestamp 1698431365
transform 1 0 52752 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2239_
timestamp 1698431365
transform 1 0 53648 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2240_
timestamp 1698431365
transform -1 0 57792 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2241_
timestamp 1698431365
transform 1 0 56448 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2242_
timestamp 1698431365
transform 1 0 56448 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2243_
timestamp 1698431365
transform -1 0 57792 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2244_
timestamp 1698431365
transform -1 0 57680 0 1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2245_
timestamp 1698431365
transform -1 0 44240 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2246_
timestamp 1698431365
transform -1 0 56224 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2247_
timestamp 1698431365
transform -1 0 58352 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2248_
timestamp 1698431365
transform 1 0 55552 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2249_
timestamp 1698431365
transform -1 0 58352 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2250_
timestamp 1698431365
transform -1 0 58352 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2251_
timestamp 1698431365
transform 1 0 51856 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2252_
timestamp 1698431365
transform -1 0 56336 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2253_
timestamp 1698431365
transform -1 0 56224 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2254_
timestamp 1698431365
transform 1 0 55216 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2255_
timestamp 1698431365
transform 1 0 53760 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2256_
timestamp 1698431365
transform 1 0 54096 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2257_
timestamp 1698431365
transform 1 0 47264 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2258_
timestamp 1698431365
transform 1 0 50848 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2259_
timestamp 1698431365
transform 1 0 49728 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2260_
timestamp 1698431365
transform 1 0 51408 0 -1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2261_
timestamp 1698431365
transform 1 0 55440 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2262_
timestamp 1698431365
transform 1 0 43008 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2263_
timestamp 1698431365
transform 1 0 43680 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2264_
timestamp 1698431365
transform 1 0 46032 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2265_
timestamp 1698431365
transform -1 0 48832 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2266_
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2267_
timestamp 1698431365
transform 1 0 53872 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2268_
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2269_
timestamp 1698431365
transform 1 0 56336 0 1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2270_
timestamp 1698431365
transform -1 0 58352 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2271_
timestamp 1698431365
transform -1 0 58016 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2272_
timestamp 1698431365
transform 1 0 38528 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2273_
timestamp 1698431365
transform -1 0 40768 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2274_
timestamp 1698431365
transform -1 0 33712 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2275_
timestamp 1698431365
transform 1 0 39872 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2276_
timestamp 1698431365
transform -1 0 40544 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2277_
timestamp 1698431365
transform 1 0 53200 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2278_
timestamp 1698431365
transform 1 0 56896 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2279_
timestamp 1698431365
transform -1 0 58240 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2280_
timestamp 1698431365
transform -1 0 47376 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2281_
timestamp 1698431365
transform -1 0 48384 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2282_
timestamp 1698431365
transform 1 0 54208 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2283_
timestamp 1698431365
transform 1 0 46816 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2284_
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2285_
timestamp 1698431365
transform -1 0 56112 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2286_
timestamp 1698431365
transform 1 0 55552 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2287_
timestamp 1698431365
transform -1 0 55776 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2288_
timestamp 1698431365
transform 1 0 50288 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2289_
timestamp 1698431365
transform -1 0 52640 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2290_
timestamp 1698431365
transform 1 0 51184 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2291_
timestamp 1698431365
transform -1 0 36624 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2292_
timestamp 1698431365
transform 1 0 37520 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2293_
timestamp 1698431365
transform -1 0 41328 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2294_
timestamp 1698431365
transform -1 0 41104 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2295_
timestamp 1698431365
transform 1 0 40880 0 1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2296_
timestamp 1698431365
transform 1 0 50512 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2297_
timestamp 1698431365
transform -1 0 49616 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2298_
timestamp 1698431365
transform 1 0 47152 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2299_
timestamp 1698431365
transform -1 0 49056 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2300_
timestamp 1698431365
transform 1 0 48384 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2301_
timestamp 1698431365
transform 1 0 50960 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2302_
timestamp 1698431365
transform 1 0 52752 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2303_
timestamp 1698431365
transform -1 0 56224 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2304_
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2305_
timestamp 1698431365
transform -1 0 58352 0 1 28224
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2306_
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2307_
timestamp 1698431365
transform -1 0 56672 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2308_
timestamp 1698431365
transform -1 0 58352 0 1 9408
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2309_
timestamp 1698431365
transform -1 0 58352 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2310_
timestamp 1698431365
transform 1 0 27216 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2311_
timestamp 1698431365
transform -1 0 30352 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2312_
timestamp 1698431365
transform 1 0 29232 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2313_
timestamp 1698431365
transform -1 0 28224 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2314_
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2315_
timestamp 1698431365
transform -1 0 58240 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2316_
timestamp 1698431365
transform 1 0 53984 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2317_
timestamp 1698431365
transform 1 0 55664 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2318_
timestamp 1698431365
transform 1 0 57456 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2319_
timestamp 1698431365
transform -1 0 57904 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2320_
timestamp 1698431365
transform 1 0 50960 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2321_
timestamp 1698431365
transform 1 0 54656 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2322_
timestamp 1698431365
transform 1 0 53984 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2323_
timestamp 1698431365
transform -1 0 53088 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2324_
timestamp 1698431365
transform 1 0 50400 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2325_
timestamp 1698431365
transform 1 0 40320 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2326_
timestamp 1698431365
transform -1 0 41888 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2327_
timestamp 1698431365
transform 1 0 40992 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2328_
timestamp 1698431365
transform -1 0 39648 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2329_
timestamp 1698431365
transform -1 0 45584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2330_
timestamp 1698431365
transform -1 0 39648 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2331_
timestamp 1698431365
transform 1 0 38528 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2332_
timestamp 1698431365
transform 1 0 41328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2333_
timestamp 1698431365
transform 1 0 40768 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2334_
timestamp 1698431365
transform -1 0 43120 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2335_
timestamp 1698431365
transform -1 0 38528 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2336_
timestamp 1698431365
transform 1 0 36624 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2337_
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2338_
timestamp 1698431365
transform 1 0 41888 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2339_
timestamp 1698431365
transform 1 0 50736 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2340_
timestamp 1698431365
transform -1 0 50736 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2341_
timestamp 1698431365
transform 1 0 49392 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2342_
timestamp 1698431365
transform 1 0 49056 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2343_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2344_
timestamp 1698431365
transform 1 0 47488 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2345_
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2346_
timestamp 1698431365
transform 1 0 48048 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2347_
timestamp 1698431365
transform -1 0 48048 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2348_
timestamp 1698431365
transform 1 0 46144 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2349_
timestamp 1698431365
transform 1 0 46144 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2350_
timestamp 1698431365
transform 1 0 48720 0 1 29792
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2351_
timestamp 1698431365
transform 1 0 50960 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2352_
timestamp 1698431365
transform -1 0 57456 0 1 29792
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2353_
timestamp 1698431365
transform -1 0 57904 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2354_
timestamp 1698431365
transform 1 0 26768 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2355_
timestamp 1698431365
transform 1 0 27104 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2356_
timestamp 1698431365
transform 1 0 27888 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2357_
timestamp 1698431365
transform 1 0 27888 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2358_
timestamp 1698431365
transform 1 0 28112 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2359_
timestamp 1698431365
transform -1 0 57792 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2360_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 55328 0 1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2361_
timestamp 1698431365
transform -1 0 55664 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2362_
timestamp 1698431365
transform -1 0 55104 0 -1 31360
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2363_
timestamp 1698431365
transform -1 0 48384 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2364_
timestamp 1698431365
transform -1 0 49392 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2365_
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2366_
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2367_
timestamp 1698431365
transform -1 0 42560 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2368_
timestamp 1698431365
transform 1 0 33264 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2369_
timestamp 1698431365
transform 1 0 31696 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2370_
timestamp 1698431365
transform 1 0 32368 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2371_
timestamp 1698431365
transform -1 0 32704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2372_
timestamp 1698431365
transform -1 0 34496 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2373_
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2374_
timestamp 1698431365
transform -1 0 34048 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2375_
timestamp 1698431365
transform -1 0 32704 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2376_
timestamp 1698431365
transform -1 0 30688 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2377_
timestamp 1698431365
transform -1 0 32368 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2378_
timestamp 1698431365
transform -1 0 36400 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2379_
timestamp 1698431365
transform 1 0 35056 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2380_
timestamp 1698431365
transform -1 0 36400 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2381_
timestamp 1698431365
transform 1 0 31360 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2382_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2383_
timestamp 1698431365
transform 1 0 41776 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2384_
timestamp 1698431365
transform 1 0 44800 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2385_
timestamp 1698431365
transform 1 0 46816 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2386_
timestamp 1698431365
transform -1 0 48384 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2387_
timestamp 1698431365
transform 1 0 37856 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2388_
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2389_
timestamp 1698431365
transform 1 0 38304 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2390_
timestamp 1698431365
transform -1 0 40432 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2391_
timestamp 1698431365
transform 1 0 15232 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2392_
timestamp 1698431365
transform -1 0 35168 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2393_
timestamp 1698431365
transform 1 0 16240 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2394_
timestamp 1698431365
transform 1 0 22064 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2395_
timestamp 1698431365
transform 1 0 33488 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2396_
timestamp 1698431365
transform 1 0 36512 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2397_
timestamp 1698431365
transform 1 0 39872 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2398_
timestamp 1698431365
transform 1 0 42224 0 -1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2399_
timestamp 1698431365
transform 1 0 47376 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2400_
timestamp 1698431365
transform -1 0 51184 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2401_
timestamp 1698431365
transform -1 0 30688 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2402_
timestamp 1698431365
transform 1 0 28784 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2403_
timestamp 1698431365
transform -1 0 30128 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2404_
timestamp 1698431365
transform -1 0 27776 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2405_
timestamp 1698431365
transform -1 0 20608 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  _2406_
timestamp 1698431365
transform -1 0 50512 0 -1 29792
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2407_
timestamp 1698431365
transform 1 0 49056 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2408_
timestamp 1698431365
transform 1 0 45248 0 1 31360
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2409_
timestamp 1698431365
transform 1 0 45584 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2410_
timestamp 1698431365
transform -1 0 48384 0 -1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2411_
timestamp 1698431365
transform 1 0 41664 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2412_
timestamp 1698431365
transform -1 0 45696 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2413_
timestamp 1698431365
transform -1 0 44352 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2414_
timestamp 1698431365
transform -1 0 40208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2415_
timestamp 1698431365
transform 1 0 39200 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2416_
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2417_
timestamp 1698431365
transform 1 0 38416 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2418_
timestamp 1698431365
transform 1 0 43120 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2419_
timestamp 1698431365
transform -1 0 43568 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2420_
timestamp 1698431365
transform -1 0 32592 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2421_
timestamp 1698431365
transform -1 0 31696 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2422_
timestamp 1698431365
transform -1 0 29680 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2423_
timestamp 1698431365
transform -1 0 26432 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2424_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _2425_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26432 0 -1 21952
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2426_
timestamp 1698431365
transform 1 0 26208 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2427_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2428_
timestamp 1698431365
transform 1 0 30464 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2429_
timestamp 1698431365
transform 1 0 31808 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2430_
timestamp 1698431365
transform 1 0 33936 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2431_
timestamp 1698431365
transform -1 0 35728 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2432_
timestamp 1698431365
transform 1 0 35616 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2433_
timestamp 1698431365
transform -1 0 34272 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2434_
timestamp 1698431365
transform -1 0 23184 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2435_
timestamp 1698431365
transform -1 0 24864 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2436_
timestamp 1698431365
transform 1 0 23184 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2437_
timestamp 1698431365
transform -1 0 28448 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2438_
timestamp 1698431365
transform 1 0 27664 0 -1 26656
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2439_
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2440_
timestamp 1698431365
transform -1 0 31136 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2441_
timestamp 1698431365
transform -1 0 32256 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2442_
timestamp 1698431365
transform -1 0 19824 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2443_
timestamp 1698431365
transform 1 0 18592 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2444_
timestamp 1698431365
transform -1 0 16128 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2445_
timestamp 1698431365
transform -1 0 17584 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2446_
timestamp 1698431365
transform -1 0 20720 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2447_
timestamp 1698431365
transform -1 0 19600 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2448_
timestamp 1698431365
transform -1 0 28672 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2449_
timestamp 1698431365
transform -1 0 29680 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2450_
timestamp 1698431365
transform 1 0 28672 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2451_
timestamp 1698431365
transform 1 0 30576 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2452_
timestamp 1698431365
transform -1 0 31696 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2453_
timestamp 1698431365
transform 1 0 31136 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2454_
timestamp 1698431365
transform -1 0 31024 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2455_
timestamp 1698431365
transform 1 0 23520 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2456_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2457_
timestamp 1698431365
transform 1 0 26992 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2458_
timestamp 1698431365
transform 1 0 28336 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2459_
timestamp 1698431365
transform -1 0 26432 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2460_
timestamp 1698431365
transform 1 0 31920 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2461_
timestamp 1698431365
transform -1 0 32480 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2462_
timestamp 1698431365
transform 1 0 22512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2463_
timestamp 1698431365
transform 1 0 23408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2464_
timestamp 1698431365
transform 1 0 23520 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2465_
timestamp 1698431365
transform -1 0 31136 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2466_
timestamp 1698431365
transform 1 0 24752 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2467_
timestamp 1698431365
transform 1 0 17920 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2468_
timestamp 1698431365
transform -1 0 20832 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2469_
timestamp 1698431365
transform -1 0 19936 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2470_
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2471_
timestamp 1698431365
transform -1 0 20048 0 -1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2472_
timestamp 1698431365
transform -1 0 28784 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2473_
timestamp 1698431365
transform 1 0 27552 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2474_
timestamp 1698431365
transform -1 0 26208 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2475_
timestamp 1698431365
transform 1 0 25648 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2476_
timestamp 1698431365
transform 1 0 26208 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2477_
timestamp 1698431365
transform -1 0 27440 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2478_
timestamp 1698431365
transform -1 0 26432 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2479_
timestamp 1698431365
transform -1 0 16800 0 -1 26656
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2480_
timestamp 1698431365
transform -1 0 16128 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2481_
timestamp 1698431365
transform 1 0 14224 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2482_
timestamp 1698431365
transform -1 0 15456 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2483_
timestamp 1698431365
transform -1 0 15008 0 -1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2484_
timestamp 1698431365
transform -1 0 14112 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2485_
timestamp 1698431365
transform -1 0 16576 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2486_
timestamp 1698431365
transform -1 0 16688 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2487_
timestamp 1698431365
transform 1 0 15008 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2488_
timestamp 1698431365
transform 1 0 15568 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2489_
timestamp 1698431365
transform 1 0 14672 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2490_
timestamp 1698431365
transform 1 0 14896 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2491_
timestamp 1698431365
transform 1 0 16240 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2492_
timestamp 1698431365
transform 1 0 15344 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2493_
timestamp 1698431365
transform -1 0 18816 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2494_
timestamp 1698431365
transform 1 0 18480 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2495_
timestamp 1698431365
transform 1 0 19376 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2496_
timestamp 1698431365
transform 1 0 20160 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2497_
timestamp 1698431365
transform -1 0 20160 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2498_
timestamp 1698431365
transform -1 0 21952 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2499_
timestamp 1698431365
transform -1 0 25536 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2500_
timestamp 1698431365
transform -1 0 24864 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2501_
timestamp 1698431365
transform 1 0 21168 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2502_
timestamp 1698431365
transform -1 0 18144 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2503_
timestamp 1698431365
transform 1 0 18144 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2504_
timestamp 1698431365
transform -1 0 19936 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2505_
timestamp 1698431365
transform 1 0 23856 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2506_
timestamp 1698431365
transform -1 0 31920 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2507_
timestamp 1698431365
transform 1 0 27440 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2508_
timestamp 1698431365
transform -1 0 24864 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2509_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2510_
timestamp 1698431365
transform 1 0 20832 0 -1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2511_
timestamp 1698431365
transform 1 0 14448 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2512_
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2513_
timestamp 1698431365
transform 1 0 14560 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2514_
timestamp 1698431365
transform 1 0 16128 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2515_
timestamp 1698431365
transform 1 0 43568 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2516_
timestamp 1698431365
transform -1 0 49728 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2517_
timestamp 1698431365
transform 1 0 12096 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2518_
timestamp 1698431365
transform 1 0 11200 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _2519_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2520_
timestamp 1698431365
transform -1 0 14448 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2521_
timestamp 1698431365
transform -1 0 8848 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2522_
timestamp 1698431365
transform -1 0 6384 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2523_
timestamp 1698431365
transform -1 0 5040 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2524_
timestamp 1698431365
transform -1 0 11648 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2525_
timestamp 1698431365
transform -1 0 10080 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2526_
timestamp 1698431365
transform -1 0 10864 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2527_
timestamp 1698431365
transform -1 0 13664 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2528_
timestamp 1698431365
transform -1 0 11536 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2529_
timestamp 1698431365
transform -1 0 11088 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2530_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2531_
timestamp 1698431365
transform -1 0 10416 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2532_
timestamp 1698431365
transform 1 0 11088 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2533_
timestamp 1698431365
transform 1 0 10528 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2534_
timestamp 1698431365
transform 1 0 11312 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2535_
timestamp 1698431365
transform -1 0 11312 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2536_
timestamp 1698431365
transform 1 0 11200 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2537_
timestamp 1698431365
transform -1 0 5712 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2538_
timestamp 1698431365
transform 1 0 12544 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2539_
timestamp 1698431365
transform 1 0 12096 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2540_
timestamp 1698431365
transform -1 0 10976 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2541_
timestamp 1698431365
transform -1 0 11088 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2542_
timestamp 1698431365
transform -1 0 4704 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2543_
timestamp 1698431365
transform 1 0 2912 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2544_
timestamp 1698431365
transform -1 0 3920 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2545_
timestamp 1698431365
transform 1 0 7280 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2546_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2547_
timestamp 1698431365
transform -1 0 3808 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2548_
timestamp 1698431365
transform 1 0 2576 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2549_
timestamp 1698431365
transform -1 0 4928 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2550_
timestamp 1698431365
transform -1 0 2576 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2551_
timestamp 1698431365
transform -1 0 2688 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2552_
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2553_
timestamp 1698431365
transform -1 0 9968 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2554_
timestamp 1698431365
transform 1 0 13216 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2555_
timestamp 1698431365
transform 1 0 12432 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2556_
timestamp 1698431365
transform 1 0 12320 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2557_
timestamp 1698431365
transform -1 0 11088 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2558_
timestamp 1698431365
transform 1 0 6384 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2559_
timestamp 1698431365
transform 1 0 10080 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2560_
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2561_
timestamp 1698431365
transform -1 0 29680 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2562_
timestamp 1698431365
transform 1 0 7840 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2563_
timestamp 1698431365
transform 1 0 8400 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2564_
timestamp 1698431365
transform -1 0 7728 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2565_
timestamp 1698431365
transform 1 0 5936 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2566_
timestamp 1698431365
transform -1 0 9968 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2567_
timestamp 1698431365
transform 1 0 9968 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2568_
timestamp 1698431365
transform 1 0 13888 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2569_
timestamp 1698431365
transform 1 0 15456 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2570_
timestamp 1698431365
transform -1 0 15232 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2571_
timestamp 1698431365
transform -1 0 16016 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2572_
timestamp 1698431365
transform 1 0 15232 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2573_
timestamp 1698431365
transform -1 0 18368 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2574_
timestamp 1698431365
transform 1 0 13888 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2575_
timestamp 1698431365
transform 1 0 16352 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2576_
timestamp 1698431365
transform -1 0 12656 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2577_
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2578_
timestamp 1698431365
transform -1 0 15456 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2579_
timestamp 1698431365
transform 1 0 16128 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2580_
timestamp 1698431365
transform -1 0 6160 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2581_
timestamp 1698431365
transform -1 0 18368 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2582_
timestamp 1698431365
transform -1 0 15456 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2583_
timestamp 1698431365
transform -1 0 17024 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2584_
timestamp 1698431365
transform 1 0 15680 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2585_
timestamp 1698431365
transform -1 0 17024 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2586_
timestamp 1698431365
transform -1 0 15456 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2587_
timestamp 1698431365
transform 1 0 12544 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2588_
timestamp 1698431365
transform 1 0 14000 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2589_
timestamp 1698431365
transform -1 0 14896 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2590_
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2591_
timestamp 1698431365
transform 1 0 7504 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2592_
timestamp 1698431365
transform 1 0 8176 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2593_
timestamp 1698431365
transform -1 0 14224 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2594_
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2595_
timestamp 1698431365
transform 1 0 2576 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2596_
timestamp 1698431365
transform 1 0 3808 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2597_
timestamp 1698431365
transform 1 0 3248 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2598_
timestamp 1698431365
transform -1 0 9632 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2599_
timestamp 1698431365
transform 1 0 6944 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2600_
timestamp 1698431365
transform -1 0 8400 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2601_
timestamp 1698431365
transform 1 0 3808 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2602_
timestamp 1698431365
transform 1 0 6384 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2603_
timestamp 1698431365
transform -1 0 9184 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2604_
timestamp 1698431365
transform 1 0 4368 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2605_
timestamp 1698431365
transform 1 0 6048 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2606_
timestamp 1698431365
transform -1 0 7840 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2607_
timestamp 1698431365
transform 1 0 4256 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2608_
timestamp 1698431365
transform 1 0 5824 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2609_
timestamp 1698431365
transform -1 0 7280 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2610_
timestamp 1698431365
transform -1 0 3584 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2611_
timestamp 1698431365
transform 1 0 4256 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2612_
timestamp 1698431365
transform -1 0 10080 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2613_
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2614_
timestamp 1698431365
transform -1 0 8624 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2615_
timestamp 1698431365
transform 1 0 3248 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2616_
timestamp 1698431365
transform 1 0 7392 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2617_
timestamp 1698431365
transform -1 0 6944 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2618_
timestamp 1698431365
transform 1 0 1680 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2619_
timestamp 1698431365
transform 1 0 4256 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2620_
timestamp 1698431365
transform 1 0 10528 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2621_
timestamp 1698431365
transform 1 0 3472 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2622_
timestamp 1698431365
transform -1 0 10976 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2623_
timestamp 1698431365
transform 1 0 9744 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2624_
timestamp 1698431365
transform 1 0 10192 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2625_
timestamp 1698431365
transform 1 0 10416 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2626_
timestamp 1698431365
transform 1 0 12208 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2627_
timestamp 1698431365
transform 1 0 35728 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2628_
timestamp 1698431365
transform 1 0 11312 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2629_
timestamp 1698431365
transform 1 0 12320 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2630_
timestamp 1698431365
transform 1 0 18144 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2631_
timestamp 1698431365
transform 1 0 35056 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2632_
timestamp 1698431365
transform -1 0 37184 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2633_
timestamp 1698431365
transform 1 0 36064 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2634_
timestamp 1698431365
transform 1 0 17584 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2635_
timestamp 1698431365
transform -1 0 37744 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2636_
timestamp 1698431365
transform -1 0 38080 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2637_
timestamp 1698431365
transform 1 0 15680 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2638_
timestamp 1698431365
transform -1 0 37520 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2639_
timestamp 1698431365
transform -1 0 38976 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2640_
timestamp 1698431365
transform 1 0 17472 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2641_
timestamp 1698431365
transform 1 0 35728 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2642_
timestamp 1698431365
transform 1 0 11760 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2643_
timestamp 1698431365
transform -1 0 12208 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2644_
timestamp 1698431365
transform -1 0 11088 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2645_
timestamp 1698431365
transform 1 0 10192 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2646_
timestamp 1698431365
transform 1 0 10192 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2647_
timestamp 1698431365
transform 1 0 10752 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2648_
timestamp 1698431365
transform -1 0 12320 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2649_
timestamp 1698431365
transform 1 0 9968 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2650_
timestamp 1698431365
transform 1 0 10864 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2651_
timestamp 1698431365
transform -1 0 12544 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2652_
timestamp 1698431365
transform 1 0 10528 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2653_
timestamp 1698431365
transform 1 0 11088 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2654_
timestamp 1698431365
transform 1 0 12544 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2655_
timestamp 1698431365
transform -1 0 10192 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2656_
timestamp 1698431365
transform 1 0 10192 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2657_
timestamp 1698431365
transform -1 0 9072 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2658_
timestamp 1698431365
transform -1 0 3360 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2659_
timestamp 1698431365
transform 1 0 3696 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2660_
timestamp 1698431365
transform 1 0 3024 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2661_
timestamp 1698431365
transform 1 0 8736 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2662_
timestamp 1698431365
transform 1 0 3808 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2663_
timestamp 1698431365
transform -1 0 4368 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2664_
timestamp 1698431365
transform -1 0 3584 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2665_
timestamp 1698431365
transform -1 0 4704 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2666_
timestamp 1698431365
transform 1 0 2912 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2667_
timestamp 1698431365
transform 1 0 4368 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2668_
timestamp 1698431365
transform 1 0 1904 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2669_
timestamp 1698431365
transform 1 0 2800 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2670_
timestamp 1698431365
transform -1 0 4256 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2671_
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2672_
timestamp 1698431365
transform 1 0 2800 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2673_
timestamp 1698431365
transform -1 0 4256 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2674_
timestamp 1698431365
transform 1 0 2240 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2675_
timestamp 1698431365
transform -1 0 3472 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2676_
timestamp 1698431365
transform 1 0 2800 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2677_
timestamp 1698431365
transform -1 0 4368 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2678_
timestamp 1698431365
transform -1 0 4928 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2679_
timestamp 1698431365
transform -1 0 8960 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2680_
timestamp 1698431365
transform 1 0 2240 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2681_
timestamp 1698431365
transform -1 0 6944 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2682_
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2683_
timestamp 1698431365
transform -1 0 4480 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2684_
timestamp 1698431365
transform 1 0 9072 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2685_
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2686_
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2687_
timestamp 1698431365
transform 1 0 11088 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2688_
timestamp 1698431365
transform 1 0 18032 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2689_
timestamp 1698431365
transform 1 0 17360 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2690_
timestamp 1698431365
transform -1 0 19936 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2691_
timestamp 1698431365
transform -1 0 19264 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2692_
timestamp 1698431365
transform 1 0 10752 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2693_
timestamp 1698431365
transform -1 0 11984 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2694_
timestamp 1698431365
transform -1 0 10304 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2695_
timestamp 1698431365
transform 1 0 10864 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2696_
timestamp 1698431365
transform -1 0 18704 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2697_
timestamp 1698431365
transform 1 0 15792 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2698_
timestamp 1698431365
transform 1 0 8848 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2699_
timestamp 1698431365
transform -1 0 15456 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2700_
timestamp 1698431365
transform -1 0 15232 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2701_
timestamp 1698431365
transform 1 0 14112 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2702_
timestamp 1698431365
transform 1 0 12544 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2703_
timestamp 1698431365
transform -1 0 16464 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2704_
timestamp 1698431365
transform -1 0 15792 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2705_
timestamp 1698431365
transform 1 0 13552 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2706_
timestamp 1698431365
transform 1 0 14672 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2707_
timestamp 1698431365
transform 1 0 15792 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2708_
timestamp 1698431365
transform 1 0 19712 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2709_
timestamp 1698431365
transform 1 0 15456 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2710_
timestamp 1698431365
transform 1 0 11760 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2711_
timestamp 1698431365
transform 1 0 13664 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2712_
timestamp 1698431365
transform -1 0 15456 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2713_
timestamp 1698431365
transform -1 0 11648 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2714_
timestamp 1698431365
transform -1 0 11312 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2715_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8848 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2716_
timestamp 1698431365
transform 1 0 10080 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2717_
timestamp 1698431365
transform -1 0 47040 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2718_
timestamp 1698431365
transform 1 0 32368 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2719_
timestamp 1698431365
transform 1 0 29456 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2720_
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2721_
timestamp 1698431365
transform 1 0 25872 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2722_
timestamp 1698431365
transform 1 0 18032 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2723_
timestamp 1698431365
transform 1 0 12544 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2724_
timestamp 1698431365
transform 1 0 15904 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2725_
timestamp 1698431365
transform 1 0 15120 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2726_
timestamp 1698431365
transform 1 0 12880 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2727_
timestamp 1698431365
transform 1 0 9520 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2728_
timestamp 1698431365
transform 1 0 8736 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2729_
timestamp 1698431365
transform 1 0 5712 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2730_
timestamp 1698431365
transform 1 0 4032 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2731_
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2732_
timestamp 1698431365
transform -1 0 8736 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2733_
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2734_
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2735_
timestamp 1698431365
transform -1 0 12656 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2736_
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2737_
timestamp 1698431365
transform 1 0 4144 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2738_
timestamp 1698431365
transform -1 0 12432 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2739_
timestamp 1698431365
transform 1 0 24752 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2740_
timestamp 1698431365
transform -1 0 20048 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2741_
timestamp 1698431365
transform 1 0 1680 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2742_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2743_
timestamp 1698431365
transform -1 0 14784 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2744_
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2745_
timestamp 1698431365
transform 1 0 1792 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2746_
timestamp 1698431365
transform 1 0 2352 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2747_
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2748_
timestamp 1698431365
transform 1 0 7616 0 1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2749_
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2750_
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2751_
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2752_
timestamp 1698431365
transform 1 0 14112 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2753_
timestamp 1698431365
transform 1 0 16576 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2754_
timestamp 1698431365
transform 1 0 14672 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2755_
timestamp 1698431365
transform 1 0 18928 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2756_
timestamp 1698431365
transform 1 0 16240 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2757_
timestamp 1698431365
transform 1 0 17472 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2758_
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2759_
timestamp 1698431365
transform 1 0 13776 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2760_
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2761_
timestamp 1698431365
transform 1 0 5600 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2762_
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2763_
timestamp 1698431365
transform 1 0 5040 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2764_
timestamp 1698431365
transform 1 0 5152 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2765_
timestamp 1698431365
transform 1 0 5936 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2766_
timestamp 1698431365
transform 1 0 2688 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2767_
timestamp 1698431365
transform 1 0 9856 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2768_
timestamp 1698431365
transform 1 0 37184 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2769_
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2770_
timestamp 1698431365
transform 1 0 37296 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2771_
timestamp 1698431365
transform 1 0 37072 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2772_
timestamp 1698431365
transform 1 0 10192 0 -1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2773_
timestamp 1698431365
transform 1 0 10528 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2774_
timestamp 1698431365
transform 1 0 11200 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2775_
timestamp 1698431365
transform 1 0 9968 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2776_
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2777_
timestamp 1698431365
transform 1 0 1792 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2778_
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2779_
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2780_
timestamp 1698431365
transform 1 0 1680 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2781_
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2782_
timestamp 1698431365
transform 1 0 3136 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2783_
timestamp 1698431365
transform -1 0 11312 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2784_
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2785_
timestamp 1698431365
transform 1 0 10304 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2786_
timestamp 1698431365
transform 1 0 13776 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2787_
timestamp 1698431365
transform 1 0 16464 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2788_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2789_
timestamp 1698431365
transform 1 0 19376 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2790_
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2791_
timestamp 1698431365
transform 1 0 9632 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1361__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__A2
timestamp 1698431365
transform 1 0 48160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__A2
timestamp 1698431365
transform 1 0 46144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1371__A1
timestamp 1698431365
transform -1 0 42336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1373__A2
timestamp 1698431365
transform 1 0 51744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__I
timestamp 1698431365
transform 1 0 17808 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1377__A2
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1379__A2
timestamp 1698431365
transform -1 0 35616 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1382__A1
timestamp 1698431365
transform 1 0 41888 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1384__A1
timestamp 1698431365
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__I
timestamp 1698431365
transform -1 0 12544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1391__A1
timestamp 1698431365
transform -1 0 16352 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1391__A2
timestamp 1698431365
transform 1 0 16352 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1395__I
timestamp 1698431365
transform 1 0 17472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__A1
timestamp 1698431365
transform 1 0 7616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__A2
timestamp 1698431365
transform 1 0 7280 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__A1
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__A2
timestamp 1698431365
transform 1 0 6832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__A1
timestamp 1698431365
transform -1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__A2
timestamp 1698431365
transform 1 0 7056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__A3
timestamp 1698431365
transform 1 0 44464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1425__I
timestamp 1698431365
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__A2
timestamp 1698431365
transform 1 0 43008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1442__A2
timestamp 1698431365
transform 1 0 43456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1449__I
timestamp 1698431365
transform 1 0 47376 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1453__I
timestamp 1698431365
transform 1 0 34384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1460__I
timestamp 1698431365
transform 1 0 53200 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__I
timestamp 1698431365
transform 1 0 43568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1481__A1
timestamp 1698431365
transform 1 0 38864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1504__A1
timestamp 1698431365
transform 1 0 50848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1504__A2
timestamp 1698431365
transform 1 0 51744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A2
timestamp 1698431365
transform 1 0 46032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__B2
timestamp 1698431365
transform 1 0 42560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1534__I
timestamp 1698431365
transform 1 0 31696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1543__A1
timestamp 1698431365
transform -1 0 27328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__A1
timestamp 1698431365
transform 1 0 34608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__A2
timestamp 1698431365
transform -1 0 33488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A1
timestamp 1698431365
transform 1 0 12432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__A2
timestamp 1698431365
transform 1 0 49952 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A1
timestamp 1698431365
transform 1 0 51296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A2
timestamp 1698431365
transform 1 0 51744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1583__I
timestamp 1698431365
transform 1 0 34384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__I
timestamp 1698431365
transform -1 0 40544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A1
timestamp 1698431365
transform -1 0 19824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A2
timestamp 1698431365
transform -1 0 20272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__I
timestamp 1698431365
transform -1 0 36512 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__A1
timestamp 1698431365
transform 1 0 49840 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A2
timestamp 1698431365
transform 1 0 37744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__A2
timestamp 1698431365
transform 1 0 35056 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1614__I
timestamp 1698431365
transform -1 0 28112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A1
timestamp 1698431365
transform -1 0 28112 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__A2
timestamp 1698431365
transform 1 0 37296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__A2
timestamp 1698431365
transform 1 0 15904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__I
timestamp 1698431365
transform 1 0 47376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A2
timestamp 1698431365
transform -1 0 45360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A2
timestamp 1698431365
transform 1 0 16352 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__A2
timestamp 1698431365
transform 1 0 45696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A1
timestamp 1698431365
transform 1 0 51072 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A2
timestamp 1698431365
transform 1 0 51744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__A1
timestamp 1698431365
transform 1 0 50400 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1698431365
transform -1 0 18928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A2
timestamp 1698431365
transform -1 0 20720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__I
timestamp 1698431365
transform -1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A1
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A2
timestamp 1698431365
transform 1 0 22176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A1
timestamp 1698431365
transform 1 0 50624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__A1
timestamp 1698431365
transform -1 0 45472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__A1
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__A1
timestamp 1698431365
transform 1 0 32144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__A1
timestamp 1698431365
transform 1 0 28896 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__A2
timestamp 1698431365
transform -1 0 34048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__A2
timestamp 1698431365
transform -1 0 53984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__A3
timestamp 1698431365
transform -1 0 54208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__I
timestamp 1698431365
transform -1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__A1
timestamp 1698431365
transform -1 0 49952 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__A1
timestamp 1698431365
transform 1 0 46480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__A2
timestamp 1698431365
transform 1 0 53312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A1
timestamp 1698431365
transform -1 0 47488 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A2
timestamp 1698431365
transform 1 0 50624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__A1
timestamp 1698431365
transform 1 0 19600 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__A2
timestamp 1698431365
transform 1 0 20048 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__I
timestamp 1698431365
transform 1 0 12320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A1
timestamp 1698431365
transform 1 0 20160 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A2
timestamp 1698431365
transform -1 0 21056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__A1
timestamp 1698431365
transform 1 0 52080 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__A2
timestamp 1698431365
transform 1 0 52080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__I
timestamp 1698431365
transform 1 0 39200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A1
timestamp 1698431365
transform -1 0 38976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__A2
timestamp 1698431365
transform -1 0 38080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__I
timestamp 1698431365
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__B2
timestamp 1698431365
transform -1 0 45808 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__A1
timestamp 1698431365
transform -1 0 35168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__I
timestamp 1698431365
transform 1 0 20944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__A2
timestamp 1698431365
transform 1 0 32480 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__A2
timestamp 1698431365
transform 1 0 34832 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__A1
timestamp 1698431365
transform -1 0 45248 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__A1
timestamp 1698431365
transform 1 0 43344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__A2
timestamp 1698431365
transform 1 0 58016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__A1
timestamp 1698431365
transform -1 0 58240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__A1
timestamp 1698431365
transform -1 0 18368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__A2
timestamp 1698431365
transform -1 0 18816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A1
timestamp 1698431365
transform -1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A2
timestamp 1698431365
transform 1 0 21952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A1
timestamp 1698431365
transform 1 0 58128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A1
timestamp 1698431365
transform 1 0 58128 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__I
timestamp 1698431365
transform 1 0 13664 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__I
timestamp 1698431365
transform 1 0 31472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__A1
timestamp 1698431365
transform 1 0 35280 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__A1
timestamp 1698431365
transform 1 0 38752 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__A2
timestamp 1698431365
transform -1 0 35056 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__I
timestamp 1698431365
transform 1 0 35280 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__A2
timestamp 1698431365
transform -1 0 38192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__I
timestamp 1698431365
transform -1 0 19152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1893__A1
timestamp 1698431365
transform -1 0 35616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__A2
timestamp 1698431365
transform 1 0 34384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__A2
timestamp 1698431365
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A1
timestamp 1698431365
transform 1 0 37632 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A2
timestamp 1698431365
transform -1 0 38304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__A1
timestamp 1698431365
transform 1 0 35728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__A1
timestamp 1698431365
transform -1 0 54544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__A2
timestamp 1698431365
transform -1 0 17920 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__A1
timestamp 1698431365
transform 1 0 55104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__A2
timestamp 1698431365
transform 1 0 17808 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__A1
timestamp 1698431365
transform -1 0 33936 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__A1
timestamp 1698431365
transform 1 0 34832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__A2
timestamp 1698431365
transform -1 0 33376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1967__A2
timestamp 1698431365
transform -1 0 34048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__B
timestamp 1698431365
transform 1 0 21728 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1977__A2
timestamp 1698431365
transform -1 0 27104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A1
timestamp 1698431365
transform 1 0 31696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__I
timestamp 1698431365
transform -1 0 13776 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__I
timestamp 1698431365
transform -1 0 14000 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__A2
timestamp 1698431365
transform 1 0 22848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__A1
timestamp 1698431365
transform -1 0 30128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__A1
timestamp 1698431365
transform -1 0 22624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__A2
timestamp 1698431365
transform 1 0 25648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__A1
timestamp 1698431365
transform -1 0 24528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__A1
timestamp 1698431365
transform -1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2007__A1
timestamp 1698431365
transform -1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__A1
timestamp 1698431365
transform 1 0 26096 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A1
timestamp 1698431365
transform 1 0 34496 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__A1
timestamp 1698431365
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__A1
timestamp 1698431365
transform -1 0 35056 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__A2
timestamp 1698431365
transform -1 0 31472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A1
timestamp 1698431365
transform -1 0 22848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A1
timestamp 1698431365
transform 1 0 29344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A2
timestamp 1698431365
transform 1 0 30688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A3
timestamp 1698431365
transform 1 0 27888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A2
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A1
timestamp 1698431365
transform -1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A2
timestamp 1698431365
transform -1 0 27440 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__A2
timestamp 1698431365
transform 1 0 21840 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__A1
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__A1
timestamp 1698431365
transform -1 0 32928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A1
timestamp 1698431365
transform -1 0 26992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__I
timestamp 1698431365
transform -1 0 12656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__A1
timestamp 1698431365
transform 1 0 23856 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2082__A1
timestamp 1698431365
transform 1 0 23744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2086__A1
timestamp 1698431365
transform 1 0 21952 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2089__A1
timestamp 1698431365
transform 1 0 26880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__A2
timestamp 1698431365
transform 1 0 24416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__A2
timestamp 1698431365
transform 1 0 24864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2099__A2
timestamp 1698431365
transform 1 0 27328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2103__A1
timestamp 1698431365
transform 1 0 20160 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A2
timestamp 1698431365
transform 1 0 21728 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2121__A1
timestamp 1698431365
transform 1 0 25648 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__I
timestamp 1698431365
transform 1 0 7504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__A1
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__A2
timestamp 1698431365
transform -1 0 14896 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__I
timestamp 1698431365
transform -1 0 15904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__I
timestamp 1698431365
transform -1 0 6160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2134__A3
timestamp 1698431365
transform -1 0 6160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2164__A1
timestamp 1698431365
transform 1 0 11872 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__I
timestamp 1698431365
transform 1 0 51520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__I
timestamp 1698431365
transform 1 0 50848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2185__I
timestamp 1698431365
transform 1 0 17584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2186__A1
timestamp 1698431365
transform 1 0 45136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__A1
timestamp 1698431365
transform 1 0 50848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A1
timestamp 1698431365
transform 1 0 49392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A2
timestamp 1698431365
transform 1 0 50288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A3
timestamp 1698431365
transform 1 0 48832 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2197__A1
timestamp 1698431365
transform 1 0 51296 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2199__I
timestamp 1698431365
transform -1 0 40768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__A1
timestamp 1698431365
transform 1 0 36848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__A2
timestamp 1698431365
transform 1 0 51296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2202__I
timestamp 1698431365
transform -1 0 48496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2207__A2
timestamp 1698431365
transform 1 0 51744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2212__A1
timestamp 1698431365
transform -1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2212__B2
timestamp 1698431365
transform -1 0 47936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__A1
timestamp 1698431365
transform 1 0 44912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2226__A1
timestamp 1698431365
transform -1 0 54208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2227__I
timestamp 1698431365
transform 1 0 38304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2234__A1
timestamp 1698431365
transform 1 0 51968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__A2
timestamp 1698431365
transform 1 0 50176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2262__I
timestamp 1698431365
transform 1 0 42784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2263__A1
timestamp 1698431365
transform -1 0 43680 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2264__A1
timestamp 1698431365
transform -1 0 46144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__A1
timestamp 1698431365
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__A2
timestamp 1698431365
transform -1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2272__A1
timestamp 1698431365
transform 1 0 38304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2272__A2
timestamp 1698431365
transform 1 0 39312 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2274__I
timestamp 1698431365
transform -1 0 34944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2276__A1
timestamp 1698431365
transform 1 0 42112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2276__A2
timestamp 1698431365
transform -1 0 41888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2283__A1
timestamp 1698431365
transform 1 0 47936 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2284__A1
timestamp 1698431365
transform 1 0 48160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__A1
timestamp 1698431365
transform -1 0 35616 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__A2
timestamp 1698431365
transform 1 0 35840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2293__A2
timestamp 1698431365
transform 1 0 40992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2294__A1
timestamp 1698431365
transform -1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A1
timestamp 1698431365
transform 1 0 50176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2298__A1
timestamp 1698431365
transform 1 0 46928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2305__A1
timestamp 1698431365
transform -1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2309__A2
timestamp 1698431365
transform 1 0 58128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2310__A2
timestamp 1698431365
transform -1 0 27216 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2311__A1
timestamp 1698431365
transform -1 0 30576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2313__A1
timestamp 1698431365
transform -1 0 27664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2314__A1
timestamp 1698431365
transform -1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2314__A2
timestamp 1698431365
transform -1 0 30128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__A2
timestamp 1698431365
transform 1 0 58016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2319__A1
timestamp 1698431365
transform 1 0 58128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__A1
timestamp 1698431365
transform 1 0 39872 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2346__A1
timestamp 1698431365
transform 1 0 48832 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2347__A1
timestamp 1698431365
transform 1 0 47712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2354__A1
timestamp 1698431365
transform 1 0 26544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2354__A2
timestamp 1698431365
transform -1 0 28896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2357__A1
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2357__A2
timestamp 1698431365
transform 1 0 27664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A2
timestamp 1698431365
transform -1 0 55552 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2369__A1
timestamp 1698431365
transform -1 0 35504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2369__A2
timestamp 1698431365
transform -1 0 35392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2370__A2
timestamp 1698431365
transform 1 0 30576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2371__A1
timestamp 1698431365
transform 1 0 37408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2373__A1
timestamp 1698431365
transform -1 0 34720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2373__A2
timestamp 1698431365
transform 1 0 33936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2376__I
timestamp 1698431365
transform -1 0 31696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__A1
timestamp 1698431365
transform 1 0 37184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__I
timestamp 1698431365
transform 1 0 15008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2392__A1
timestamp 1698431365
transform -1 0 34608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2392__A2
timestamp 1698431365
transform 1 0 35728 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2393__I
timestamp 1698431365
transform 1 0 17136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2400__A1
timestamp 1698431365
transform 1 0 50848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2401__B
timestamp 1698431365
transform 1 0 30912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2402__A3
timestamp 1698431365
transform -1 0 30576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2403__A1
timestamp 1698431365
transform -1 0 31024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2405__I
timestamp 1698431365
transform 1 0 20832 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2408__A1
timestamp 1698431365
transform -1 0 43344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2408__B
timestamp 1698431365
transform 1 0 47152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__A1
timestamp 1698431365
transform -1 0 25872 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2424__A1
timestamp 1698431365
transform -1 0 31136 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2424__A2
timestamp 1698431365
transform 1 0 31360 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2425__A1
timestamp 1698431365
transform 1 0 34720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2425__A2
timestamp 1698431365
transform 1 0 34384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2434__A1
timestamp 1698431365
transform -1 0 22064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__A1
timestamp 1698431365
transform 1 0 24752 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__A1
timestamp 1698431365
transform 1 0 29232 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A1
timestamp 1698431365
transform -1 0 32480 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__A1
timestamp 1698431365
transform 1 0 17920 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__A2
timestamp 1698431365
transform -1 0 21504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__I
timestamp 1698431365
transform 1 0 16352 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A1
timestamp 1698431365
transform 1 0 17584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2446__A2
timestamp 1698431365
transform 1 0 20720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__A1
timestamp 1698431365
transform -1 0 20272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2450__A1
timestamp 1698431365
transform 1 0 30576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__A1
timestamp 1698431365
transform 1 0 17248 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__A2
timestamp 1698431365
transform -1 0 17920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2468__A2
timestamp 1698431365
transform -1 0 21616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__A1
timestamp 1698431365
transform 1 0 20160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2474__A1
timestamp 1698431365
transform -1 0 25648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2474__A2
timestamp 1698431365
transform 1 0 25760 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2493__A1
timestamp 1698431365
transform 1 0 18032 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A2
timestamp 1698431365
transform 1 0 22288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2512__A1
timestamp 1698431365
transform 1 0 17024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__I
timestamp 1698431365
transform 1 0 56000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2517__I
timestamp 1698431365
transform -1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__I
timestamp 1698431365
transform 1 0 11312 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__A2
timestamp 1698431365
transform 1 0 34608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A3
timestamp 1698431365
transform 1 0 11984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A4
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2521__A1
timestamp 1698431365
transform -1 0 7616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2524__C
timestamp 1698431365
transform -1 0 10304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2525__A1
timestamp 1698431365
transform -1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__C
timestamp 1698431365
transform -1 0 9856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2527__A1
timestamp 1698431365
transform 1 0 13888 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2527__A2
timestamp 1698431365
transform 1 0 13664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2528__A1
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2528__A2
timestamp 1698431365
transform -1 0 5936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__A1
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__I
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2542__A1
timestamp 1698431365
transform -1 0 3808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__C
timestamp 1698431365
transform 1 0 4032 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__A1
timestamp 1698431365
transform -1 0 2352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__A1
timestamp 1698431365
transform -1 0 2576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2550__A1
timestamp 1698431365
transform -1 0 4592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2552__A1
timestamp 1698431365
transform 1 0 5152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__A1
timestamp 1698431365
transform 1 0 10192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2557__A1
timestamp 1698431365
transform -1 0 7392 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2559__A1
timestamp 1698431365
transform -1 0 8848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2559__C
timestamp 1698431365
transform -1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__A2
timestamp 1698431365
transform 1 0 33712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__I
timestamp 1698431365
transform 1 0 8512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__C
timestamp 1698431365
transform -1 0 7280 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2566__I
timestamp 1698431365
transform 1 0 9744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2567__A1
timestamp 1698431365
transform 1 0 9072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2570__A1
timestamp 1698431365
transform -1 0 11648 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__A1
timestamp 1698431365
transform -1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__C
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__A1
timestamp 1698431365
transform 1 0 15008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__A1
timestamp 1698431365
transform -1 0 15680 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__C
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__A1
timestamp 1698431365
transform -1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__A1
timestamp 1698431365
transform 1 0 14336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__A1
timestamp 1698431365
transform 1 0 16352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__A1
timestamp 1698431365
transform 1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__C
timestamp 1698431365
transform 1 0 17024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__A1
timestamp 1698431365
transform 1 0 14112 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__A1
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__C
timestamp 1698431365
transform 1 0 14560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__A1
timestamp 1698431365
transform 1 0 15456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__A1
timestamp 1698431365
transform -1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__C
timestamp 1698431365
transform 1 0 15904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2587__A1
timestamp 1698431365
transform -1 0 11536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__A1
timestamp 1698431365
transform -1 0 13776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__A1
timestamp 1698431365
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__I
timestamp 1698431365
transform -1 0 8176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2594__A3
timestamp 1698431365
transform -1 0 10416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__C
timestamp 1698431365
transform -1 0 3808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__A1
timestamp 1698431365
transform 1 0 5152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__I
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__A1
timestamp 1698431365
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__A1
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__A1
timestamp 1698431365
transform 1 0 8512 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2623__I
timestamp 1698431365
transform -1 0 9968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__A2
timestamp 1698431365
transform 1 0 35728 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__A1
timestamp 1698431365
transform 1 0 18928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2631__I
timestamp 1698431365
transform 1 0 36288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__A2
timestamp 1698431365
transform 1 0 38416 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2633__A2
timestamp 1698431365
transform 1 0 38864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__A1
timestamp 1698431365
transform 1 0 15680 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__A2
timestamp 1698431365
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2636__A2
timestamp 1698431365
transform 1 0 38752 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__A1
timestamp 1698431365
transform 1 0 15456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__A2
timestamp 1698431365
transform 1 0 38304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__A2
timestamp 1698431365
transform 1 0 39648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__A1
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__A2
timestamp 1698431365
transform -1 0 35728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2643__A1
timestamp 1698431365
transform 1 0 12432 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__A1
timestamp 1698431365
transform 1 0 9968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2646__I
timestamp 1698431365
transform 1 0 9968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__A1
timestamp 1698431365
transform -1 0 12768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__A1
timestamp 1698431365
transform 1 0 9744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__A1
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2655__A1
timestamp 1698431365
transform 1 0 9408 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__C
timestamp 1698431365
transform 1 0 5040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__I
timestamp 1698431365
transform 1 0 4704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2675__A1
timestamp 1698431365
transform -1 0 4704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2677__A2
timestamp 1698431365
transform 1 0 10640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__A1
timestamp 1698431365
transform 1 0 11088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__B
timestamp 1698431365
transform 1 0 10304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2681__A2
timestamp 1698431365
transform 1 0 7168 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__A1
timestamp 1698431365
transform 1 0 7168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2683__B
timestamp 1698431365
transform -1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2684__A2
timestamp 1698431365
transform 1 0 9856 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__A1
timestamp 1698431365
transform -1 0 5936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2686__B
timestamp 1698431365
transform 1 0 8848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__A1
timestamp 1698431365
transform 1 0 16800 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__A1
timestamp 1698431365
transform -1 0 18816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__C
timestamp 1698431365
transform 1 0 17248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__A1
timestamp 1698431365
transform -1 0 19488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__A1
timestamp 1698431365
transform 1 0 9744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__B
timestamp 1698431365
transform 1 0 10640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__A1
timestamp 1698431365
transform -1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__A1
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__A1
timestamp 1698431365
transform 1 0 16688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2702__A1
timestamp 1698431365
transform 1 0 12320 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__A1
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__A1
timestamp 1698431365
transform 1 0 13328 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__A1
timestamp 1698431365
transform 1 0 13664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2708__C
timestamp 1698431365
transform 1 0 20160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__A1
timestamp 1698431365
transform 1 0 12544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__A1
timestamp 1698431365
transform -1 0 16464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__A1
timestamp 1698431365
transform 1 0 10192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2714__B
timestamp 1698431365
transform -1 0 10416 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2717__CLK
timestamp 1698431365
transform 1 0 51408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2718__CLK
timestamp 1698431365
transform 1 0 32144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2719__CLK
timestamp 1698431365
transform 1 0 30128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2720__CLK
timestamp 1698431365
transform 1 0 26656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2721__CLK
timestamp 1698431365
transform 1 0 24640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2722__CLK
timestamp 1698431365
transform 1 0 18480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2723__CLK
timestamp 1698431365
transform 1 0 14336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2725__CLK
timestamp 1698431365
transform 1 0 14896 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__CLK
timestamp 1698431365
transform 1 0 16128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__CLK
timestamp 1698431365
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2728__CLK
timestamp 1698431365
transform 1 0 11872 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2729__CLK
timestamp 1698431365
transform 1 0 11088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2730__CLK
timestamp 1698431365
transform 1 0 5040 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__CLK
timestamp 1698431365
transform 1 0 13664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__CLK
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__CLK
timestamp 1698431365
transform 1 0 7280 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__CLK
timestamp 1698431365
transform 1 0 6384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__CLK
timestamp 1698431365
transform 1 0 12432 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__CLK
timestamp 1698431365
transform 1 0 4368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2737__CLK
timestamp 1698431365
transform -1 0 6384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2738__CLK
timestamp 1698431365
transform -1 0 7280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2739__CLK
timestamp 1698431365
transform 1 0 35056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2740__CLK
timestamp 1698431365
transform 1 0 11984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2741__CLK
timestamp 1698431365
transform 1 0 3920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2742__CLK
timestamp 1698431365
transform 1 0 20384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2744__CLK
timestamp 1698431365
transform 1 0 4816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2760__CLK
timestamp 1698431365
transform 1 0 5712 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2791__CLK
timestamp 1698431365
transform 1 0 9408 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform -1 0 30352 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout54_I
timestamp 1698431365
transform 1 0 1904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout55_I
timestamp 1698431365
transform -1 0 6832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout63_I
timestamp 1698431365
transform -1 0 2016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout66_I
timestamp 1698431365
transform -1 0 2016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout67_I
timestamp 1698431365
transform -1 0 10080 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout72_I
timestamp 1698431365
transform -1 0 5040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout73_I
timestamp 1698431365
transform 1 0 35616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout74_I
timestamp 1698431365
transform 1 0 20272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 2800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 5936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 47040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 52080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 8960 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 11984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 6384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 3136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 11536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 6160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 6608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 3472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 5824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 8848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 6608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 6160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 6608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 5040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 7056 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 2688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 35056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 34160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 37856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 7728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 11984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 56000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 56896 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 56448 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 55552 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 51296 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 42896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 43008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 41664 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output37_I
timestamp 1698431365
transform 1 0 56560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_rebuffer2_I
timestamp 1698431365
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698431365
transform -1 0 26768 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698431365
transform -1 0 27552 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout54
timestamp 1698431365
transform 1 0 2576 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout55
timestamp 1698431365
transform 1 0 8512 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout56
timestamp 1698431365
transform -1 0 2352 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout57
timestamp 1698431365
transform -1 0 12320 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout58
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout59
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout60
timestamp 1698431365
transform 1 0 5040 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout61
timestamp 1698431365
transform 1 0 4368 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout62
timestamp 1698431365
transform -1 0 2688 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout63
timestamp 1698431365
transform 1 0 1792 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout64
timestamp 1698431365
transform -1 0 2240 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout65
timestamp 1698431365
transform -1 0 5152 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout66
timestamp 1698431365
transform 1 0 2016 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout67
timestamp 1698431365
transform -1 0 11648 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout68
timestamp 1698431365
transform -1 0 2688 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout69
timestamp 1698431365
transform 1 0 13888 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout70
timestamp 1698431365
transform 1 0 13888 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout71
timestamp 1698431365
transform -1 0 2800 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout72
timestamp 1698431365
transform 1 0 3248 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout73
timestamp 1698431365
transform 1 0 35840 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout74
timestamp 1698431365
transform -1 0 21168 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout75
timestamp 1698431365
transform 1 0 2576 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_10 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_19
timestamp 1698431365
transform 1 0 3472 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_27
timestamp 1698431365
transform 1 0 4368 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_38
timestamp 1698431365
transform 1 0 5600 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_41
timestamp 1698431365
transform 1 0 5936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_45
timestamp 1698431365
transform 1 0 6384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_49
timestamp 1698431365
transform 1 0 6832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_53
timestamp 1698431365
transform 1 0 7280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_63
timestamp 1698431365
transform 1 0 8400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_65
timestamp 1698431365
transform 1 0 8624 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_99
timestamp 1698431365
transform 1 0 12432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_167
timestamp 1698431365
transform 1 0 20048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_184
timestamp 1698431365
transform 1 0 21952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_208
timestamp 1698431365
transform 1 0 24640 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_269
timestamp 1698431365
transform 1 0 31472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698431365
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_276
timestamp 1698431365
transform 1 0 32256 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_283
timestamp 1698431365
transform 1 0 33040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_287
timestamp 1698431365
transform 1 0 33488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_291
timestamp 1698431365
transform 1 0 33936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_295
timestamp 1698431365
transform 1 0 34384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_299
timestamp 1698431365
transform 1 0 34832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_303
timestamp 1698431365
transform 1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_316 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_336
timestamp 1698431365
transform 1 0 38976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_350
timestamp 1698431365
transform 1 0 40544 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_370
timestamp 1698431365
transform 1 0 42784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_381
timestamp 1698431365
transform 1 0 44016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_385
timestamp 1698431365
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_400
timestamp 1698431365
transform 1 0 46144 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_420 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48384 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_436
timestamp 1698431365
transform 1 0 50176 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_440
timestamp 1698431365
transform 1 0 50624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_448
timestamp 1698431365
transform 1 0 51520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_450
timestamp 1698431365
transform 1 0 51744 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_461
timestamp 1698431365
transform 1 0 52976 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_469
timestamp 1698431365
transform 1 0 53872 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_473
timestamp 1698431365
transform 1 0 54320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_475
timestamp 1698431365
transform 1 0 54544 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_486
timestamp 1698431365
transform 1 0 55776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_490
timestamp 1698431365
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_492
timestamp 1698431365
transform 1 0 56448 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_505
timestamp 1698431365
transform 1 0 57904 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_18
timestamp 1698431365
transform 1 0 3360 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_22
timestamp 1698431365
transform 1 0 3808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_24
timestamp 1698431365
transform 1 0 4032 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_54
timestamp 1698431365
transform 1 0 7392 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_65
timestamp 1698431365
transform 1 0 8624 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_74
timestamp 1698431365
transform 1 0 9632 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_172
timestamp 1698431365
transform 1 0 20608 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_218
timestamp 1698431365
transform 1 0 25760 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_295
timestamp 1698431365
transform 1 0 34384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_299
timestamp 1698431365
transform 1 0 34832 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_303
timestamp 1698431365
transform 1 0 35280 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_319
timestamp 1698431365
transform 1 0 37072 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_323
timestamp 1698431365
transform 1 0 37520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_325
timestamp 1698431365
transform 1 0 37744 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_341
timestamp 1698431365
transform 1 0 39536 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_376
timestamp 1698431365
transform 1 0 43456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_406
timestamp 1698431365
transform 1 0 46816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_418
timestamp 1698431365
transform 1 0 48160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_438
timestamp 1698431365
transform 1 0 50400 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_446
timestamp 1698431365
transform 1 0 51296 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_456 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 52416 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_488
timestamp 1698431365
transform 1 0 56000 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_508
timestamp 1698431365
transform 1 0 58240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_18
timestamp 1698431365
transform 1 0 3360 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_21
timestamp 1698431365
transform 1 0 3696 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_25
timestamp 1698431365
transform 1 0 4144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_64
timestamp 1698431365
transform 1 0 8512 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_91
timestamp 1698431365
transform 1 0 11536 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_97
timestamp 1698431365
transform 1 0 12208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_130
timestamp 1698431365
transform 1 0 15904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_132
timestamp 1698431365
transform 1 0 16128 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_179
timestamp 1698431365
transform 1 0 21392 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_238
timestamp 1698431365
transform 1 0 28000 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_299
timestamp 1698431365
transform 1 0 34832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_303
timestamp 1698431365
transform 1 0 35280 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_312
timestamp 1698431365
transform 1 0 36288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698431365
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_340
timestamp 1698431365
transform 1 0 39424 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_358
timestamp 1698431365
transform 1 0 41440 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_371
timestamp 1698431365
transform 1 0 42896 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_393
timestamp 1698431365
transform 1 0 45360 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_401
timestamp 1698431365
transform 1 0 46256 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_419
timestamp 1698431365
transform 1 0 48272 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_434
timestamp 1698431365
transform 1 0 49952 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_475
timestamp 1698431365
transform 1 0 54544 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_503
timestamp 1698431365
transform 1 0 57680 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_507
timestamp 1698431365
transform 1 0 58128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_4
timestamp 1698431365
transform 1 0 1792 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_7
timestamp 1698431365
transform 1 0 2128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_76
timestamp 1698431365
transform 1 0 9856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_91
timestamp 1698431365
transform 1 0 11536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_93
timestamp 1698431365
transform 1 0 11760 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_115
timestamp 1698431365
transform 1 0 14224 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_167
timestamp 1698431365
transform 1 0 20048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_228
timestamp 1698431365
transform 1 0 26880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_287
timestamp 1698431365
transform 1 0 33488 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_323
timestamp 1698431365
transform 1 0 37520 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_325
timestamp 1698431365
transform 1 0 37744 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_338
timestamp 1698431365
transform 1 0 39200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_340
timestamp 1698431365
transform 1 0 39424 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698431365
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_411
timestamp 1698431365
transform 1 0 47376 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_479
timestamp 1698431365
transform 1 0 54992 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_483
timestamp 1698431365
transform 1 0 55440 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1698431365
transform 1 0 4928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_51
timestamp 1698431365
transform 1 0 7056 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_53
timestamp 1698431365
transform 1 0 7280 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_87
timestamp 1698431365
transform 1 0 11088 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_91
timestamp 1698431365
transform 1 0 11536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_119
timestamp 1698431365
transform 1 0 14672 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_121
timestamp 1698431365
transform 1 0 14896 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_234
timestamp 1698431365
transform 1 0 27552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_236
timestamp 1698431365
transform 1 0 27776 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_289
timestamp 1698431365
transform 1 0 33712 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_295
timestamp 1698431365
transform 1 0 34384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_297
timestamp 1698431365
transform 1 0 34608 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_314
timestamp 1698431365
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_321
timestamp 1698431365
transform 1 0 37296 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_369
timestamp 1698431365
transform 1 0 42672 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_384
timestamp 1698431365
transform 1 0 44352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_418
timestamp 1698431365
transform 1 0 48160 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_420
timestamp 1698431365
transform 1 0 48384 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_440
timestamp 1698431365
transform 1 0 50624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_444
timestamp 1698431365
transform 1 0 51072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_448
timestamp 1698431365
transform 1 0 51520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_452
timestamp 1698431365
transform 1 0 51968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_454
timestamp 1698431365
transform 1 0 52192 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_474
timestamp 1698431365
transform 1 0 54432 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_482
timestamp 1698431365
transform 1 0 55328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_6
timestamp 1698431365
transform 1 0 2016 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_25
timestamp 1698431365
transform 1 0 4144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_29
timestamp 1698431365
transform 1 0 4592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_33
timestamp 1698431365
transform 1 0 5040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_55
timestamp 1698431365
transform 1 0 7504 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_64
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_101
timestamp 1698431365
transform 1 0 12656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_115
timestamp 1698431365
transform 1 0 14224 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_251
timestamp 1698431365
transform 1 0 29456 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_298
timestamp 1698431365
transform 1 0 34720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_315
timestamp 1698431365
transform 1 0 36624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_319
timestamp 1698431365
transform 1 0 37072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_323
timestamp 1698431365
transform 1 0 37520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_327
timestamp 1698431365
transform 1 0 37968 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_349
timestamp 1698431365
transform 1 0 40432 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_391
timestamp 1698431365
transform 1 0 45136 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_395
timestamp 1698431365
transform 1 0 45584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_409
timestamp 1698431365
transform 1 0 47152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_444
timestamp 1698431365
transform 1 0 51072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_482
timestamp 1698431365
transform 1 0 55328 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_506
timestamp 1698431365
transform 1 0 58016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_31
timestamp 1698431365
transform 1 0 4816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_60
timestamp 1698431365
transform 1 0 8064 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_64
timestamp 1698431365
transform 1 0 8512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_96
timestamp 1698431365
transform 1 0 12096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_149
timestamp 1698431365
transform 1 0 18032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_199
timestamp 1698431365
transform 1 0 23632 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_226
timestamp 1698431365
transform 1 0 26656 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_269
timestamp 1698431365
transform 1 0 31472 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_271
timestamp 1698431365
transform 1 0 31696 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_312
timestamp 1698431365
transform 1 0 36288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698431365
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_382
timestamp 1698431365
transform 1 0 44128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_384
timestamp 1698431365
transform 1 0 44352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_415
timestamp 1698431365
transform 1 0 47824 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_442
timestamp 1698431365
transform 1 0 50848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_450
timestamp 1698431365
transform 1 0 51744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_454
timestamp 1698431365
transform 1 0 52192 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_461
timestamp 1698431365
transform 1 0 52976 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_468
timestamp 1698431365
transform 1 0 53760 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_9
timestamp 1698431365
transform 1 0 2352 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_17
timestamp 1698431365
transform 1 0 3248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_19
timestamp 1698431365
transform 1 0 3472 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_22
timestamp 1698431365
transform 1 0 3808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_26
timestamp 1698431365
transform 1 0 4256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_30
timestamp 1698431365
transform 1 0 4704 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_33
timestamp 1698431365
transform 1 0 5040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_129
timestamp 1698431365
transform 1 0 15792 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_131
timestamp 1698431365
transform 1 0 16016 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_183
timestamp 1698431365
transform 1 0 21840 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_214
timestamp 1698431365
transform 1 0 25312 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_230
timestamp 1698431365
transform 1 0 27104 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_263
timestamp 1698431365
transform 1 0 30800 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_272
timestamp 1698431365
transform 1 0 31808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_291
timestamp 1698431365
transform 1 0 33936 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_293
timestamp 1698431365
transform 1 0 34160 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_302
timestamp 1698431365
transform 1 0 35168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_337
timestamp 1698431365
transform 1 0 39088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_347
timestamp 1698431365
transform 1 0 40208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_349
timestamp 1698431365
transform 1 0 40432 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_358
timestamp 1698431365
transform 1 0 41440 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_376
timestamp 1698431365
transform 1 0 43456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_383
timestamp 1698431365
transform 1 0 44240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_387
timestamp 1698431365
transform 1 0 44688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_405
timestamp 1698431365
transform 1 0 46704 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_419
timestamp 1698431365
transform 1 0 48272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_437
timestamp 1698431365
transform 1 0 50288 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_441
timestamp 1698431365
transform 1 0 50736 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_473
timestamp 1698431365
transform 1 0 54320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_475
timestamp 1698431365
transform 1 0 54544 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_489
timestamp 1698431365
transform 1 0 56112 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_505
timestamp 1698431365
transform 1 0 57904 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_31
timestamp 1698431365
transform 1 0 4816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_39
timestamp 1698431365
transform 1 0 5712 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_92
timestamp 1698431365
transform 1 0 11648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_94
timestamp 1698431365
transform 1 0 11872 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_97
timestamp 1698431365
transform 1 0 12208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_131
timestamp 1698431365
transform 1 0 16016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_133
timestamp 1698431365
transform 1 0 16240 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_165
timestamp 1698431365
transform 1 0 19824 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_286
timestamp 1698431365
transform 1 0 33376 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_309
timestamp 1698431365
transform 1 0 35952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_329
timestamp 1698431365
transform 1 0 38192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_383
timestamp 1698431365
transform 1 0 44240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_416
timestamp 1698431365
transform 1 0 47936 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_446
timestamp 1698431365
transform 1 0 51296 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_454
timestamp 1698431365
transform 1 0 52192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_465
timestamp 1698431365
transform 1 0 53424 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_473
timestamp 1698431365
transform 1 0 54320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_8
timestamp 1698431365
transform 1 0 2240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_65
timestamp 1698431365
transform 1 0 8624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_67
timestamp 1698431365
transform 1 0 8848 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_74
timestamp 1698431365
transform 1 0 9632 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_126
timestamp 1698431365
transform 1 0 15456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_132
timestamp 1698431365
transform 1 0 16128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_157
timestamp 1698431365
transform 1 0 18928 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_208
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_217
timestamp 1698431365
transform 1 0 25648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_247
timestamp 1698431365
transform 1 0 29008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_249
timestamp 1698431365
transform 1 0 29232 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_268
timestamp 1698431365
transform 1 0 31360 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_270
timestamp 1698431365
transform 1 0 31584 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_273
timestamp 1698431365
transform 1 0 31920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_277
timestamp 1698431365
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_288
timestamp 1698431365
transform 1 0 33600 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_292
timestamp 1698431365
transform 1 0 34048 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_322
timestamp 1698431365
transform 1 0 37408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_330
timestamp 1698431365
transform 1 0 38304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_334
timestamp 1698431365
transform 1 0 38752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_394
timestamp 1698431365
transform 1 0 45472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_410
timestamp 1698431365
transform 1 0 47264 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_418
timestamp 1698431365
transform 1 0 48160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_435
timestamp 1698431365
transform 1 0 50064 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_439
timestamp 1698431365
transform 1 0 50512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_441
timestamp 1698431365
transform 1 0 50736 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_454
timestamp 1698431365
transform 1 0 52192 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_462
timestamp 1698431365
transform 1 0 53088 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_466
timestamp 1698431365
transform 1 0 53536 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_504
timestamp 1698431365
transform 1 0 57792 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698431365
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_77
timestamp 1698431365
transform 1 0 9968 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_113
timestamp 1698431365
transform 1 0 14000 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_143
timestamp 1698431365
transform 1 0 17360 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_145
timestamp 1698431365
transform 1 0 17584 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_208
timestamp 1698431365
transform 1 0 24640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_210
timestamp 1698431365
transform 1 0 24864 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_249
timestamp 1698431365
transform 1 0 29232 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_299
timestamp 1698431365
transform 1 0 34832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_358
timestamp 1698431365
transform 1 0 41440 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_362
timestamp 1698431365
transform 1 0 41888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_366
timestamp 1698431365
transform 1 0 42336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_370
timestamp 1698431365
transform 1 0 42784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_374
timestamp 1698431365
transform 1 0 43232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_378
timestamp 1698431365
transform 1 0 43680 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_382
timestamp 1698431365
transform 1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_389
timestamp 1698431365
transform 1 0 44912 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_400
timestamp 1698431365
transform 1 0 46144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_402
timestamp 1698431365
transform 1 0 46368 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_423
timestamp 1698431365
transform 1 0 48720 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_427
timestamp 1698431365
transform 1 0 49168 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_446
timestamp 1698431365
transform 1 0 51296 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_453
timestamp 1698431365
transform 1 0 52080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_473
timestamp 1698431365
transform 1 0 54320 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_39
timestamp 1698431365
transform 1 0 5712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_64
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_78
timestamp 1698431365
transform 1 0 10080 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_86
timestamp 1698431365
transform 1 0 10976 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_121
timestamp 1698431365
transform 1 0 14896 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_125
timestamp 1698431365
transform 1 0 15344 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_152
timestamp 1698431365
transform 1 0 18368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_154
timestamp 1698431365
transform 1 0 18592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_186
timestamp 1698431365
transform 1 0 22176 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_244
timestamp 1698431365
transform 1 0 28672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_248
timestamp 1698431365
transform 1 0 29120 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_252
timestamp 1698431365
transform 1 0 29568 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_277
timestamp 1698431365
transform 1 0 32368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_293
timestamp 1698431365
transform 1 0 34160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_297
timestamp 1698431365
transform 1 0 34608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_301
timestamp 1698431365
transform 1 0 35056 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_305
timestamp 1698431365
transform 1 0 35504 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_307
timestamp 1698431365
transform 1 0 35728 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_328
timestamp 1698431365
transform 1 0 38080 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_336
timestamp 1698431365
transform 1 0 38976 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_376
timestamp 1698431365
transform 1 0 43456 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_412
timestamp 1698431365
transform 1 0 47488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_450
timestamp 1698431365
transform 1 0 51744 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_503
timestamp 1698431365
transform 1 0 57680 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_507
timestamp 1698431365
transform 1 0 58128 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_4
timestamp 1698431365
transform 1 0 1792 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_41
timestamp 1698431365
transform 1 0 5936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_113
timestamp 1698431365
transform 1 0 14000 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_117
timestamp 1698431365
transform 1 0 14448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_131
timestamp 1698431365
transform 1 0 16016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_162
timestamp 1698431365
transform 1 0 19488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_164
timestamp 1698431365
transform 1 0 19712 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_170
timestamp 1698431365
transform 1 0 20384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_172
timestamp 1698431365
transform 1 0 20608 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_181
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_184
timestamp 1698431365
transform 1 0 21952 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_188
timestamp 1698431365
transform 1 0 22400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_235
timestamp 1698431365
transform 1 0 27664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_239
timestamp 1698431365
transform 1 0 28112 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_268
timestamp 1698431365
transform 1 0 31360 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_272
timestamp 1698431365
transform 1 0 31808 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_308
timestamp 1698431365
transform 1 0 35840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_312
timestamp 1698431365
transform 1 0 36288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_362
timestamp 1698431365
transform 1 0 41888 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_370
timestamp 1698431365
transform 1 0 42784 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_374
timestamp 1698431365
transform 1 0 43232 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_376
timestamp 1698431365
transform 1 0 43456 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_403
timestamp 1698431365
transform 1 0 46480 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_428
timestamp 1698431365
transform 1 0 49280 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_442
timestamp 1698431365
transform 1 0 50848 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_473
timestamp 1698431365
transform 1 0 54320 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_4
timestamp 1698431365
transform 1 0 1792 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_50
timestamp 1698431365
transform 1 0 6944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_54
timestamp 1698431365
transform 1 0 7392 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_87
timestamp 1698431365
transform 1 0 11088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_89
timestamp 1698431365
transform 1 0 11312 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_111
timestamp 1698431365
transform 1 0 13776 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_152
timestamp 1698431365
transform 1 0 18368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_156
timestamp 1698431365
transform 1 0 18816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_160
timestamp 1698431365
transform 1 0 19264 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_162
timestamp 1698431365
transform 1 0 19488 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_165
timestamp 1698431365
transform 1 0 19824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_169
timestamp 1698431365
transform 1 0 20272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_173
timestamp 1698431365
transform 1 0 20720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_203
timestamp 1698431365
transform 1 0 24080 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_207
timestamp 1698431365
transform 1 0 24528 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_226
timestamp 1698431365
transform 1 0 26656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_230
timestamp 1698431365
transform 1 0 27104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_234
timestamp 1698431365
transform 1 0 27552 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_266
timestamp 1698431365
transform 1 0 31136 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_298
timestamp 1698431365
transform 1 0 34720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_302
timestamp 1698431365
transform 1 0 35168 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_308
timestamp 1698431365
transform 1 0 35840 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_325
timestamp 1698431365
transform 1 0 37744 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_341
timestamp 1698431365
transform 1 0 39536 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_381
timestamp 1698431365
transform 1 0 44016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_417
timestamp 1698431365
transform 1 0 48048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_419
timestamp 1698431365
transform 1 0 48272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_435
timestamp 1698431365
transform 1 0 50064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_439
timestamp 1698431365
transform 1 0 50512 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_484
timestamp 1698431365
transform 1 0 55552 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_507
timestamp 1698431365
transform 1 0 58128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_43
timestamp 1698431365
transform 1 0 6160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_47
timestamp 1698431365
transform 1 0 6608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_51
timestamp 1698431365
transform 1 0 7056 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_93
timestamp 1698431365
transform 1 0 11760 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_95
timestamp 1698431365
transform 1 0 11984 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_109
timestamp 1698431365
transform 1 0 13552 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_112
timestamp 1698431365
transform 1 0 13888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_116
timestamp 1698431365
transform 1 0 14336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_138
timestamp 1698431365
transform 1 0 16800 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_142
timestamp 1698431365
transform 1 0 17248 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_194
timestamp 1698431365
transform 1 0 23072 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_220
timestamp 1698431365
transform 1 0 25984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_222
timestamp 1698431365
transform 1 0 26208 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_229
timestamp 1698431365
transform 1 0 26992 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_233
timestamp 1698431365
transform 1 0 27440 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_260
timestamp 1698431365
transform 1 0 30464 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_268
timestamp 1698431365
transform 1 0 31360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_276
timestamp 1698431365
transform 1 0 32256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_280
timestamp 1698431365
transform 1 0 32704 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_294
timestamp 1698431365
transform 1 0 34272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_296
timestamp 1698431365
transform 1 0 34496 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_321
timestamp 1698431365
transform 1 0 37296 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_329
timestamp 1698431365
transform 1 0 38192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_349
timestamp 1698431365
transform 1 0 40432 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_366
timestamp 1698431365
transform 1 0 42336 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_374
timestamp 1698431365
transform 1 0 43232 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_378
timestamp 1698431365
transform 1 0 43680 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_395
timestamp 1698431365
transform 1 0 45584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_397
timestamp 1698431365
transform 1 0 45808 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_414
timestamp 1698431365
transform 1 0 47712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_427
timestamp 1698431365
transform 1 0 49168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_431
timestamp 1698431365
transform 1 0 49616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_435
timestamp 1698431365
transform 1 0 50064 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_439
timestamp 1698431365
transform 1 0 50512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_453
timestamp 1698431365
transform 1 0 52080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_465
timestamp 1698431365
transform 1 0 53424 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_473
timestamp 1698431365
transform 1 0 54320 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_481
timestamp 1698431365
transform 1 0 55216 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_31
timestamp 1698431365
transform 1 0 4816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_33
timestamp 1698431365
transform 1 0 5040 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_43
timestamp 1698431365
transform 1 0 6160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_63
timestamp 1698431365
transform 1 0 8400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_67
timestamp 1698431365
transform 1 0 8848 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_74
timestamp 1698431365
transform 1 0 9632 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_87
timestamp 1698431365
transform 1 0 11088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_120
timestamp 1698431365
transform 1 0 14784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_124
timestamp 1698431365
transform 1 0 15232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_128
timestamp 1698431365
transform 1 0 15680 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_132
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698431365
transform 1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_150
timestamp 1698431365
transform 1 0 18144 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_154
timestamp 1698431365
transform 1 0 18592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_156
timestamp 1698431365
transform 1 0 18816 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_159
timestamp 1698431365
transform 1 0 19152 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_167
timestamp 1698431365
transform 1 0 20048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_169
timestamp 1698431365
transform 1 0 20272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_189
timestamp 1698431365
transform 1 0 22512 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_217
timestamp 1698431365
transform 1 0 25648 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_235
timestamp 1698431365
transform 1 0 27664 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_260
timestamp 1698431365
transform 1 0 30464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_264
timestamp 1698431365
transform 1 0 30912 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_272
timestamp 1698431365
transform 1 0 31808 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698431365
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_286
timestamp 1698431365
transform 1 0 33376 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_305
timestamp 1698431365
transform 1 0 35504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_307
timestamp 1698431365
transform 1 0 35728 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_343
timestamp 1698431365
transform 1 0 39760 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_347
timestamp 1698431365
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_369
timestamp 1698431365
transform 1 0 42672 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_396
timestamp 1698431365
transform 1 0 45696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_398
timestamp 1698431365
transform 1 0 45920 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_409
timestamp 1698431365
transform 1 0 47152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_413
timestamp 1698431365
transform 1 0 47600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_505
timestamp 1698431365
transform 1 0 57904 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_31
timestamp 1698431365
transform 1 0 4816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_56
timestamp 1698431365
transform 1 0 7616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_58
timestamp 1698431365
transform 1 0 7840 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_73
timestamp 1698431365
transform 1 0 9520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_77
timestamp 1698431365
transform 1 0 9968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_87
timestamp 1698431365
transform 1 0 11088 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_111
timestamp 1698431365
transform 1 0 13776 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_114
timestamp 1698431365
transform 1 0 14112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_118
timestamp 1698431365
transform 1 0 14560 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_148
timestamp 1698431365
transform 1 0 17920 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_155
timestamp 1698431365
transform 1 0 18704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_159
timestamp 1698431365
transform 1 0 19152 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_165
timestamp 1698431365
transform 1 0 19824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_169
timestamp 1698431365
transform 1 0 20272 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_179
timestamp 1698431365
transform 1 0 21392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_203
timestamp 1698431365
transform 1 0 24080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_205
timestamp 1698431365
transform 1 0 24304 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_224
timestamp 1698431365
transform 1 0 26432 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_249
timestamp 1698431365
transform 1 0 29232 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_269
timestamp 1698431365
transform 1 0 31472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_293
timestamp 1698431365
transform 1 0 34160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_297
timestamp 1698431365
transform 1 0 34608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_301
timestamp 1698431365
transform 1 0 35056 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_305
timestamp 1698431365
transform 1 0 35504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_309
timestamp 1698431365
transform 1 0 35952 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_325
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_329
timestamp 1698431365
transform 1 0 38192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_333
timestamp 1698431365
transform 1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_337
timestamp 1698431365
transform 1 0 39088 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_339
timestamp 1698431365
transform 1 0 39312 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_346
timestamp 1698431365
transform 1 0 40096 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_350
timestamp 1698431365
transform 1 0 40544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_352
timestamp 1698431365
transform 1 0 40768 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_384
timestamp 1698431365
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_409
timestamp 1698431365
transform 1 0 47152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_413
timestamp 1698431365
transform 1 0 47600 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_440
timestamp 1698431365
transform 1 0 50624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_444
timestamp 1698431365
transform 1 0 51072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_448
timestamp 1698431365
transform 1 0 51520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_452
timestamp 1698431365
transform 1 0 51968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_454
timestamp 1698431365
transform 1 0 52192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_463
timestamp 1698431365
transform 1 0 53200 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_479
timestamp 1698431365
transform 1 0 54992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_43
timestamp 1698431365
transform 1 0 6160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_47
timestamp 1698431365
transform 1 0 6608 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_80
timestamp 1698431365
transform 1 0 10304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_82
timestamp 1698431365
transform 1 0 10528 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_97
timestamp 1698431365
transform 1 0 12208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_99
timestamp 1698431365
transform 1 0 12432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_110
timestamp 1698431365
transform 1 0 13664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_126
timestamp 1698431365
transform 1 0 15456 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_171
timestamp 1698431365
transform 1 0 20496 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_201
timestamp 1698431365
transform 1 0 23856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_225
timestamp 1698431365
transform 1 0 26544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_227
timestamp 1698431365
transform 1 0 26768 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_243
timestamp 1698431365
transform 1 0 28560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_245
timestamp 1698431365
transform 1 0 28784 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_263
timestamp 1698431365
transform 1 0 30800 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_269
timestamp 1698431365
transform 1 0 31472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_273
timestamp 1698431365
transform 1 0 31920 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_293
timestamp 1698431365
transform 1 0 34160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_303
timestamp 1698431365
transform 1 0 35280 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_359
timestamp 1698431365
transform 1 0 41552 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_363
timestamp 1698431365
transform 1 0 42000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_382
timestamp 1698431365
transform 1 0 44128 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_390
timestamp 1698431365
transform 1 0 45024 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_403
timestamp 1698431365
transform 1 0 46480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_405
timestamp 1698431365
transform 1 0 46704 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_417
timestamp 1698431365
transform 1 0 48048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_432
timestamp 1698431365
transform 1 0 49728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_436
timestamp 1698431365
transform 1 0 50176 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_440
timestamp 1698431365
transform 1 0 50624 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_453
timestamp 1698431365
transform 1 0 52080 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_455
timestamp 1698431365
transform 1 0 52304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_482
timestamp 1698431365
transform 1 0 55328 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_505
timestamp 1698431365
transform 1 0 57904 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_14
timestamp 1698431365
transform 1 0 2912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_18
timestamp 1698431365
transform 1 0 3360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_43
timestamp 1698431365
transform 1 0 6160 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_47
timestamp 1698431365
transform 1 0 6608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_59
timestamp 1698431365
transform 1 0 7952 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_63
timestamp 1698431365
transform 1 0 8400 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_66
timestamp 1698431365
transform 1 0 8736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_68
timestamp 1698431365
transform 1 0 8960 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_112
timestamp 1698431365
transform 1 0 13888 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_126
timestamp 1698431365
transform 1 0 15456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_139
timestamp 1698431365
transform 1 0 16912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_141
timestamp 1698431365
transform 1 0 17136 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_144
timestamp 1698431365
transform 1 0 17472 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_150
timestamp 1698431365
transform 1 0 18144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_152
timestamp 1698431365
transform 1 0 18368 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_165
timestamp 1698431365
transform 1 0 19824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_167
timestamp 1698431365
transform 1 0 20048 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_227
timestamp 1698431365
transform 1 0 26768 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_272
timestamp 1698431365
transform 1 0 31808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_274
timestamp 1698431365
transform 1 0 32032 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_287
timestamp 1698431365
transform 1 0 33488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_289
timestamp 1698431365
transform 1 0 33712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_350
timestamp 1698431365
transform 1 0 40544 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_354
timestamp 1698431365
transform 1 0 40992 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_393
timestamp 1698431365
transform 1 0 45360 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_399
timestamp 1698431365
transform 1 0 46032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_401
timestamp 1698431365
transform 1 0 46256 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_408
timestamp 1698431365
transform 1 0 47040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_410
timestamp 1698431365
transform 1 0 47264 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_417
timestamp 1698431365
transform 1 0 48048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_421
timestamp 1698431365
transform 1 0 48496 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_448
timestamp 1698431365
transform 1 0 51520 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_452
timestamp 1698431365
transform 1 0 51968 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_454
timestamp 1698431365
transform 1 0 52192 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_459
timestamp 1698431365
transform 1 0 52752 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_508
timestamp 1698431365
transform 1 0 58240 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_8
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_10
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_51
timestamp 1698431365
transform 1 0 7056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_86
timestamp 1698431365
transform 1 0 10976 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_97
timestamp 1698431365
transform 1 0 12208 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_99
timestamp 1698431365
transform 1 0 12432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_172
timestamp 1698431365
transform 1 0 20608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_174
timestamp 1698431365
transform 1 0 20832 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_201
timestamp 1698431365
transform 1 0 23856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_229
timestamp 1698431365
transform 1 0 26992 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_245
timestamp 1698431365
transform 1 0 28784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_302
timestamp 1698431365
transform 1 0 35168 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_306
timestamp 1698431365
transform 1 0 35616 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_310
timestamp 1698431365
transform 1 0 36064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_314
timestamp 1698431365
transform 1 0 36512 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_328
timestamp 1698431365
transform 1 0 38080 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_332
timestamp 1698431365
transform 1 0 38528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_336
timestamp 1698431365
transform 1 0 38976 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_344
timestamp 1698431365
transform 1 0 39872 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_356
timestamp 1698431365
transform 1 0 41216 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_371
timestamp 1698431365
transform 1 0 42896 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_375
timestamp 1698431365
transform 1 0 43344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_377
timestamp 1698431365
transform 1 0 43568 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_394
timestamp 1698431365
transform 1 0 45472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_398
timestamp 1698431365
transform 1 0 45920 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_417
timestamp 1698431365
transform 1 0 48048 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_419
timestamp 1698431365
transform 1 0 48272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_442
timestamp 1698431365
transform 1 0 50848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_469
timestamp 1698431365
transform 1 0 53872 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_505
timestamp 1698431365
transform 1 0 57904 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_31
timestamp 1698431365
transform 1 0 4816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_57
timestamp 1698431365
transform 1 0 7728 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_74
timestamp 1698431365
transform 1 0 9632 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_115
timestamp 1698431365
transform 1 0 14224 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_121
timestamp 1698431365
transform 1 0 14896 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_125
timestamp 1698431365
transform 1 0 15344 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_133
timestamp 1698431365
transform 1 0 16240 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_137
timestamp 1698431365
transform 1 0 16688 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_140
timestamp 1698431365
transform 1 0 17024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_149
timestamp 1698431365
transform 1 0 18032 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_153
timestamp 1698431365
transform 1 0 18480 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_204
timestamp 1698431365
transform 1 0 24192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_208
timestamp 1698431365
transform 1 0 24640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_212
timestamp 1698431365
transform 1 0 25088 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_226
timestamp 1698431365
transform 1 0 26656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_230
timestamp 1698431365
transform 1 0 27104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_232
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_255
timestamp 1698431365
transform 1 0 29904 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_259
timestamp 1698431365
transform 1 0 30352 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_275
timestamp 1698431365
transform 1 0 32144 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_299
timestamp 1698431365
transform 1 0 34832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_348
timestamp 1698431365
transform 1 0 40320 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_352
timestamp 1698431365
transform 1 0 40768 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_383
timestamp 1698431365
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_393
timestamp 1698431365
transform 1 0 45360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_419
timestamp 1698431365
transform 1 0 48272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_421
timestamp 1698431365
transform 1 0 48496 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_434
timestamp 1698431365
transform 1 0 49952 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_438
timestamp 1698431365
transform 1 0 50400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_445
timestamp 1698431365
transform 1 0 51184 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_471
timestamp 1698431365
transform 1 0 54096 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_475
timestamp 1698431365
transform 1 0 54544 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_505
timestamp 1698431365
transform 1 0 57904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_14
timestamp 1698431365
transform 1 0 2912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_25
timestamp 1698431365
transform 1 0 4144 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_41
timestamp 1698431365
transform 1 0 5936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_45
timestamp 1698431365
transform 1 0 6384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_49
timestamp 1698431365
transform 1 0 6832 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_53
timestamp 1698431365
transform 1 0 7280 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_57
timestamp 1698431365
transform 1 0 7728 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698431365
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_74
timestamp 1698431365
transform 1 0 9632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_77
timestamp 1698431365
transform 1 0 9968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_95
timestamp 1698431365
transform 1 0 11984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_105
timestamp 1698431365
transform 1 0 13104 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_155
timestamp 1698431365
transform 1 0 18704 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_166
timestamp 1698431365
transform 1 0 19936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_170
timestamp 1698431365
transform 1 0 20384 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_176
timestamp 1698431365
transform 1 0 21056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_178
timestamp 1698431365
transform 1 0 21280 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_203
timestamp 1698431365
transform 1 0 24080 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_262
timestamp 1698431365
transform 1 0 30688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_266
timestamp 1698431365
transform 1 0 31136 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_270
timestamp 1698431365
transform 1 0 31584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_286
timestamp 1698431365
transform 1 0 33376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_336
timestamp 1698431365
transform 1 0 38976 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_340
timestamp 1698431365
transform 1 0 39424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_344
timestamp 1698431365
transform 1 0 39872 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_348
timestamp 1698431365
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_357
timestamp 1698431365
transform 1 0 41328 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_411
timestamp 1698431365
transform 1 0 47376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_413
timestamp 1698431365
transform 1 0 47600 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_433
timestamp 1698431365
transform 1 0 49840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_440
timestamp 1698431365
transform 1 0 50624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_444
timestamp 1698431365
transform 1 0 51072 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_448
timestamp 1698431365
transform 1 0 51520 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_452
timestamp 1698431365
transform 1 0 51968 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_464
timestamp 1698431365
transform 1 0 53312 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_474
timestamp 1698431365
transform 1 0 54432 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_482
timestamp 1698431365
transform 1 0 55328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_484
timestamp 1698431365
transform 1 0 55552 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_504
timestamp 1698431365
transform 1 0 57792 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_508
timestamp 1698431365
transform 1 0 58240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_31
timestamp 1698431365
transform 1 0 4816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_74
timestamp 1698431365
transform 1 0 9632 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_82
timestamp 1698431365
transform 1 0 10528 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_99
timestamp 1698431365
transform 1 0 12432 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_103
timestamp 1698431365
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_109
timestamp 1698431365
transform 1 0 13552 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_126
timestamp 1698431365
transform 1 0 15456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_128
timestamp 1698431365
transform 1 0 15680 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_179
timestamp 1698431365
transform 1 0 21392 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_192
timestamp 1698431365
transform 1 0 22848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_194
timestamp 1698431365
transform 1 0 23072 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_293
timestamp 1698431365
transform 1 0 34160 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_297
timestamp 1698431365
transform 1 0 34608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_301
timestamp 1698431365
transform 1 0 35056 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_418
timestamp 1698431365
transform 1 0 48160 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_422
timestamp 1698431365
transform 1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_424
timestamp 1698431365
transform 1 0 48832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_434
timestamp 1698431365
transform 1 0 49952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_446
timestamp 1698431365
transform 1 0 51296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_450
timestamp 1698431365
transform 1 0 51744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_454
timestamp 1698431365
transform 1 0 52192 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_479
timestamp 1698431365
transform 1 0 54992 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_18
timestamp 1698431365
transform 1 0 3360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_20
timestamp 1698431365
transform 1 0 3584 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_33
timestamp 1698431365
transform 1 0 5040 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_49
timestamp 1698431365
transform 1 0 6832 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_53
timestamp 1698431365
transform 1 0 7280 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_74
timestamp 1698431365
transform 1 0 9632 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_109
timestamp 1698431365
transform 1 0 13552 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_111
timestamp 1698431365
transform 1 0 13776 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_134
timestamp 1698431365
transform 1 0 16352 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698431365
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_146
timestamp 1698431365
transform 1 0 17696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_160
timestamp 1698431365
transform 1 0 19264 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_198
timestamp 1698431365
transform 1 0 23520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_202
timestamp 1698431365
transform 1 0 23968 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_216
timestamp 1698431365
transform 1 0 25536 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_267
timestamp 1698431365
transform 1 0 31248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_271
timestamp 1698431365
transform 1 0 31696 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_292
timestamp 1698431365
transform 1 0 34048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_320
timestamp 1698431365
transform 1 0 37184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_348
timestamp 1698431365
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_362
timestamp 1698431365
transform 1 0 41888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_409
timestamp 1698431365
transform 1 0 47152 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_470
timestamp 1698431365
transform 1 0 53984 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_477
timestamp 1698431365
transform 1 0 54768 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_481
timestamp 1698431365
transform 1 0 55216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_489
timestamp 1698431365
transform 1 0 56112 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_494
timestamp 1698431365
transform 1 0 56672 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_508
timestamp 1698431365
transform 1 0 58240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_6
timestamp 1698431365
transform 1 0 2016 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_21
timestamp 1698431365
transform 1 0 3696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_23
timestamp 1698431365
transform 1 0 3920 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_30
timestamp 1698431365
transform 1 0 4704 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_39
timestamp 1698431365
transform 1 0 5712 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_63
timestamp 1698431365
transform 1 0 8400 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_73
timestamp 1698431365
transform 1 0 9520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_77
timestamp 1698431365
transform 1 0 9968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_95
timestamp 1698431365
transform 1 0 11984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_97
timestamp 1698431365
transform 1 0 12208 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_135
timestamp 1698431365
transform 1 0 16464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_139
timestamp 1698431365
transform 1 0 16912 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_155
timestamp 1698431365
transform 1 0 18704 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_159
timestamp 1698431365
transform 1 0 19152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_162
timestamp 1698431365
transform 1 0 19488 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_166
timestamp 1698431365
transform 1 0 19936 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_168
timestamp 1698431365
transform 1 0 20160 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_196
timestamp 1698431365
transform 1 0 23296 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_200
timestamp 1698431365
transform 1 0 23744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_296
timestamp 1698431365
transform 1 0 34496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_300
timestamp 1698431365
transform 1 0 34944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_304
timestamp 1698431365
transform 1 0 35392 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_313
timestamp 1698431365
transform 1 0 36400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_332
timestamp 1698431365
transform 1 0 38528 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_336
timestamp 1698431365
transform 1 0 38976 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_342
timestamp 1698431365
transform 1 0 39648 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_346
timestamp 1698431365
transform 1 0 40096 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_376
timestamp 1698431365
transform 1 0 43456 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_380
timestamp 1698431365
transform 1 0 43904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_382
timestamp 1698431365
transform 1 0 44128 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_404
timestamp 1698431365
transform 1 0 46592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_406
timestamp 1698431365
transform 1 0 46816 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_430
timestamp 1698431365
transform 1 0 49504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_453
timestamp 1698431365
transform 1 0 52080 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_461
timestamp 1698431365
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_465
timestamp 1698431365
transform 1 0 53424 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_482
timestamp 1698431365
transform 1 0 55328 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_504
timestamp 1698431365
transform 1 0 57792 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_508
timestamp 1698431365
transform 1 0 58240 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_31
timestamp 1698431365
transform 1 0 4816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_103
timestamp 1698431365
transform 1 0 12880 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_109
timestamp 1698431365
transform 1 0 13552 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_118
timestamp 1698431365
transform 1 0 14560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_120
timestamp 1698431365
transform 1 0 14784 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_131
timestamp 1698431365
transform 1 0 16016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_135
timestamp 1698431365
transform 1 0 16464 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_177
timestamp 1698431365
transform 1 0 21168 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_181
timestamp 1698431365
transform 1 0 21616 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_183
timestamp 1698431365
transform 1 0 21840 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_186
timestamp 1698431365
transform 1 0 22176 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_194
timestamp 1698431365
transform 1 0 23072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_196
timestamp 1698431365
transform 1 0 23296 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_214
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_242
timestamp 1698431365
transform 1 0 28448 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_244
timestamp 1698431365
transform 1 0 28672 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_253
timestamp 1698431365
transform 1 0 29680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_255
timestamp 1698431365
transform 1 0 29904 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_273
timestamp 1698431365
transform 1 0 31920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_289
timestamp 1698431365
transform 1 0 33712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_318
timestamp 1698431365
transform 1 0 36960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698431365
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_328
timestamp 1698431365
transform 1 0 38080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_344
timestamp 1698431365
transform 1 0 39872 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_348
timestamp 1698431365
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_362
timestamp 1698431365
transform 1 0 41888 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_396
timestamp 1698431365
transform 1 0 45696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_400
timestamp 1698431365
transform 1 0 46144 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_404
timestamp 1698431365
transform 1 0 46592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_406
timestamp 1698431365
transform 1 0 46816 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_434
timestamp 1698431365
transform 1 0 49952 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_438
timestamp 1698431365
transform 1 0 50400 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_458
timestamp 1698431365
transform 1 0 52640 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_466
timestamp 1698431365
transform 1 0 53536 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_470
timestamp 1698431365
transform 1 0 53984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_485
timestamp 1698431365
transform 1 0 55664 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_489
timestamp 1698431365
transform 1 0 56112 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_504
timestamp 1698431365
transform 1 0 57792 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_4
timestamp 1698431365
transform 1 0 1792 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_20
timestamp 1698431365
transform 1 0 3584 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_63
timestamp 1698431365
transform 1 0 8400 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_71
timestamp 1698431365
transform 1 0 9296 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_74
timestamp 1698431365
transform 1 0 9632 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_78
timestamp 1698431365
transform 1 0 10080 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_92
timestamp 1698431365
transform 1 0 11648 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_98
timestamp 1698431365
transform 1 0 12320 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_102
timestamp 1698431365
transform 1 0 12768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_136
timestamp 1698431365
transform 1 0 16576 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_140
timestamp 1698431365
transform 1 0 17024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_166
timestamp 1698431365
transform 1 0 19936 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_200
timestamp 1698431365
transform 1 0 23744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_204
timestamp 1698431365
transform 1 0 24192 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_210
timestamp 1698431365
transform 1 0 24864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_216
timestamp 1698431365
transform 1 0 25536 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_265
timestamp 1698431365
transform 1 0 31024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_267
timestamp 1698431365
transform 1 0 31248 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_294
timestamp 1698431365
transform 1 0 34272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_298
timestamp 1698431365
transform 1 0 34720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_300
timestamp 1698431365
transform 1 0 34944 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_313
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_365
timestamp 1698431365
transform 1 0 42224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_373
timestamp 1698431365
transform 1 0 43120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_375
timestamp 1698431365
transform 1 0 43344 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_378
timestamp 1698431365
transform 1 0 43680 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_382
timestamp 1698431365
transform 1 0 44128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_400
timestamp 1698431365
transform 1 0 46144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_402
timestamp 1698431365
transform 1 0 46368 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_411
timestamp 1698431365
transform 1 0 47376 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_436
timestamp 1698431365
transform 1 0 50176 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_462
timestamp 1698431365
transform 1 0 53088 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_466
timestamp 1698431365
transform 1 0 53536 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_474
timestamp 1698431365
transform 1 0 54432 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_478
timestamp 1698431365
transform 1 0 54880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_12
timestamp 1698431365
transform 1 0 2688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_32
timestamp 1698431365
transform 1 0 4928 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_36
timestamp 1698431365
transform 1 0 5376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_67
timestamp 1698431365
transform 1 0 8848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_76
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_78
timestamp 1698431365
transform 1 0 10080 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_110
timestamp 1698431365
transform 1 0 13664 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_118
timestamp 1698431365
transform 1 0 14560 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_132
timestamp 1698431365
transform 1 0 16128 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_167
timestamp 1698431365
transform 1 0 20048 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_171
timestamp 1698431365
transform 1 0 20496 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_173
timestamp 1698431365
transform 1 0 20720 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_197
timestamp 1698431365
transform 1 0 23408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_224
timestamp 1698431365
transform 1 0 26432 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_228
timestamp 1698431365
transform 1 0 26880 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_244
timestamp 1698431365
transform 1 0 28672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_246
timestamp 1698431365
transform 1 0 28896 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_267
timestamp 1698431365
transform 1 0 31248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_320
timestamp 1698431365
transform 1 0 37184 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_324
timestamp 1698431365
transform 1 0 37632 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_373
timestamp 1698431365
transform 1 0 43120 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_377
timestamp 1698431365
transform 1 0 43568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_404
timestamp 1698431365
transform 1 0 46592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_408
timestamp 1698431365
transform 1 0 47040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_442
timestamp 1698431365
transform 1 0 50848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_459
timestamp 1698431365
transform 1 0 52752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_505
timestamp 1698431365
transform 1 0 57904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_33
timestamp 1698431365
transform 1 0 5040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_49
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_51
timestamp 1698431365
transform 1 0 7056 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_67
timestamp 1698431365
transform 1 0 8848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_75
timestamp 1698431365
transform 1 0 9744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_97
timestamp 1698431365
transform 1 0 12208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_109
timestamp 1698431365
transform 1 0 13552 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_118
timestamp 1698431365
transform 1 0 14560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_120
timestamp 1698431365
transform 1 0 14784 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_139
timestamp 1698431365
transform 1 0 16912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_143
timestamp 1698431365
transform 1 0 17360 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_151
timestamp 1698431365
transform 1 0 18256 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_153
timestamp 1698431365
transform 1 0 18480 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_166
timestamp 1698431365
transform 1 0 19936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_170
timestamp 1698431365
transform 1 0 20384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_240
timestamp 1698431365
transform 1 0 28224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_242
timestamp 1698431365
transform 1 0 28448 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_310
timestamp 1698431365
transform 1 0 36064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_375
timestamp 1698431365
transform 1 0 43344 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_379
timestamp 1698431365
transform 1 0 43792 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_412
timestamp 1698431365
transform 1 0 47488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_416
timestamp 1698431365
transform 1 0 47936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_432
timestamp 1698431365
transform 1 0 49728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_451
timestamp 1698431365
transform 1 0 51856 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_475
timestamp 1698431365
transform 1 0 54544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_477
timestamp 1698431365
transform 1 0 54768 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_8
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_12
timestamp 1698431365
transform 1 0 2688 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_21
timestamp 1698431365
transform 1 0 3696 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_32
timestamp 1698431365
transform 1 0 4928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_40
timestamp 1698431365
transform 1 0 5824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_74
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_111
timestamp 1698431365
transform 1 0 13776 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_113
timestamp 1698431365
transform 1 0 14000 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_166
timestamp 1698431365
transform 1 0 19936 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_168
timestamp 1698431365
transform 1 0 20160 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_174
timestamp 1698431365
transform 1 0 20832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_176
timestamp 1698431365
transform 1 0 21056 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_185
timestamp 1698431365
transform 1 0 22064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_218
timestamp 1698431365
transform 1 0 25760 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_226
timestamp 1698431365
transform 1 0 26656 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_230
timestamp 1698431365
transform 1 0 27104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_232
timestamp 1698431365
transform 1 0 27328 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_297
timestamp 1698431365
transform 1 0 34608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_301
timestamp 1698431365
transform 1 0 35056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_305
timestamp 1698431365
transform 1 0 35504 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_321
timestamp 1698431365
transform 1 0 37296 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_325
timestamp 1698431365
transform 1 0 37744 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_333
timestamp 1698431365
transform 1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_335
timestamp 1698431365
transform 1 0 38864 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_357
timestamp 1698431365
transform 1 0 41328 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_373
timestamp 1698431365
transform 1 0 43120 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_381
timestamp 1698431365
transform 1 0 44016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_388
timestamp 1698431365
transform 1 0 44800 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_414
timestamp 1698431365
transform 1 0 47712 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_418
timestamp 1698431365
transform 1 0 48160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_451
timestamp 1698431365
transform 1 0 51856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_473
timestamp 1698431365
transform 1 0 54320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_475
timestamp 1698431365
transform 1 0 54544 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_482
timestamp 1698431365
transform 1 0 55328 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_504
timestamp 1698431365
transform 1 0 57792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_508
timestamp 1698431365
transform 1 0 58240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_31
timestamp 1698431365
transform 1 0 4816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_66
timestamp 1698431365
transform 1 0 8736 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_74
timestamp 1698431365
transform 1 0 9632 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_76
timestamp 1698431365
transform 1 0 9856 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_98
timestamp 1698431365
transform 1 0 12320 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_102
timestamp 1698431365
transform 1 0 12768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_123
timestamp 1698431365
transform 1 0 15120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_138
timestamp 1698431365
transform 1 0 16800 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_144
timestamp 1698431365
transform 1 0 17472 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_169
timestamp 1698431365
transform 1 0 20272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_181
timestamp 1698431365
transform 1 0 21616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_207
timestamp 1698431365
transform 1 0 24528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_211
timestamp 1698431365
transform 1 0 24976 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_251
timestamp 1698431365
transform 1 0 29456 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_257
timestamp 1698431365
transform 1 0 30128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_278
timestamp 1698431365
transform 1 0 32480 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_282
timestamp 1698431365
transform 1 0 32928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_286
timestamp 1698431365
transform 1 0 33376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_288
timestamp 1698431365
transform 1 0 33600 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_302
timestamp 1698431365
transform 1 0 35168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_304
timestamp 1698431365
transform 1 0 35392 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_329
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_333
timestamp 1698431365
transform 1 0 38640 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_336
timestamp 1698431365
transform 1 0 38976 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_348
timestamp 1698431365
transform 1 0 40320 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_356
timestamp 1698431365
transform 1 0 41216 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_360
timestamp 1698431365
transform 1 0 41664 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_381
timestamp 1698431365
transform 1 0 44016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_395
timestamp 1698431365
transform 1 0 45584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_397
timestamp 1698431365
transform 1 0 45808 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_422
timestamp 1698431365
transform 1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_429
timestamp 1698431365
transform 1 0 49392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_431
timestamp 1698431365
transform 1 0 49616 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_434
timestamp 1698431365
transform 1 0 49952 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_462
timestamp 1698431365
transform 1 0 53088 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_468
timestamp 1698431365
transform 1 0 53760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_472
timestamp 1698431365
transform 1 0 54208 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_20
timestamp 1698431365
transform 1 0 3584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_28
timestamp 1698431365
transform 1 0 4480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_32
timestamp 1698431365
transform 1 0 4928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_36
timestamp 1698431365
transform 1 0 5376 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_44
timestamp 1698431365
transform 1 0 6272 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_48
timestamp 1698431365
transform 1 0 6720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_56
timestamp 1698431365
transform 1 0 7616 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_78
timestamp 1698431365
transform 1 0 10080 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_87
timestamp 1698431365
transform 1 0 11088 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_146
timestamp 1698431365
transform 1 0 17696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_148
timestamp 1698431365
transform 1 0 17920 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_176
timestamp 1698431365
transform 1 0 21056 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_180
timestamp 1698431365
transform 1 0 21504 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_184
timestamp 1698431365
transform 1 0 21952 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_190
timestamp 1698431365
transform 1 0 22624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_194
timestamp 1698431365
transform 1 0 23072 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_224
timestamp 1698431365
transform 1 0 26432 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_228
timestamp 1698431365
transform 1 0 26880 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_247
timestamp 1698431365
transform 1 0 29008 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_255
timestamp 1698431365
transform 1 0 29904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_286
timestamp 1698431365
transform 1 0 33376 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_307
timestamp 1698431365
transform 1 0 35728 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_311
timestamp 1698431365
transform 1 0 36176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_313
timestamp 1698431365
transform 1 0 36400 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_347
timestamp 1698431365
transform 1 0 40208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_358
timestamp 1698431365
transform 1 0 41440 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_362
timestamp 1698431365
transform 1 0 41888 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_385
timestamp 1698431365
transform 1 0 44464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_387
timestamp 1698431365
transform 1 0 44688 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_463
timestamp 1698431365
transform 1 0 53200 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_467
timestamp 1698431365
transform 1 0 53648 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698431365
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_12
timestamp 1698431365
transform 1 0 2688 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_31
timestamp 1698431365
transform 1 0 4816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_45
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_47
timestamp 1698431365
transform 1 0 6608 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_68
timestamp 1698431365
transform 1 0 8960 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_132
timestamp 1698431365
transform 1 0 16128 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_148
timestamp 1698431365
transform 1 0 17920 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_152
timestamp 1698431365
transform 1 0 18368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_166
timestamp 1698431365
transform 1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_170
timestamp 1698431365
transform 1 0 20384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_199
timestamp 1698431365
transform 1 0 23632 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_221
timestamp 1698431365
transform 1 0 26096 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_240
timestamp 1698431365
transform 1 0 28224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_271
timestamp 1698431365
transform 1 0 31696 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_279
timestamp 1698431365
transform 1 0 32592 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_292
timestamp 1698431365
transform 1 0 34048 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_294
timestamp 1698431365
transform 1 0 34272 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_297
timestamp 1698431365
transform 1 0 34608 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_305
timestamp 1698431365
transform 1 0 35504 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_322
timestamp 1698431365
transform 1 0 37408 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_326
timestamp 1698431365
transform 1 0 37856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_330
timestamp 1698431365
transform 1 0 38304 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_373
timestamp 1698431365
transform 1 0 43120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_397
timestamp 1698431365
transform 1 0 45808 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_399
timestamp 1698431365
transform 1 0 46032 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_439
timestamp 1698431365
transform 1 0 50512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_32
timestamp 1698431365
transform 1 0 4928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_63
timestamp 1698431365
transform 1 0 8400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_67
timestamp 1698431365
transform 1 0 8848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_69
timestamp 1698431365
transform 1 0 9072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_76
timestamp 1698431365
transform 1 0 9856 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_106
timestamp 1698431365
transform 1 0 13216 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_113
timestamp 1698431365
transform 1 0 14000 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_127
timestamp 1698431365
transform 1 0 15568 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_135
timestamp 1698431365
transform 1 0 16464 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_181
timestamp 1698431365
transform 1 0 21616 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_185
timestamp 1698431365
transform 1 0 22064 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_193
timestamp 1698431365
transform 1 0 22960 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_197
timestamp 1698431365
transform 1 0 23408 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_228
timestamp 1698431365
transform 1 0 26880 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_230
timestamp 1698431365
transform 1 0 27104 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_299
timestamp 1698431365
transform 1 0 34832 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_301
timestamp 1698431365
transform 1 0 35056 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_332
timestamp 1698431365
transform 1 0 38528 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_336
timestamp 1698431365
transform 1 0 38976 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_368
timestamp 1698431365
transform 1 0 42560 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_398
timestamp 1698431365
transform 1 0 45920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_402
timestamp 1698431365
transform 1 0 46368 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_410
timestamp 1698431365
transform 1 0 47264 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_439
timestamp 1698431365
transform 1 0 50512 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_505
timestamp 1698431365
transform 1 0 57904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_16
timestamp 1698431365
transform 1 0 3136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_18
timestamp 1698431365
transform 1 0 3360 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_24
timestamp 1698431365
transform 1 0 4032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_42
timestamp 1698431365
transform 1 0 6048 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_44
timestamp 1698431365
transform 1 0 6272 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_50
timestamp 1698431365
transform 1 0 6944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_62
timestamp 1698431365
transform 1 0 8288 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_66
timestamp 1698431365
transform 1 0 8736 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_74
timestamp 1698431365
transform 1 0 9632 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_92
timestamp 1698431365
transform 1 0 11648 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_100
timestamp 1698431365
transform 1 0 12544 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_111
timestamp 1698431365
transform 1 0 13776 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_138
timestamp 1698431365
transform 1 0 16800 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_142
timestamp 1698431365
transform 1 0 17248 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_170
timestamp 1698431365
transform 1 0 20384 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_228
timestamp 1698431365
transform 1 0 26880 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_232
timestamp 1698431365
transform 1 0 27328 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_253
timestamp 1698431365
transform 1 0 29680 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_257
timestamp 1698431365
transform 1 0 30128 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_265
timestamp 1698431365
transform 1 0 31024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_273
timestamp 1698431365
transform 1 0 31920 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_275
timestamp 1698431365
transform 1 0 32144 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_278
timestamp 1698431365
transform 1 0 32480 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_294
timestamp 1698431365
transform 1 0 34272 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_310
timestamp 1698431365
transform 1 0 36064 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_325
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_329
timestamp 1698431365
transform 1 0 38192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_353
timestamp 1698431365
transform 1 0 40880 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_389
timestamp 1698431365
transform 1 0 44912 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_392
timestamp 1698431365
transform 1 0 45248 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698431365
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_476
timestamp 1698431365
transform 1 0 54656 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_507
timestamp 1698431365
transform 1 0 58128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_10
timestamp 1698431365
transform 1 0 2464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_105
timestamp 1698431365
transform 1 0 13104 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_113
timestamp 1698431365
transform 1 0 14000 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_117
timestamp 1698431365
transform 1 0 14448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_132
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_144
timestamp 1698431365
transform 1 0 17472 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_147
timestamp 1698431365
transform 1 0 17808 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_167
timestamp 1698431365
transform 1 0 20048 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_172
timestamp 1698431365
transform 1 0 20608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_176
timestamp 1698431365
transform 1 0 21056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_180
timestamp 1698431365
transform 1 0 21504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_182
timestamp 1698431365
transform 1 0 21728 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_216
timestamp 1698431365
transform 1 0 25536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_218
timestamp 1698431365
transform 1 0 25760 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_231
timestamp 1698431365
transform 1 0 27216 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_235
timestamp 1698431365
transform 1 0 27664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_237
timestamp 1698431365
transform 1 0 27888 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_259
timestamp 1698431365
transform 1 0 30352 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_263
timestamp 1698431365
transform 1 0 30800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_265
timestamp 1698431365
transform 1 0 31024 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_278
timestamp 1698431365
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_288
timestamp 1698431365
transform 1 0 33600 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_305
timestamp 1698431365
transform 1 0 35504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_307
timestamp 1698431365
transform 1 0 35728 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_336
timestamp 1698431365
transform 1 0 38976 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_360
timestamp 1698431365
transform 1 0 41664 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_364
timestamp 1698431365
transform 1 0 42112 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_389
timestamp 1698431365
transform 1 0 44912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_486
timestamp 1698431365
transform 1 0 55776 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_504
timestamp 1698431365
transform 1 0 57792 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_508
timestamp 1698431365
transform 1 0 58240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_10
timestamp 1698431365
transform 1 0 2464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_19
timestamp 1698431365
transform 1 0 3472 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_42
timestamp 1698431365
transform 1 0 6048 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_58
timestamp 1698431365
transform 1 0 7840 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_65
timestamp 1698431365
transform 1 0 8624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_74
timestamp 1698431365
transform 1 0 9632 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_78
timestamp 1698431365
transform 1 0 10080 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_87
timestamp 1698431365
transform 1 0 11088 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_103
timestamp 1698431365
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_111
timestamp 1698431365
transform 1 0 13776 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_113
timestamp 1698431365
transform 1 0 14000 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_137
timestamp 1698431365
transform 1 0 16688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_139
timestamp 1698431365
transform 1 0 16912 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_145
timestamp 1698431365
transform 1 0 17584 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_147
timestamp 1698431365
transform 1 0 17808 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_173
timestamp 1698431365
transform 1 0 20720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_200
timestamp 1698431365
transform 1 0 23744 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_209
timestamp 1698431365
transform 1 0 24752 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_213
timestamp 1698431365
transform 1 0 25200 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_237
timestamp 1698431365
transform 1 0 27888 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_282
timestamp 1698431365
transform 1 0 32928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_301
timestamp 1698431365
transform 1 0 35056 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_330
timestamp 1698431365
transform 1 0 38304 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_352
timestamp 1698431365
transform 1 0 40768 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_358
timestamp 1698431365
transform 1 0 41440 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_373
timestamp 1698431365
transform 1 0 43120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_375
timestamp 1698431365
transform 1 0 43344 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698431365
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_440
timestamp 1698431365
transform 1 0 50624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_444
timestamp 1698431365
transform 1 0 51072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_448
timestamp 1698431365
transform 1 0 51520 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_506
timestamp 1698431365
transform 1 0 58016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_508
timestamp 1698431365
transform 1 0 58240 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_50
timestamp 1698431365
transform 1 0 6944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_54
timestamp 1698431365
transform 1 0 7392 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_80
timestamp 1698431365
transform 1 0 10304 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_96
timestamp 1698431365
transform 1 0 12096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_165
timestamp 1698431365
transform 1 0 19824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_169
timestamp 1698431365
transform 1 0 20272 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_175
timestamp 1698431365
transform 1 0 20944 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_199
timestamp 1698431365
transform 1 0 23632 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_203
timestamp 1698431365
transform 1 0 24080 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_207
timestamp 1698431365
transform 1 0 24528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698431365
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_225
timestamp 1698431365
transform 1 0 26544 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_233
timestamp 1698431365
transform 1 0 27440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_255
timestamp 1698431365
transform 1 0 29904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_278
timestamp 1698431365
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_288
timestamp 1698431365
transform 1 0 33600 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_292
timestamp 1698431365
transform 1 0 34048 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_298
timestamp 1698431365
transform 1 0 34720 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_306
timestamp 1698431365
transform 1 0 35616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_310
timestamp 1698431365
transform 1 0 36064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_342
timestamp 1698431365
transform 1 0 39648 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_365
timestamp 1698431365
transform 1 0 42224 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_371
timestamp 1698431365
transform 1 0 42896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_407
timestamp 1698431365
transform 1 0 46928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_411
timestamp 1698431365
transform 1 0 47376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_413
timestamp 1698431365
transform 1 0 47600 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_480
timestamp 1698431365
transform 1 0 55104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_484
timestamp 1698431365
transform 1 0 55552 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_505
timestamp 1698431365
transform 1 0 57904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_31
timestamp 1698431365
transform 1 0 4816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_41
timestamp 1698431365
transform 1 0 5936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_49
timestamp 1698431365
transform 1 0 6832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_53
timestamp 1698431365
transform 1 0 7280 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_57
timestamp 1698431365
transform 1 0 7728 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_59
timestamp 1698431365
transform 1 0 7952 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_89
timestamp 1698431365
transform 1 0 11312 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_93
timestamp 1698431365
transform 1 0 11760 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_97
timestamp 1698431365
transform 1 0 12208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_114
timestamp 1698431365
transform 1 0 14112 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_182
timestamp 1698431365
transform 1 0 21728 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_186
timestamp 1698431365
transform 1 0 22176 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_215
timestamp 1698431365
transform 1 0 25424 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_219
timestamp 1698431365
transform 1 0 25872 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_223
timestamp 1698431365
transform 1 0 26320 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_262
timestamp 1698431365
transform 1 0 30688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_266
timestamp 1698431365
transform 1 0 31136 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_301
timestamp 1698431365
transform 1 0 35056 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_307
timestamp 1698431365
transform 1 0 35728 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_448
timestamp 1698431365
transform 1 0 51520 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_452
timestamp 1698431365
transform 1 0 51968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_454
timestamp 1698431365
transform 1 0 52192 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_459
timestamp 1698431365
transform 1 0 52752 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_477
timestamp 1698431365
transform 1 0 54768 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_481
timestamp 1698431365
transform 1 0 55216 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_10
timestamp 1698431365
transform 1 0 2464 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_32
timestamp 1698431365
transform 1 0 4928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_34
timestamp 1698431365
transform 1 0 5152 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_45
timestamp 1698431365
transform 1 0 6384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_55
timestamp 1698431365
transform 1 0 7504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_63
timestamp 1698431365
transform 1 0 8400 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_65
timestamp 1698431365
transform 1 0 8624 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_68
timestamp 1698431365
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_74
timestamp 1698431365
transform 1 0 9632 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_81
timestamp 1698431365
transform 1 0 10416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_85
timestamp 1698431365
transform 1 0 10864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_89
timestamp 1698431365
transform 1 0 11312 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_93
timestamp 1698431365
transform 1 0 11760 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_96
timestamp 1698431365
transform 1 0 12096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_129
timestamp 1698431365
transform 1 0 15792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_131
timestamp 1698431365
transform 1 0 16016 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_138
timestamp 1698431365
transform 1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_148
timestamp 1698431365
transform 1 0 17920 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_152
timestamp 1698431365
transform 1 0 18368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_176
timestamp 1698431365
transform 1 0 21056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_178
timestamp 1698431365
transform 1 0 21280 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_199
timestamp 1698431365
transform 1 0 23632 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_209
timestamp 1698431365
transform 1 0 24752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_225
timestamp 1698431365
transform 1 0 26544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_229
timestamp 1698431365
transform 1 0 26992 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_242
timestamp 1698431365
transform 1 0 28448 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_246
timestamp 1698431365
transform 1 0 28896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_248
timestamp 1698431365
transform 1 0 29120 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_257
timestamp 1698431365
transform 1 0 30128 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_261
timestamp 1698431365
transform 1 0 30576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_265
timestamp 1698431365
transform 1 0 31024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_267
timestamp 1698431365
transform 1 0 31248 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_319
timestamp 1698431365
transform 1 0 37072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_348
timestamp 1698431365
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_364
timestamp 1698431365
transform 1 0 42112 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_366
timestamp 1698431365
transform 1 0 42336 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_416
timestamp 1698431365
transform 1 0 47936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_432
timestamp 1698431365
transform 1 0 49728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_478
timestamp 1698431365
transform 1 0 54880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_482
timestamp 1698431365
transform 1 0 55328 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_504
timestamp 1698431365
transform 1 0 57792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_506
timestamp 1698431365
transform 1 0 58016 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_26
timestamp 1698431365
transform 1 0 4256 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_30
timestamp 1698431365
transform 1 0 4704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_109
timestamp 1698431365
transform 1 0 13552 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_116
timestamp 1698431365
transform 1 0 14336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_120
timestamp 1698431365
transform 1 0 14784 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_152
timestamp 1698431365
transform 1 0 18368 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_160
timestamp 1698431365
transform 1 0 19264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_174
timestamp 1698431365
transform 1 0 20832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_194
timestamp 1698431365
transform 1 0 23072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_227
timestamp 1698431365
transform 1 0 26768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_229
timestamp 1698431365
transform 1 0 26992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_236
timestamp 1698431365
transform 1 0 27776 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_255
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_269
timestamp 1698431365
transform 1 0 31472 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_273
timestamp 1698431365
transform 1 0 31920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_277
timestamp 1698431365
transform 1 0 32368 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_287
timestamp 1698431365
transform 1 0 33488 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_296
timestamp 1698431365
transform 1 0 34496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_310
timestamp 1698431365
transform 1 0 36064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_328
timestamp 1698431365
transform 1 0 38080 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_452
timestamp 1698431365
transform 1 0 51968 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_454
timestamp 1698431365
transform 1 0 52192 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_465
timestamp 1698431365
transform 1 0 53424 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_467
timestamp 1698431365
transform 1 0 53648 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_504
timestamp 1698431365
transform 1 0 57792 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_508
timestamp 1698431365
transform 1 0 58240 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_53
timestamp 1698431365
transform 1 0 7280 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_65
timestamp 1698431365
transform 1 0 8624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_74
timestamp 1698431365
transform 1 0 9632 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_85
timestamp 1698431365
transform 1 0 10864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_138
timestamp 1698431365
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_146
timestamp 1698431365
transform 1 0 17696 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_194
timestamp 1698431365
transform 1 0 23072 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_196
timestamp 1698431365
transform 1 0 23296 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_216
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_248
timestamp 1698431365
transform 1 0 29120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_250
timestamp 1698431365
transform 1 0 29344 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_292
timestamp 1698431365
transform 1 0 34048 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_298
timestamp 1698431365
transform 1 0 34720 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_302
timestamp 1698431365
transform 1 0 35168 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_358
timestamp 1698431365
transform 1 0 41440 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_362
timestamp 1698431365
transform 1 0 41888 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_366
timestamp 1698431365
transform 1 0 42336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_418
timestamp 1698431365
transform 1 0 48160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_445
timestamp 1698431365
transform 1 0 51184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_473
timestamp 1698431365
transform 1 0 54320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_482
timestamp 1698431365
transform 1 0 55328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_486
timestamp 1698431365
transform 1 0 55776 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_497
timestamp 1698431365
transform 1 0 57008 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_505
timestamp 1698431365
transform 1 0 57904 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_31
timestamp 1698431365
transform 1 0 4816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_33
timestamp 1698431365
transform 1 0 5040 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_36
timestamp 1698431365
transform 1 0 5376 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_38
timestamp 1698431365
transform 1 0 5600 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_70
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_72
timestamp 1698431365
transform 1 0 9408 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_108
timestamp 1698431365
transform 1 0 13440 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_112
timestamp 1698431365
transform 1 0 13888 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_114
timestamp 1698431365
transform 1 0 14112 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_125
timestamp 1698431365
transform 1 0 15344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_127
timestamp 1698431365
transform 1 0 15568 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_130
timestamp 1698431365
transform 1 0 15904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_134
timestamp 1698431365
transform 1 0 16352 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_148
timestamp 1698431365
transform 1 0 17920 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_152
timestamp 1698431365
transform 1 0 18368 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_165
timestamp 1698431365
transform 1 0 19824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_167
timestamp 1698431365
transform 1 0 20048 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_185
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_187
timestamp 1698431365
transform 1 0 22288 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_200
timestamp 1698431365
transform 1 0 23744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_206
timestamp 1698431365
transform 1 0 24416 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_224
timestamp 1698431365
transform 1 0 26432 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_269
timestamp 1698431365
transform 1 0 31472 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_271
timestamp 1698431365
transform 1 0 31696 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_274
timestamp 1698431365
transform 1 0 32032 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_276
timestamp 1698431365
transform 1 0 32256 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_360
timestamp 1698431365
transform 1 0 41664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_370
timestamp 1698431365
transform 1 0 42784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_376
timestamp 1698431365
transform 1 0 43456 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_378
timestamp 1698431365
transform 1 0 43680 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_416
timestamp 1698431365
transform 1 0 47936 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_432
timestamp 1698431365
transform 1 0 49728 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_434
timestamp 1698431365
transform 1 0 49952 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_441
timestamp 1698431365
transform 1 0 50736 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_444
timestamp 1698431365
transform 1 0 51072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_446
timestamp 1698431365
transform 1 0 51296 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_471
timestamp 1698431365
transform 1 0 54096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_475
timestamp 1698431365
transform 1 0 54544 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_486
timestamp 1698431365
transform 1 0 55776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_490
timestamp 1698431365
transform 1 0 56224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_494
timestamp 1698431365
transform 1 0 56672 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_498
timestamp 1698431365
transform 1 0 57120 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_506
timestamp 1698431365
transform 1 0 58016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_508
timestamp 1698431365
transform 1 0 58240 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 3472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 8400 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698431365
transform 1 0 47264 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input4
timestamp 1698431365
transform 1 0 52080 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 14560 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input6
timestamp 1698431365
transform 1 0 3360 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 2912 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 2240 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 1904 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input16
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input17
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input18
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input19
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input20
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input21
timestamp 1698431365
transform 1 0 2240 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 30800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input25
timestamp 1698431365
transform -1 0 33040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 37856 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 10416 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input29
timestamp 1698431365
transform -1 0 55776 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 54096 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 50736 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input32
timestamp 1698431365
transform -1 0 49056 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 48160 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 47264 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 42112 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform -1 0 41440 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output37 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 56784 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output38
timestamp 1698431365
transform 1 0 18704 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output39
timestamp 1698431365
transform 1 0 16800 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output40
timestamp 1698431365
transform 1 0 14224 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output41 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output42
timestamp 1698431365
transform 1 0 9744 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output43
timestamp 1698431365
transform 1 0 7504 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output44
timestamp 1698431365
transform 1 0 5264 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output45
timestamp 1698431365
transform -1 0 4032 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output46
timestamp 1698431365
transform -1 0 37408 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output47
timestamp 1698431365
transform -1 0 36064 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output48
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output49
timestamp 1698431365
transform -1 0 31472 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output50
timestamp 1698431365
transform -1 0 28000 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output51
timestamp 1698431365
transform 1 0 24864 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output52
timestamp 1698431365
transform 1 0 22624 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output53
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_43 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_44
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_45
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer1
timestamp 1698431365
transform -1 0 52304 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer2
timestamp 1698431365
transform -1 0 22960 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer3
timestamp 1698431365
transform 1 0 28112 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer4
timestamp 1698431365
transform 1 0 31472 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer5
timestamp 1698431365
transform -1 0 24864 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer6
timestamp 1698431365
transform -1 0 48384 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer7
timestamp 1698431365
transform -1 0 55776 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer8
timestamp 1698431365
transform 1 0 19152 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer9
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer10
timestamp 1698431365
transform 1 0 38528 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer11
timestamp 1698431365
transform -1 0 42224 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer12
timestamp 1698431365
transform -1 0 40880 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  rebuffer13
timestamp 1698431365
transform -1 0 28000 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  rebuffer14
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer15
timestamp 1698431365
transform -1 0 42896 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer16
timestamp 1698431365
transform 1 0 42224 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer17
timestamp 1698431365
transform -1 0 42672 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer18 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33600 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer19
timestamp 1698431365
transform -1 0 25536 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer20
timestamp 1698431365
transform -1 0 40208 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer21
timestamp 1698431365
transform -1 0 42000 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer22
timestamp 1698431365
transform 1 0 39536 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer23
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer24
timestamp 1698431365
transform 1 0 40096 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer25
timestamp 1698431365
transform -1 0 42896 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_86 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_87
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_88
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_89
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_104
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_105
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_106
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_109
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_110
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_111
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_112
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_113
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_114
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_115
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_116
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_117
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_118
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_119
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_120
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_121
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_122
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_123
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_124
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_125
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_126
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_127
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_128
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_129
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_130
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_131
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_132
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_133
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_134
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_135
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_136
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_137
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_138
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_139
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_140
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_141
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_142
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_143
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_144
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_145
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_146
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_147
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_148
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_149
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_150
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_151
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_152
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_153
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_154
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_155
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_156
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_157
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_158
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_159
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_160
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_161
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_162
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_163
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_164
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_165
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_166
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_167
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_168
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_169
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_170
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_171
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_172
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_173
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_174
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_175
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_176
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_177
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_178
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_179
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_180
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_181
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_183
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_184
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_185
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_186
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_187
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_188
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_189
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_190
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_191
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_192
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_193
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_194
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_195
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_196
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_197
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_198
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_199
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_200
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_201
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_202
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_203
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_204
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_205
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_206
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_207
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_208
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_209
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_210
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_211
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_212
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_213
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_214
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_215
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_216
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_217
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_218
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_219
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_220
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_221
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_222
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_223
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_224
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_225
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_226
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_227
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_228
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_229
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_230
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_231
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_232
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_233
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_234
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_235
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_236
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_237
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_238
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_239
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_240
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_241
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_242
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_243
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_244
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_245
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_246
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_247
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_248
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_249
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_250
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_251
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_252
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_253
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_254
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_255
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_256
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_257
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_258
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_259
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_260
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_261
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_262
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_263
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_264
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_265
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_266
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_267
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_268
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_269
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_270
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_271
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_272
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_273
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_274
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_275
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_276
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_277
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_278
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_279
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_280
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_281
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_282
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_283
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_284
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_285
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_286
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_287
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_288
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_289
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_290
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_291
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_292
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_293
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_294
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_295
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_296
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_297
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_298
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_299
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_300
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_301
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_302
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_303
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_304
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_305
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_306
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_307
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_308
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_309
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_310
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_311
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_312
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_313
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_314
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_315
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_316
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_317
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_318
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_319
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_320
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_321
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_322
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_323
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_324
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_325
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_326
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_327
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_328
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_329
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_330
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_331
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_332
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_333
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_334
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_335
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_336
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_337
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_338
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_339
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_340
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_341
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_342
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_343
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_344
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_345
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_346
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_347
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_348
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_349
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_350
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_351
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_352
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_353
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_354
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_355
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_356
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_357
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_358
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_359
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_360
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_361
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_362
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_363
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_364
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_365
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_366
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_367
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_368
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_369
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_370
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_371
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_372
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_373
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_374
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_375
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_376
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_377
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_378
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_379
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_380
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_381
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_382
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_383
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_384
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_385
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_386
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_387
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_388
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_389
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_390
timestamp 1698431365
transform 1 0 16576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_391
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_392
timestamp 1698431365
transform 1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_393
timestamp 1698431365
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_394
timestamp 1698431365
transform 1 0 31808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_395
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_396
timestamp 1698431365
transform 1 0 39424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_397
timestamp 1698431365
transform 1 0 43232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_398
timestamp 1698431365
transform 1 0 47040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_399
timestamp 1698431365
transform 1 0 50848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_400
timestamp 1698431365
transform 1 0 54656 0 1 36064
box -86 -86 310 870
<< labels >>
flabel metal2 s 56672 39200 56784 40000 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 8337 3076 8657 36908 0 FreeSans 1280 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 22644 3076 22964 36908 0 FreeSans 1280 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 36951 3076 37271 36908 0 FreeSans 1280 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 51258 3076 51578 36908 0 FreeSans 1280 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 15490 3076 15810 36908 0 FreeSans 1280 90 0 0 vss
port 2 nsew ground bidirectional
flabel metal4 s 29797 3076 30117 36908 0 FreeSans 1280 90 0 0 vss
port 2 nsew ground bidirectional
flabel metal4 s 44104 3076 44424 36908 0 FreeSans 1280 90 0 0 vss
port 2 nsew ground bidirectional
flabel metal4 s 58411 3076 58731 36908 0 FreeSans 1280 90 0 0 vss
port 2 nsew ground bidirectional
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 wb_clk_i
port 3 nsew signal input
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 wb_rst_i
port 4 nsew signal input
flabel metal2 s 56896 0 57008 800 0 FreeSans 448 90 0 0 wbs_ack_o
port 5 nsew signal tristate
flabel metal2 s 47040 0 47152 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 6 nsew signal input
flabel metal2 s 51968 0 52080 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 7 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 8 nsew signal input
flabel metal3 s 0 37184 800 37296 0 FreeSans 448 0 0 0 wbs_dat_i[0]
port 9 nsew signal input
flabel metal3 s 0 25984 800 26096 0 FreeSans 448 0 0 0 wbs_dat_i[10]
port 10 nsew signal input
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 wbs_dat_i[11]
port 11 nsew signal input
flabel metal3 s 0 23744 800 23856 0 FreeSans 448 0 0 0 wbs_dat_i[12]
port 12 nsew signal input
flabel metal3 s 0 22624 800 22736 0 FreeSans 448 0 0 0 wbs_dat_i[13]
port 13 nsew signal input
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 wbs_dat_i[14]
port 14 nsew signal input
flabel metal3 s 0 20384 800 20496 0 FreeSans 448 0 0 0 wbs_dat_i[15]
port 15 nsew signal input
flabel metal3 s 0 19264 800 19376 0 FreeSans 448 0 0 0 wbs_dat_i[16]
port 16 nsew signal input
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 wbs_dat_i[17]
port 17 nsew signal input
flabel metal3 s 0 17024 800 17136 0 FreeSans 448 0 0 0 wbs_dat_i[18]
port 18 nsew signal input
flabel metal3 s 0 15904 800 16016 0 FreeSans 448 0 0 0 wbs_dat_i[19]
port 19 nsew signal input
flabel metal3 s 0 36064 800 36176 0 FreeSans 448 0 0 0 wbs_dat_i[1]
port 20 nsew signal input
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 wbs_dat_i[20]
port 21 nsew signal input
flabel metal3 s 0 13664 800 13776 0 FreeSans 448 0 0 0 wbs_dat_i[21]
port 22 nsew signal input
flabel metal3 s 0 12544 800 12656 0 FreeSans 448 0 0 0 wbs_dat_i[22]
port 23 nsew signal input
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 wbs_dat_i[23]
port 24 nsew signal input
flabel metal3 s 0 10304 800 10416 0 FreeSans 448 0 0 0 wbs_dat_i[24]
port 25 nsew signal input
flabel metal3 s 0 9184 800 9296 0 FreeSans 448 0 0 0 wbs_dat_i[25]
port 26 nsew signal input
flabel metal3 s 0 8064 800 8176 0 FreeSans 448 0 0 0 wbs_dat_i[26]
port 27 nsew signal input
flabel metal3 s 0 6944 800 7056 0 FreeSans 448 0 0 0 wbs_dat_i[27]
port 28 nsew signal input
flabel metal3 s 0 5824 800 5936 0 FreeSans 448 0 0 0 wbs_dat_i[28]
port 29 nsew signal input
flabel metal3 s 0 4704 800 4816 0 FreeSans 448 0 0 0 wbs_dat_i[29]
port 30 nsew signal input
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 wbs_dat_i[2]
port 31 nsew signal input
flabel metal3 s 0 3584 800 3696 0 FreeSans 448 0 0 0 wbs_dat_i[30]
port 32 nsew signal input
flabel metal3 s 0 2464 800 2576 0 FreeSans 448 0 0 0 wbs_dat_i[31]
port 33 nsew signal input
flabel metal3 s 0 33824 800 33936 0 FreeSans 448 0 0 0 wbs_dat_i[3]
port 34 nsew signal input
flabel metal3 s 0 32704 800 32816 0 FreeSans 448 0 0 0 wbs_dat_i[4]
port 35 nsew signal input
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 wbs_dat_i[5]
port 36 nsew signal input
flabel metal3 s 0 30464 800 30576 0 FreeSans 448 0 0 0 wbs_dat_i[6]
port 37 nsew signal input
flabel metal3 s 0 29344 800 29456 0 FreeSans 448 0 0 0 wbs_dat_i[7]
port 38 nsew signal input
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 wbs_dat_i[8]
port 39 nsew signal input
flabel metal3 s 0 27104 800 27216 0 FreeSans 448 0 0 0 wbs_dat_i[9]
port 40 nsew signal input
flabel metal2 s 27328 0 27440 800 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 41 nsew signal input
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 42 nsew signal input
flabel metal2 s 37184 0 37296 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 43 nsew signal input
flabel metal2 s 42112 0 42224 800 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 44 nsew signal input
flabel metal2 s 12544 0 12656 800 0 FreeSans 448 90 0 0 wbs_stb_i
port 45 nsew signal input
flabel metal2 s 22400 0 22512 800 0 FreeSans 448 90 0 0 wbs_we_i
port 46 nsew signal input
flabel metal2 s 18592 39200 18704 40000 0 FreeSans 448 90 0 0 x_end[0]
port 47 nsew signal tristate
flabel metal2 s 16352 39200 16464 40000 0 FreeSans 448 90 0 0 x_end[1]
port 48 nsew signal tristate
flabel metal2 s 14112 39200 14224 40000 0 FreeSans 448 90 0 0 x_end[2]
port 49 nsew signal tristate
flabel metal2 s 11872 39200 11984 40000 0 FreeSans 448 90 0 0 x_end[3]
port 50 nsew signal tristate
flabel metal2 s 9632 39200 9744 40000 0 FreeSans 448 90 0 0 x_end[4]
port 51 nsew signal tristate
flabel metal2 s 7392 39200 7504 40000 0 FreeSans 448 90 0 0 x_end[5]
port 52 nsew signal tristate
flabel metal2 s 5152 39200 5264 40000 0 FreeSans 448 90 0 0 x_end[6]
port 53 nsew signal tristate
flabel metal2 s 2912 39200 3024 40000 0 FreeSans 448 90 0 0 x_end[7]
port 54 nsew signal tristate
flabel metal2 s 36512 39200 36624 40000 0 FreeSans 448 90 0 0 x_start[0]
port 55 nsew signal tristate
flabel metal2 s 34272 39200 34384 40000 0 FreeSans 448 90 0 0 x_start[1]
port 56 nsew signal tristate
flabel metal2 s 32032 39200 32144 40000 0 FreeSans 448 90 0 0 x_start[2]
port 57 nsew signal tristate
flabel metal2 s 29792 39200 29904 40000 0 FreeSans 448 90 0 0 x_start[3]
port 58 nsew signal tristate
flabel metal2 s 27552 39200 27664 40000 0 FreeSans 448 90 0 0 x_start[4]
port 59 nsew signal tristate
flabel metal2 s 25312 39200 25424 40000 0 FreeSans 448 90 0 0 x_start[5]
port 60 nsew signal tristate
flabel metal2 s 23072 39200 23184 40000 0 FreeSans 448 90 0 0 x_start[6]
port 61 nsew signal tristate
flabel metal2 s 20832 39200 20944 40000 0 FreeSans 448 90 0 0 x_start[7]
port 62 nsew signal tristate
flabel metal2 s 54432 39200 54544 40000 0 FreeSans 448 90 0 0 y[0]
port 63 nsew signal input
flabel metal2 s 52192 39200 52304 40000 0 FreeSans 448 90 0 0 y[1]
port 64 nsew signal input
flabel metal2 s 49952 39200 50064 40000 0 FreeSans 448 90 0 0 y[2]
port 65 nsew signal input
flabel metal2 s 47712 39200 47824 40000 0 FreeSans 448 90 0 0 y[3]
port 66 nsew signal input
flabel metal2 s 45472 39200 45584 40000 0 FreeSans 448 90 0 0 y[4]
port 67 nsew signal input
flabel metal2 s 43232 39200 43344 40000 0 FreeSans 448 90 0 0 y[5]
port 68 nsew signal input
flabel metal2 s 40992 39200 41104 40000 0 FreeSans 448 90 0 0 y[6]
port 69 nsew signal input
flabel metal2 s 38752 39200 38864 40000 0 FreeSans 448 90 0 0 y[7]
port 70 nsew signal input
rlabel metal1 29960 36848 29960 36848 0 vdd
rlabel via1 30037 36064 30037 36064 0 vss
rlabel metal3 47656 36344 47656 36344 0 _0000_
rlabel metal2 33208 35336 33208 35336 0 _0001_
rlabel metal2 29736 35168 29736 35168 0 _0002_
rlabel metal2 28392 35560 28392 35560 0 _0003_
rlabel metal2 27272 35168 27272 35168 0 _0004_
rlabel metal2 19096 35168 19096 35168 0 _0005_
rlabel metal2 13608 33600 13608 33600 0 _0006_
rlabel metal2 16800 33432 16800 33432 0 _0007_
rlabel metal2 16072 35392 16072 35392 0 _0008_
rlabel metal2 13832 35168 13832 35168 0 _0009_
rlabel metal2 12152 35056 12152 35056 0 _0010_
rlabel metal2 9912 34552 9912 34552 0 _0011_
rlabel metal2 7896 35336 7896 35336 0 _0012_
rlabel metal2 4984 35840 4984 35840 0 _0013_
rlabel metal2 2632 34328 2632 34328 0 _0014_
rlabel metal2 7000 34552 7000 34552 0 _0015_
rlabel metal2 2464 16184 2464 16184 0 _0016_
rlabel metal2 3864 17024 3864 17024 0 _0017_
rlabel metal3 10472 12824 10472 12824 0 _0018_
rlabel metal2 2520 7896 2520 7896 0 _0019_
rlabel metal2 4984 3808 4984 3808 0 _0020_
rlabel metal2 11480 3864 11480 3864 0 _0021_
rlabel metal3 28336 3416 28336 3416 0 _0022_
rlabel metal2 19096 3864 19096 3864 0 _0023_
rlabel metal2 2632 6888 2632 6888 0 _0024_
rlabel metal2 18200 9072 18200 9072 0 _0025_
rlabel metal2 9800 8960 9800 8960 0 _0026_
rlabel metal2 10584 10080 10584 10080 0 _0027_
rlabel metal3 13104 15176 13104 15176 0 _0028_
rlabel metal2 2520 15148 2520 15148 0 _0029_
rlabel metal2 2800 11144 2800 11144 0 _0030_
rlabel metal2 3304 10920 3304 10920 0 _0031_
rlabel metal2 2464 9912 2464 9912 0 _0032_
rlabel metal2 8736 6664 8736 6664 0 _0033_
rlabel metal2 12376 12936 12376 12936 0 _0034_
rlabel metal2 10360 9352 10360 9352 0 _0035_
rlabel metal2 6440 19824 6440 19824 0 _0036_
rlabel metal2 15064 12096 15064 12096 0 _0037_
rlabel metal2 17528 11144 17528 11144 0 _0038_
rlabel metal2 15624 16296 15624 16296 0 _0039_
rlabel metal2 18088 12936 18088 12936 0 _0040_
rlabel metal2 16520 13496 16520 13496 0 _0041_
rlabel metal2 16744 16072 16744 16072 0 _0042_
rlabel metal2 18200 17024 18200 17024 0 _0043_
rlabel metal2 14728 18592 14728 18592 0 _0044_
rlabel metal2 2520 18872 2520 18872 0 _0045_
rlabel metal2 6608 24024 6608 24024 0 _0046_
rlabel metal2 6440 26712 6440 26712 0 _0047_
rlabel metal2 6048 22456 6048 22456 0 _0048_
rlabel metal2 5768 29008 5768 29008 0 _0049_
rlabel metal2 7504 29960 7504 29960 0 _0050_
rlabel metal2 4424 29960 4424 29960 0 _0051_
rlabel metal2 10752 30296 10752 30296 0 _0052_
rlabel metal3 37520 16856 37520 16856 0 _0053_
rlabel metal2 37464 15624 37464 15624 0 _0054_
rlabel metal2 38248 17696 38248 17696 0 _0055_
rlabel metal3 37016 19320 37016 19320 0 _0056_
rlabel metal2 11144 25032 11144 25032 0 _0057_
rlabel metal2 11256 26600 11256 26600 0 _0058_
rlabel metal2 12152 28168 12152 28168 0 _0059_
rlabel metal2 10472 29008 10472 29008 0 _0060_
rlabel metal2 3304 20440 3304 20440 0 _0061_
rlabel metal2 3192 25144 3192 25144 0 _0062_
rlabel metal2 3080 26684 3080 26684 0 _0063_
rlabel metal2 3080 22736 3080 22736 0 _0064_
rlabel metal2 3080 28952 3080 28952 0 _0065_
rlabel metal2 2520 32984 2520 32984 0 _0066_
rlabel metal2 4088 31976 4088 31976 0 _0067_
rlabel metal3 10024 32760 10024 32760 0 _0068_
rlabel metal3 22680 20216 22680 20216 0 _0069_
rlabel metal2 11256 21000 11256 21000 0 _0070_
rlabel metal2 15064 20328 15064 20328 0 _0071_
rlabel metal3 16800 20888 16800 20888 0 _0072_
rlabel metal2 18200 22568 18200 22568 0 _0073_
rlabel metal2 20272 21448 20272 21448 0 _0074_
rlabel metal2 14056 23576 14056 23576 0 _0075_
rlabel metal2 11032 22736 11032 22736 0 _0076_
rlabel metal2 48496 17640 48496 17640 0 _0077_
rlabel metal2 49784 21616 49784 21616 0 _0078_
rlabel metal2 49560 7504 49560 7504 0 _0079_
rlabel metal2 19544 19040 19544 19040 0 _0080_
rlabel metal3 48160 16744 48160 16744 0 _0081_
rlabel metal2 49560 7000 49560 7000 0 _0082_
rlabel metal2 49336 6384 49336 6384 0 _0083_
rlabel metal3 20272 22232 20272 22232 0 _0084_
rlabel metal2 44968 20440 44968 20440 0 _0085_
rlabel metal2 48832 5880 48832 5880 0 _0086_
rlabel metal2 49784 5376 49784 5376 0 _0087_
rlabel metal3 47432 5880 47432 5880 0 _0088_
rlabel metal3 48832 5768 48832 5768 0 _0089_
rlabel metal2 49000 5488 49000 5488 0 _0090_
rlabel metal2 51016 4984 51016 4984 0 _0091_
rlabel metal3 51744 6664 51744 6664 0 _0092_
rlabel metal2 51912 6440 51912 6440 0 _0093_
rlabel metal3 21280 18984 21280 18984 0 _0094_
rlabel metal3 38640 7224 38640 7224 0 _0095_
rlabel metal2 52920 20048 52920 20048 0 _0096_
rlabel metal3 46648 20104 46648 20104 0 _0097_
rlabel metal3 51072 19320 51072 19320 0 _0098_
rlabel metal3 43960 22064 43960 22064 0 _0099_
rlabel metal3 52360 19208 52360 19208 0 _0100_
rlabel metal2 53648 16408 53648 16408 0 _0101_
rlabel metal2 53592 6384 53592 6384 0 _0102_
rlabel metal3 53592 6552 53592 6552 0 _0103_
rlabel metal2 52248 4704 52248 4704 0 _0104_
rlabel metal2 51464 5320 51464 5320 0 _0105_
rlabel metal3 49504 5096 49504 5096 0 _0106_
rlabel metal2 46424 8288 46424 8288 0 _0107_
rlabel metal2 47432 8680 47432 8680 0 _0108_
rlabel metal2 45248 9240 45248 9240 0 _0109_
rlabel metal3 45808 8008 45808 8008 0 _0110_
rlabel metal2 46536 8456 46536 8456 0 _0111_
rlabel metal2 48552 7000 48552 7000 0 _0112_
rlabel metal2 49224 4984 49224 4984 0 _0113_
rlabel metal2 51912 4424 51912 4424 0 _0114_
rlabel metal2 56952 5152 56952 5152 0 _0115_
rlabel metal2 54264 5320 54264 5320 0 _0116_
rlabel metal2 54432 5096 54432 5096 0 _0117_
rlabel metal2 55832 5544 55832 5544 0 _0118_
rlabel metal2 54376 7056 54376 7056 0 _0119_
rlabel metal2 54936 7728 54936 7728 0 _0120_
rlabel metal2 57176 7448 57176 7448 0 _0121_
rlabel metal2 36904 24640 36904 24640 0 _0122_
rlabel metal2 47432 20216 47432 20216 0 _0123_
rlabel metal2 46200 20776 46200 20776 0 _0124_
rlabel metal2 55944 19768 55944 19768 0 _0125_
rlabel metal2 53200 19432 53200 19432 0 _0126_
rlabel metal2 52304 19432 52304 19432 0 _0127_
rlabel metal2 55944 20552 55944 20552 0 _0128_
rlabel metal3 52416 20776 52416 20776 0 _0129_
rlabel metal2 49224 20776 49224 20776 0 _0130_
rlabel metal2 52920 20608 52920 20608 0 _0131_
rlabel metal2 53144 20496 53144 20496 0 _0132_
rlabel metal2 53704 20888 53704 20888 0 _0133_
rlabel metal2 56168 20552 56168 20552 0 _0134_
rlabel metal2 56616 19768 56616 19768 0 _0135_
rlabel metal2 57456 19432 57456 19432 0 _0136_
rlabel metal2 57624 6216 57624 6216 0 _0137_
rlabel metal3 57400 5880 57400 5880 0 _0138_
rlabel metal2 44072 8736 44072 8736 0 _0139_
rlabel metal2 40376 9576 40376 9576 0 _0140_
rlabel metal2 55720 6104 55720 6104 0 _0141_
rlabel metal2 57848 6272 57848 6272 0 _0142_
rlabel metal3 56168 8232 56168 8232 0 _0143_
rlabel metal2 58072 7560 58072 7560 0 _0144_
rlabel metal2 57176 9128 57176 9128 0 _0145_
rlabel metal2 57904 11480 57904 11480 0 _0146_
rlabel metal2 55496 20720 55496 20720 0 _0147_
rlabel metal2 55720 20132 55720 20132 0 _0148_
rlabel metal2 56896 20776 56896 20776 0 _0149_
rlabel metal2 54264 20608 54264 20608 0 _0150_
rlabel metal2 55720 22064 55720 22064 0 _0151_
rlabel metal2 50288 22344 50288 22344 0 _0152_
rlabel metal2 52248 22232 52248 22232 0 _0153_
rlabel metal3 52248 22120 52248 22120 0 _0154_
rlabel metal3 54824 21672 54824 21672 0 _0155_
rlabel metal2 56112 22568 56112 22568 0 _0156_
rlabel metal2 26152 21896 26152 21896 0 _0157_
rlabel metal2 54264 22624 54264 22624 0 _0158_
rlabel metal2 47208 23464 47208 23464 0 _0159_
rlabel via2 48552 23016 48552 23016 0 _0160_
rlabel metal2 54488 22736 54488 22736 0 _0161_
rlabel metal2 56728 22792 56728 22792 0 _0162_
rlabel metal2 57288 22176 57288 22176 0 _0163_
rlabel metal3 56336 21560 56336 21560 0 _0164_
rlabel metal2 56280 9744 56280 9744 0 _0165_
rlabel metal2 41776 11144 41776 11144 0 _0166_
rlabel metal2 39984 10024 39984 10024 0 _0167_
rlabel metal2 35168 21784 35168 21784 0 _0168_
rlabel metal2 40152 10248 40152 10248 0 _0169_
rlabel metal2 38920 22344 38920 22344 0 _0170_
rlabel metal2 53984 21112 53984 21112 0 _0171_
rlabel metal2 57848 21840 57848 21840 0 _0172_
rlabel metal2 57960 29456 57960 29456 0 _0173_
rlabel metal3 47432 23688 47432 23688 0 _0174_
rlabel metal3 51240 23128 51240 23128 0 _0175_
rlabel metal3 53536 28616 53536 28616 0 _0176_
rlabel metal3 48440 26600 48440 26600 0 _0177_
rlabel metal2 51912 28392 51912 28392 0 _0178_
rlabel metal2 55608 21952 55608 21952 0 _0179_
rlabel metal2 55720 24136 55720 24136 0 _0180_
rlabel metal2 55384 27832 55384 27832 0 _0181_
rlabel metal2 51296 22344 51296 22344 0 _0182_
rlabel metal2 51912 22624 51912 22624 0 _0183_
rlabel metal2 51576 22120 51576 22120 0 _0184_
rlabel metal2 36344 21840 36344 21840 0 _0185_
rlabel metal2 41384 21896 41384 21896 0 _0186_
rlabel metal2 40656 22120 40656 22120 0 _0187_
rlabel metal2 40488 21504 40488 21504 0 _0188_
rlabel metal2 43344 22456 43344 22456 0 _0189_
rlabel metal2 51632 26152 51632 26152 0 _0190_
rlabel metal2 49112 24696 49112 24696 0 _0191_
rlabel metal2 48552 24080 48552 24080 0 _0192_
rlabel metal2 47880 25088 47880 25088 0 _0193_
rlabel metal2 51912 26992 51912 26992 0 _0194_
rlabel metal2 52136 27440 52136 27440 0 _0195_
rlabel metal3 54096 27832 54096 27832 0 _0196_
rlabel metal2 54600 28336 54600 28336 0 _0197_
rlabel metal2 55832 29792 55832 29792 0 _0198_
rlabel metal2 54712 30296 54712 30296 0 _0199_
rlabel metal2 57680 10472 57680 10472 0 _0200_
rlabel metal2 55888 8456 55888 8456 0 _0201_
rlabel metal2 54936 31808 54936 31808 0 _0202_
rlabel metal3 34356 26824 34356 26824 0 _0203_
rlabel metal2 28056 24920 28056 24920 0 _0204_
rlabel metal2 29176 24920 29176 24920 0 _0205_
rlabel metal3 28560 25480 28560 25480 0 _0206_
rlabel metal2 28504 32424 28504 32424 0 _0207_
rlabel metal2 57568 29736 57568 29736 0 _0208_
rlabel metal2 56728 30240 56728 30240 0 _0209_
rlabel metal2 56392 29400 56392 29400 0 _0210_
rlabel metal2 57736 29680 57736 29680 0 _0211_
rlabel metal2 53704 31136 53704 31136 0 _0212_
rlabel metal2 54376 28168 54376 28168 0 _0213_
rlabel metal2 54824 26152 54824 26152 0 _0214_
rlabel metal2 51576 29400 51576 29400 0 _0215_
rlabel metal2 51912 27608 51912 27608 0 _0216_
rlabel metal2 50680 27552 50680 27552 0 _0217_
rlabel metal2 41048 21840 41048 21840 0 _0218_
rlabel metal2 41608 22288 41608 22288 0 _0219_
rlabel metal2 41048 23352 41048 23352 0 _0220_
rlabel metal2 39144 21840 39144 21840 0 _0221_
rlabel metal3 42112 21448 42112 21448 0 _0222_
rlabel metal2 38696 22344 38696 22344 0 _0223_
rlabel metal2 40936 23688 40936 23688 0 _0224_
rlabel metal3 42392 24808 42392 24808 0 _0225_
rlabel metal2 41272 24304 41272 24304 0 _0226_
rlabel metal2 42616 25200 42616 25200 0 _0227_
rlabel metal2 38472 23296 38472 23296 0 _0228_
rlabel metal2 38808 25200 38808 25200 0 _0229_
rlabel metal2 42448 24696 42448 24696 0 _0230_
rlabel metal2 50904 27720 50904 27720 0 _0231_
rlabel metal2 51576 28280 51576 28280 0 _0232_
rlabel metal2 49784 28392 49784 28392 0 _0233_
rlabel metal2 53368 29680 53368 29680 0 _0234_
rlabel metal2 49448 29064 49448 29064 0 _0235_
rlabel metal3 43064 24864 43064 24864 0 _0236_
rlabel metal2 48216 24640 48216 24640 0 _0237_
rlabel metal2 48832 24584 48832 24584 0 _0238_
rlabel metal2 47208 27048 47208 27048 0 _0239_
rlabel metal2 46984 27496 46984 27496 0 _0240_
rlabel metal2 48216 28280 48216 28280 0 _0241_
rlabel metal2 49224 29512 49224 29512 0 _0242_
rlabel metal3 53816 29400 53816 29400 0 _0243_
rlabel metal2 53816 30240 53816 30240 0 _0244_
rlabel metal2 55272 31304 55272 31304 0 _0245_
rlabel metal2 56392 36288 56392 36288 0 _0246_
rlabel metal2 27944 33712 27944 33712 0 _0247_
rlabel metal2 28280 34552 28280 34552 0 _0248_
rlabel metal2 29064 32536 29064 32536 0 _0249_
rlabel metal3 29120 33432 29120 33432 0 _0250_
rlabel metal2 56616 31416 56616 31416 0 _0251_
rlabel metal2 50904 32200 50904 32200 0 _0252_
rlabel metal2 51688 30240 51688 30240 0 _0253_
rlabel metal2 48104 31584 48104 31584 0 _0254_
rlabel metal2 48104 30240 48104 30240 0 _0255_
rlabel metal2 49112 29120 49112 29120 0 _0256_
rlabel metal3 48552 31752 48552 31752 0 _0257_
rlabel metal2 43512 30072 43512 30072 0 _0258_
rlabel metal2 42280 26096 42280 26096 0 _0259_
rlabel metal2 16744 21056 16744 21056 0 _0260_
rlabel metal2 29568 23128 29568 23128 0 _0261_
rlabel metal3 32312 21560 32312 21560 0 _0262_
rlabel metal2 32424 22064 32424 22064 0 _0263_
rlabel metal2 33432 21728 33432 21728 0 _0264_
rlabel metal2 33040 21560 33040 21560 0 _0265_
rlabel metal2 32648 23128 32648 23128 0 _0266_
rlabel metal3 32816 24696 32816 24696 0 _0267_
rlabel metal3 22176 22120 22176 22120 0 _0268_
rlabel metal3 32592 23800 32592 23800 0 _0269_
rlabel metal2 15512 21616 15512 21616 0 _0270_
rlabel metal2 35560 23688 35560 23688 0 _0271_
rlabel metal3 32704 23912 32704 23912 0 _0272_
rlabel metal2 32816 24696 32816 24696 0 _0273_
rlabel metal2 42000 25480 42000 25480 0 _0274_
rlabel metal2 42504 31304 42504 31304 0 _0275_
rlabel metal3 46928 27832 46928 27832 0 _0276_
rlabel metal2 47376 27272 47376 27272 0 _0277_
rlabel metal2 41272 27888 41272 27888 0 _0278_
rlabel metal3 38696 24808 38696 24808 0 _0279_
rlabel metal2 39144 24976 39144 24976 0 _0280_
rlabel metal3 39424 24584 39424 24584 0 _0281_
rlabel metal2 39816 27720 39816 27720 0 _0282_
rlabel metal2 15960 25200 15960 25200 0 _0283_
rlabel metal2 34328 27384 34328 27384 0 _0284_
rlabel metal2 16744 24304 16744 24304 0 _0285_
rlabel metal2 33768 27384 33768 27384 0 _0286_
rlabel metal3 36960 27832 36960 27832 0 _0287_
rlabel metal3 40600 28616 40600 28616 0 _0288_
rlabel metal3 43344 30968 43344 30968 0 _0289_
rlabel metal2 46648 32200 46648 32200 0 _0290_
rlabel metal2 50120 30520 50120 30520 0 _0291_
rlabel metal3 43736 32816 43736 32816 0 _0292_
rlabel metal2 45640 31864 45640 31864 0 _0293_
rlabel metal2 29792 32760 29792 32760 0 _0294_
rlabel metal3 28504 34328 28504 34328 0 _0295_
rlabel metal3 16856 16856 16856 16856 0 _0296_
rlabel metal2 46424 30296 46424 30296 0 _0297_
rlabel metal3 48160 31976 48160 31976 0 _0298_
rlabel metal2 20216 32872 20216 32872 0 _0299_
rlabel metal2 46760 31696 46760 31696 0 _0300_
rlabel metal3 42308 31080 42308 31080 0 _0301_
rlabel metal2 43008 30296 43008 30296 0 _0302_
rlabel metal2 44296 30576 44296 30576 0 _0303_
rlabel metal3 39816 30240 39816 30240 0 _0304_
rlabel metal2 39928 28280 39928 28280 0 _0305_
rlabel metal3 40600 27944 40600 27944 0 _0306_
rlabel metal3 39928 28056 39928 28056 0 _0307_
rlabel metal3 38668 28392 38668 28392 0 _0308_
rlabel metal2 43848 27552 43848 27552 0 _0309_
rlabel metal2 32200 27832 32200 27832 0 _0310_
rlabel metal2 32256 24920 32256 24920 0 _0311_
rlabel metal2 31192 22624 31192 22624 0 _0312_
rlabel metal2 26824 23716 26824 23716 0 _0313_
rlabel metal2 25928 21840 25928 21840 0 _0314_
rlabel metal3 24920 22120 24920 22120 0 _0315_
rlabel metal2 26824 21952 26824 21952 0 _0316_
rlabel metal2 27776 23240 27776 23240 0 _0317_
rlabel metal3 30464 25480 30464 25480 0 _0318_
rlabel metal2 31584 25592 31584 25592 0 _0319_
rlabel metal3 31976 26264 31976 26264 0 _0320_
rlabel metal2 34440 27328 34440 27328 0 _0321_
rlabel metal2 28504 26628 28504 26628 0 _0322_
rlabel metal2 35896 23408 35896 23408 0 _0323_
rlabel metal2 25480 27720 25480 27720 0 _0324_
rlabel metal2 23576 26628 23576 26628 0 _0325_
rlabel metal2 24304 26488 24304 26488 0 _0326_
rlabel metal3 25312 26936 25312 26936 0 _0327_
rlabel metal2 26040 27440 26040 27440 0 _0328_
rlabel metal2 31080 26572 31080 26572 0 _0329_
rlabel metal2 30296 28616 30296 28616 0 _0330_
rlabel metal2 29512 30296 29512 30296 0 _0331_
rlabel metal2 20328 31584 20328 31584 0 _0332_
rlabel metal2 17752 33768 17752 33768 0 _0333_
rlabel metal2 15176 19376 15176 19376 0 _0334_
rlabel metal3 17696 31752 17696 31752 0 _0335_
rlabel metal2 19600 31752 19600 31752 0 _0336_
rlabel metal2 14728 32368 14728 32368 0 _0337_
rlabel metal3 28896 30856 28896 30856 0 _0338_
rlabel metal2 29176 30576 29176 30576 0 _0339_
rlabel metal2 14840 31472 14840 31472 0 _0340_
rlabel metal2 31752 27832 31752 27832 0 _0341_
rlabel metal2 30632 28672 30632 28672 0 _0342_
rlabel metal2 30520 28840 30520 28840 0 _0343_
rlabel metal2 14728 29624 14728 29624 0 _0344_
rlabel metal3 24976 27720 24976 27720 0 _0345_
rlabel metal2 25872 27832 25872 27832 0 _0346_
rlabel metal2 28336 27720 28336 27720 0 _0347_
rlabel metal3 28616 27664 28616 27664 0 _0348_
rlabel metal2 15736 27160 15736 27160 0 _0349_
rlabel metal2 32424 26544 32424 26544 0 _0350_
rlabel metal2 16408 26376 16408 26376 0 _0351_
rlabel metal2 23688 25032 23688 25032 0 _0352_
rlabel metal2 24136 25480 24136 25480 0 _0353_
rlabel metal3 21728 24696 21728 24696 0 _0354_
rlabel metal2 25928 22176 25928 22176 0 _0355_
rlabel metal2 19768 24528 19768 24528 0 _0356_
rlabel metal2 19488 25480 19488 25480 0 _0357_
rlabel metal3 19264 26824 19264 26824 0 _0358_
rlabel metal2 18760 25928 18760 25928 0 _0359_
rlabel metal2 18312 24808 18312 24808 0 _0360_
rlabel metal3 19040 26152 19040 26152 0 _0361_
rlabel metal2 28168 23912 28168 23912 0 _0362_
rlabel metal2 25368 23408 25368 23408 0 _0363_
rlabel metal2 25872 22344 25872 22344 0 _0364_
rlabel metal2 26264 22344 26264 22344 0 _0365_
rlabel metal2 27272 22624 27272 22624 0 _0366_
rlabel metal2 25368 24640 25368 24640 0 _0367_
rlabel metal2 21336 25872 21336 25872 0 _0368_
rlabel metal2 15176 27944 15176 27944 0 _0369_
rlabel metal2 14896 29288 14896 29288 0 _0370_
rlabel metal2 15736 31136 15736 31136 0 _0371_
rlabel metal3 13776 31752 13776 31752 0 _0372_
rlabel metal2 13048 32760 13048 32760 0 _0373_
rlabel metal2 15176 32480 15176 32480 0 _0374_
rlabel metal2 16184 31808 16184 31808 0 _0375_
rlabel metal2 15288 33040 15288 33040 0 _0376_
rlabel metal2 15512 30856 15512 30856 0 _0377_
rlabel metal2 14952 30688 14952 30688 0 _0378_
rlabel metal2 16072 26236 16072 26236 0 _0379_
rlabel metal2 16184 27160 16184 27160 0 _0380_
rlabel metal2 15624 27552 15624 27552 0 _0381_
rlabel metal3 18872 27832 18872 27832 0 _0382_
rlabel metal3 19768 27384 19768 27384 0 _0383_
rlabel metal2 20104 27552 20104 27552 0 _0384_
rlabel metal3 20160 27720 20160 27720 0 _0385_
rlabel metal3 16912 27720 16912 27720 0 _0386_
rlabel metal2 21448 25032 21448 25032 0 _0387_
rlabel metal3 24920 23688 24920 23688 0 _0388_
rlabel metal2 24360 24416 24360 24416 0 _0389_
rlabel metal2 21448 25816 21448 25816 0 _0390_
rlabel metal2 19768 23744 19768 23744 0 _0391_
rlabel metal2 19040 23800 19040 23800 0 _0392_
rlabel metal3 20552 24024 20552 24024 0 _0393_
rlabel metal2 24136 22792 24136 22792 0 _0394_
rlabel metal2 31416 23520 31416 23520 0 _0395_
rlabel metal2 24472 23296 24472 23296 0 _0396_
rlabel metal2 23520 23240 23520 23240 0 _0397_
rlabel metal2 23072 24808 23072 24808 0 _0398_
rlabel metal2 22904 25032 22904 25032 0 _0399_
rlabel metal2 16464 28056 16464 28056 0 _0400_
rlabel metal2 14952 32256 14952 32256 0 _0401_
rlabel metal2 15736 33768 15736 33768 0 _0402_
rlabel metal3 55440 36176 55440 36176 0 _0403_
rlabel metal2 11816 17584 11816 17584 0 _0404_
rlabel metal2 12152 16632 12152 16632 0 _0405_
rlabel metal2 11088 2296 11088 2296 0 _0406_
rlabel metal2 10696 10528 10696 10528 0 _0407_
rlabel metal3 9912 10024 9912 10024 0 _0408_
rlabel metal3 5208 18424 5208 18424 0 _0409_
rlabel metal2 4200 18648 4200 18648 0 _0410_
rlabel metal3 9856 8904 9856 8904 0 _0411_
rlabel metal3 9240 16968 9240 16968 0 _0412_
rlabel metal2 10808 16632 10808 16632 0 _0413_
rlabel metal2 10584 18872 10584 18872 0 _0414_
rlabel metal2 10136 15960 10136 15960 0 _0415_
rlabel metal2 11256 14616 11256 14616 0 _0416_
rlabel metal2 11592 14056 11592 14056 0 _0417_
rlabel metal3 11816 14392 11816 14392 0 _0418_
rlabel metal2 11704 19712 11704 19712 0 _0419_
rlabel metal2 11368 16128 11368 16128 0 _0420_
rlabel metal2 11760 15288 11760 15288 0 _0421_
rlabel metal2 18984 19600 18984 19600 0 _0422_
rlabel metal3 13944 16856 13944 16856 0 _0423_
rlabel metal2 2520 12152 2520 12152 0 _0424_
rlabel metal2 2576 13832 2576 13832 0 _0425_
rlabel metal2 4200 14784 4200 14784 0 _0426_
rlabel metal2 3304 13496 3304 13496 0 _0427_
rlabel metal2 7784 17304 7784 17304 0 _0428_
rlabel metal2 3080 11424 3080 11424 0 _0429_
rlabel metal2 3080 13216 3080 13216 0 _0430_
rlabel metal2 2128 11592 2128 11592 0 _0431_
rlabel metal2 9240 11984 9240 11984 0 _0432_
rlabel metal3 13272 13720 13272 13720 0 _0433_
rlabel metal2 12600 16296 12600 16296 0 _0434_
rlabel metal2 10696 12600 10696 12600 0 _0435_
rlabel metal2 16856 15148 16856 15148 0 _0436_
rlabel metal2 2744 19544 2744 19544 0 _0437_
rlabel metal3 24640 13496 24640 13496 0 _0438_
rlabel metal2 8848 20888 8848 20888 0 _0439_
rlabel metal2 7560 18872 7560 18872 0 _0440_
rlabel metal2 7224 19264 7224 19264 0 _0441_
rlabel metal3 9800 18424 9800 18424 0 _0442_
rlabel metal2 15400 17192 15400 17192 0 _0443_
rlabel metal2 15848 13160 15848 13160 0 _0444_
rlabel metal3 16128 14392 16128 14392 0 _0445_
rlabel metal2 15288 13216 15288 13216 0 _0446_
rlabel metal2 17640 12320 17640 12320 0 _0447_
rlabel metal2 16520 17360 16520 17360 0 _0448_
rlabel metal2 15064 17360 15064 17360 0 _0449_
rlabel metal2 13440 17640 13440 17640 0 _0450_
rlabel metal2 13832 17192 13832 17192 0 _0451_
rlabel metal2 17640 13888 17640 13888 0 _0452_
rlabel metal2 16296 17136 16296 17136 0 _0453_
rlabel metal2 16296 13608 16296 13608 0 _0454_
rlabel metal2 16184 16632 16184 16632 0 _0455_
rlabel metal2 14952 17696 14952 17696 0 _0456_
rlabel metal2 13048 17360 13048 17360 0 _0457_
rlabel metal2 13832 19096 13832 19096 0 _0458_
rlabel metal2 13720 19040 13720 19040 0 _0459_
rlabel metal3 9632 26936 9632 26936 0 _0460_
rlabel metal2 8680 19936 8680 19936 0 _0461_
rlabel metal2 2856 19208 2856 19208 0 _0462_
rlabel metal2 3416 18592 3416 18592 0 _0463_
rlabel metal2 4032 17752 4032 17752 0 _0464_
rlabel metal2 7056 27832 7056 27832 0 _0465_
rlabel metal2 7448 28280 7448 28280 0 _0466_
rlabel metal2 6888 23856 6888 23856 0 _0467_
rlabel metal2 6440 24192 6440 24192 0 _0468_
rlabel metal3 7616 26264 7616 26264 0 _0469_
rlabel metal2 4928 24920 4928 24920 0 _0470_
rlabel metal2 6328 23240 6328 23240 0 _0471_
rlabel metal3 5376 22232 5376 22232 0 _0472_
rlabel metal3 6384 28616 6384 28616 0 _0473_
rlabel metal3 2632 32648 2632 32648 0 _0474_
rlabel metal3 5152 28616 5152 28616 0 _0475_
rlabel metal2 6104 28840 6104 28840 0 _0476_
rlabel metal2 7896 30856 7896 30856 0 _0477_
rlabel metal2 7672 30184 7672 30184 0 _0478_
rlabel metal3 5600 30072 5600 30072 0 _0479_
rlabel metal2 4424 30632 4424 30632 0 _0480_
rlabel metal2 10584 30632 10584 30632 0 _0481_
rlabel metal3 6188 29960 6188 29960 0 _0482_
rlabel metal2 10472 19208 10472 19208 0 _0483_
rlabel metal2 9128 21168 9128 21168 0 _0484_
rlabel metal2 11928 20216 11928 20216 0 _0485_
rlabel metal2 23240 17528 23240 17528 0 _0486_
rlabel metal3 36456 16856 36456 16856 0 _0487_
rlabel metal2 11816 19992 11816 19992 0 _0488_
rlabel metal2 17976 17640 17976 17640 0 _0489_
rlabel metal2 18648 15456 18648 15456 0 _0490_
rlabel metal2 36456 16464 36456 16464 0 _0491_
rlabel metal3 36904 15960 36904 15960 0 _0492_
rlabel metal3 18088 17304 18088 17304 0 _0493_
rlabel metal2 37520 18424 37520 18424 0 _0494_
rlabel metal3 27552 2184 27552 2184 0 _0495_
rlabel metal2 36232 19544 36232 19544 0 _0496_
rlabel metal3 18088 18256 18088 18256 0 _0497_
rlabel metal2 12208 20664 12208 20664 0 _0498_
rlabel metal3 11480 25368 11480 25368 0 _0499_
rlabel metal2 10696 27496 10696 27496 0 _0500_
rlabel metal2 10808 25368 10808 25368 0 _0501_
rlabel metal2 10920 27888 10920 27888 0 _0502_
rlabel metal3 11536 27048 11536 27048 0 _0503_
rlabel metal2 10696 27048 10696 27048 0 _0504_
rlabel metal3 11760 28616 11760 28616 0 _0505_
rlabel metal2 11032 28336 11032 28336 0 _0506_
rlabel metal2 12824 28784 12824 28784 0 _0507_
rlabel metal2 10024 28840 10024 28840 0 _0508_
rlabel metal2 3192 22960 3192 22960 0 _0509_
rlabel metal2 2184 23912 2184 23912 0 _0510_
rlabel metal3 3920 19768 3920 19768 0 _0511_
rlabel metal2 4760 28112 4760 28112 0 _0512_
rlabel metal2 4144 28504 4144 28504 0 _0513_
rlabel metal2 3416 24976 3416 24976 0 _0514_
rlabel metal2 3080 24304 3080 24304 0 _0515_
rlabel metal2 3528 25536 3528 25536 0 _0516_
rlabel metal3 4648 26152 4648 26152 0 _0517_
rlabel metal2 2408 25088 2408 25088 0 _0518_
rlabel metal2 3416 22680 3416 22680 0 _0519_
rlabel metal2 2968 23016 2968 23016 0 _0520_
rlabel metal3 3528 28616 3528 28616 0 _0521_
rlabel metal3 5208 31640 5208 31640 0 _0522_
rlabel metal2 2856 29512 2856 29512 0 _0523_
rlabel metal2 2744 33264 2744 33264 0 _0524_
rlabel metal2 2408 33376 2408 33376 0 _0525_
rlabel metal3 4536 31976 4536 31976 0 _0526_
rlabel metal3 5208 32536 5208 32536 0 _0527_
rlabel metal3 5264 30184 5264 30184 0 _0528_
rlabel metal2 9576 31836 9576 31836 0 _0529_
rlabel metal2 5992 32088 5992 32088 0 _0530_
rlabel metal2 17528 20160 17528 20160 0 _0531_
rlabel metal3 18816 21672 18816 21672 0 _0532_
rlabel metal3 18536 19768 18536 19768 0 _0533_
rlabel metal3 11564 20776 11564 20776 0 _0534_
rlabel metal2 11704 21392 11704 21392 0 _0535_
rlabel metal2 15960 21840 15960 21840 0 _0536_
rlabel metal2 10920 21056 10920 21056 0 _0537_
rlabel metal2 15064 21056 15064 21056 0 _0538_
rlabel metal2 15512 20776 15512 20776 0 _0539_
rlabel metal2 15288 22512 15288 22512 0 _0540_
rlabel metal2 15288 23016 15288 23016 0 _0541_
rlabel metal3 15288 22232 15288 22232 0 _0542_
rlabel metal2 16296 22400 16296 22400 0 _0543_
rlabel metal2 15008 22344 15008 22344 0 _0544_
rlabel metal2 14728 22400 14728 22400 0 _0545_
rlabel metal2 16296 21056 16296 21056 0 _0546_
rlabel metal3 15064 23128 15064 23128 0 _0547_
rlabel metal2 13720 23184 13720 23184 0 _0548_
rlabel metal2 10920 22512 10920 22512 0 _0549_
rlabel metal2 11144 23016 11144 23016 0 _0550_
rlabel metal3 18928 3752 18928 3752 0 _0551_
rlabel metal2 29176 7952 29176 7952 0 _0552_
rlabel metal2 20552 10640 20552 10640 0 _0553_
rlabel metal2 31304 8344 31304 8344 0 _0554_
rlabel metal2 42280 10472 42280 10472 0 _0555_
rlabel metal2 39704 9408 39704 9408 0 _0556_
rlabel metal2 42616 9072 42616 9072 0 _0557_
rlabel metal2 13608 31920 13608 31920 0 _0558_
rlabel metal2 44968 34496 44968 34496 0 _0559_
rlabel metal3 14252 29400 14252 29400 0 _0560_
rlabel metal3 45976 35560 45976 35560 0 _0561_
rlabel metal2 8008 28224 8008 28224 0 _0562_
rlabel metal2 42280 35224 42280 35224 0 _0563_
rlabel metal2 44072 35336 44072 35336 0 _0564_
rlabel metal2 8904 33152 8904 33152 0 _0565_
rlabel metal2 43848 34888 43848 34888 0 _0566_
rlabel metal2 41776 20664 41776 20664 0 _0567_
rlabel metal2 19040 7560 19040 7560 0 _0568_
rlabel metal2 36456 32592 36456 32592 0 _0569_
rlabel metal2 39592 35280 39592 35280 0 _0570_
rlabel metal2 18088 34664 18088 34664 0 _0571_
rlabel metal2 39928 35616 39928 35616 0 _0572_
rlabel metal2 7392 18984 7392 18984 0 _0573_
rlabel metal3 8568 28392 8568 28392 0 _0574_
rlabel metal2 40152 35224 40152 35224 0 _0575_
rlabel metal2 8176 22568 8176 22568 0 _0576_
rlabel metal3 40656 35448 40656 35448 0 _0577_
rlabel metal2 20664 10248 20664 10248 0 _0578_
rlabel metal2 20440 4368 20440 4368 0 _0579_
rlabel metal3 18088 4424 18088 4424 0 _0580_
rlabel metal2 18536 4536 18536 4536 0 _0581_
rlabel metal2 17864 6608 17864 6608 0 _0582_
rlabel metal3 4648 6104 4648 6104 0 _0583_
rlabel metal2 19768 10640 19768 10640 0 _0584_
rlabel metal2 6776 9296 6776 9296 0 _0585_
rlabel metal2 7784 6608 7784 6608 0 _0586_
rlabel metal3 22960 10696 22960 10696 0 _0587_
rlabel metal2 25816 7000 25816 7000 0 _0588_
rlabel metal2 5992 11312 5992 11312 0 _0589_
rlabel metal2 13160 28784 13160 28784 0 _0590_
rlabel metal2 6832 30632 6832 30632 0 _0591_
rlabel metal2 4872 13160 4872 13160 0 _0592_
rlabel metal2 7448 12992 7448 12992 0 _0593_
rlabel metal2 6776 10024 6776 10024 0 _0594_
rlabel metal2 6552 13272 6552 13272 0 _0595_
rlabel metal2 5768 11032 5768 11032 0 _0596_
rlabel metal2 6328 10472 6328 10472 0 _0597_
rlabel metal2 8008 10640 8008 10640 0 _0598_
rlabel metal3 17640 8120 17640 8120 0 _0599_
rlabel metal2 20216 7280 20216 7280 0 _0600_
rlabel metal3 12824 3304 12824 3304 0 _0601_
rlabel metal2 18312 5432 18312 5432 0 _0602_
rlabel metal2 19992 7000 19992 7000 0 _0603_
rlabel metal3 10864 5992 10864 5992 0 _0604_
rlabel metal2 11144 6048 11144 6048 0 _0605_
rlabel metal3 15960 2520 15960 2520 0 _0606_
rlabel metal2 20664 6664 20664 6664 0 _0607_
rlabel metal2 33320 3976 33320 3976 0 _0608_
rlabel metal2 35784 10528 35784 10528 0 _0609_
rlabel metal2 43512 12544 43512 12544 0 _0610_
rlabel metal2 22344 4872 22344 4872 0 _0611_
rlabel metal2 24752 4424 24752 4424 0 _0612_
rlabel metal2 23352 5376 23352 5376 0 _0613_
rlabel metal2 42056 9464 42056 9464 0 _0614_
rlabel metal2 41440 15400 41440 15400 0 _0615_
rlabel metal2 46536 6608 46536 6608 0 _0616_
rlabel metal3 46088 7448 46088 7448 0 _0617_
rlabel metal2 26488 7840 26488 7840 0 _0618_
rlabel metal2 42168 9800 42168 9800 0 _0619_
rlabel metal2 44184 6720 44184 6720 0 _0620_
rlabel metal2 43288 7112 43288 7112 0 _0621_
rlabel metal2 22792 4816 22792 4816 0 _0622_
rlabel metal3 25928 4312 25928 4312 0 _0623_
rlabel metal3 18872 4200 18872 4200 0 _0624_
rlabel metal2 25256 5824 25256 5824 0 _0625_
rlabel metal2 17080 5656 17080 5656 0 _0626_
rlabel metal2 22568 5992 22568 5992 0 _0627_
rlabel metal3 15288 5152 15288 5152 0 _0628_
rlabel metal2 21672 6720 21672 6720 0 _0629_
rlabel metal2 26600 4648 26600 4648 0 _0630_
rlabel metal2 28504 3976 28504 3976 0 _0631_
rlabel metal2 33432 6552 33432 6552 0 _0632_
rlabel metal3 33208 16856 33208 16856 0 _0633_
rlabel metal2 42616 7952 42616 7952 0 _0634_
rlabel metal3 42728 9688 42728 9688 0 _0635_
rlabel metal2 46200 7728 46200 7728 0 _0636_
rlabel metal2 47656 8344 47656 8344 0 _0637_
rlabel metal2 48888 16912 48888 16912 0 _0638_
rlabel metal3 40936 15400 40936 15400 0 _0639_
rlabel metal2 48720 13832 48720 13832 0 _0640_
rlabel metal2 45752 15792 45752 15792 0 _0641_
rlabel metal2 49560 18872 49560 18872 0 _0642_
rlabel metal2 50456 15680 50456 15680 0 _0643_
rlabel metal2 48944 14280 48944 14280 0 _0644_
rlabel metal2 45472 23688 45472 23688 0 _0645_
rlabel metal2 43064 17080 43064 17080 0 _0646_
rlabel metal2 46872 17136 46872 17136 0 _0647_
rlabel metal2 48104 13664 48104 13664 0 _0648_
rlabel metal2 47040 11368 47040 11368 0 _0649_
rlabel metal2 45248 23688 45248 23688 0 _0650_
rlabel metal2 43960 14504 43960 14504 0 _0651_
rlabel metal2 49560 17528 49560 17528 0 _0652_
rlabel metal2 49504 23912 49504 23912 0 _0653_
rlabel metal2 48048 26376 48048 26376 0 _0654_
rlabel metal2 44576 18424 44576 18424 0 _0655_
rlabel metal3 44240 11256 44240 11256 0 _0656_
rlabel metal2 46704 19096 46704 19096 0 _0657_
rlabel metal2 44688 24024 44688 24024 0 _0658_
rlabel metal2 44968 14224 44968 14224 0 _0659_
rlabel metal2 45640 16800 45640 16800 0 _0660_
rlabel metal2 46704 11480 46704 11480 0 _0661_
rlabel metal2 47544 10080 47544 10080 0 _0662_
rlabel metal2 47432 9520 47432 9520 0 _0663_
rlabel metal2 47208 12152 47208 12152 0 _0664_
rlabel metal2 46984 14560 46984 14560 0 _0665_
rlabel metal2 45752 11648 45752 11648 0 _0666_
rlabel metal2 45752 11312 45752 11312 0 _0667_
rlabel metal2 45976 11256 45976 11256 0 _0668_
rlabel metal2 48720 10024 48720 10024 0 _0669_
rlabel metal2 47208 5040 47208 5040 0 _0670_
rlabel metal2 26152 11536 26152 11536 0 _0671_
rlabel metal3 33880 10584 33880 10584 0 _0672_
rlabel metal2 21448 32928 21448 32928 0 _0673_
rlabel metal3 41328 4312 41328 4312 0 _0674_
rlabel metal3 44072 7448 44072 7448 0 _0675_
rlabel metal2 42392 7728 42392 7728 0 _0676_
rlabel metal2 41496 4424 41496 4424 0 _0677_
rlabel metal3 32256 4424 32256 4424 0 _0678_
rlabel metal3 15792 8904 15792 8904 0 _0679_
rlabel metal2 18088 6384 18088 6384 0 _0680_
rlabel metal2 17752 8288 17752 8288 0 _0681_
rlabel metal2 23632 5992 23632 5992 0 _0682_
rlabel metal3 21224 2856 21224 2856 0 _0683_
rlabel metal2 26264 5488 26264 5488 0 _0684_
rlabel metal2 26712 5432 26712 5432 0 _0685_
rlabel metal2 29848 7056 29848 7056 0 _0686_
rlabel metal2 30296 13160 30296 13160 0 _0687_
rlabel metal2 30800 7224 30800 7224 0 _0688_
rlabel metal3 31864 6552 31864 6552 0 _0689_
rlabel metal2 40824 3976 40824 3976 0 _0690_
rlabel metal2 46648 4760 46648 4760 0 _0691_
rlabel metal2 47992 5376 47992 5376 0 _0692_
rlabel metal2 46480 18536 46480 18536 0 _0693_
rlabel metal2 47432 13160 47432 13160 0 _0694_
rlabel metal2 47208 18480 47208 18480 0 _0695_
rlabel metal2 40992 15960 40992 15960 0 _0696_
rlabel metal2 50232 16268 50232 16268 0 _0697_
rlabel metal2 49112 14000 49112 14000 0 _0698_
rlabel metal2 49672 14000 49672 14000 0 _0699_
rlabel metal2 49784 13384 49784 13384 0 _0700_
rlabel metal2 49224 16128 49224 16128 0 _0701_
rlabel metal2 40936 15512 40936 15512 0 _0702_
rlabel metal2 41048 18256 41048 18256 0 _0703_
rlabel metal3 47768 16184 47768 16184 0 _0704_
rlabel metal3 47600 16968 47600 16968 0 _0705_
rlabel metal3 49112 16072 49112 16072 0 _0706_
rlabel metal2 49392 11368 49392 11368 0 _0707_
rlabel metal2 51632 11592 51632 11592 0 _0708_
rlabel metal2 52584 9744 52584 9744 0 _0709_
rlabel metal2 49784 9408 49784 9408 0 _0710_
rlabel metal3 48440 8120 48440 8120 0 _0711_
rlabel metal2 47880 7728 47880 7728 0 _0712_
rlabel metal2 22792 11088 22792 11088 0 _0713_
rlabel metal2 45416 8512 45416 8512 0 _0714_
rlabel metal2 46536 9856 46536 9856 0 _0715_
rlabel metal2 44296 10696 44296 10696 0 _0716_
rlabel metal2 46200 12768 46200 12768 0 _0717_
rlabel metal3 45528 9688 45528 9688 0 _0718_
rlabel metal2 46704 9800 46704 9800 0 _0719_
rlabel metal2 46312 9856 46312 9856 0 _0720_
rlabel metal2 46536 9240 46536 9240 0 _0721_
rlabel metal2 46312 8848 46312 8848 0 _0722_
rlabel metal2 46984 9632 46984 9632 0 _0723_
rlabel metal2 49336 9072 49336 9072 0 _0724_
rlabel metal2 50008 8512 50008 8512 0 _0725_
rlabel metal2 47432 3696 47432 3696 0 _0726_
rlabel metal2 26264 12040 26264 12040 0 _0727_
rlabel metal3 33600 14280 33600 14280 0 _0728_
rlabel metal3 41272 6048 41272 6048 0 _0729_
rlabel metal3 35168 5208 35168 5208 0 _0730_
rlabel metal2 37576 5768 37576 5768 0 _0731_
rlabel metal2 30632 5656 30632 5656 0 _0732_
rlabel metal2 17864 7952 17864 7952 0 _0733_
rlabel metal2 31080 8288 31080 8288 0 _0734_
rlabel metal2 33768 7784 33768 7784 0 _0735_
rlabel metal2 31192 6496 31192 6496 0 _0736_
rlabel metal3 30296 8904 30296 8904 0 _0737_
rlabel metal2 32312 5488 32312 5488 0 _0738_
rlabel metal2 40152 4536 40152 4536 0 _0739_
rlabel metal2 28840 5824 28840 5824 0 _0740_
rlabel metal3 30968 5880 30968 5880 0 _0741_
rlabel metal2 26376 6944 26376 6944 0 _0742_
rlabel metal2 26712 8344 26712 8344 0 _0743_
rlabel metal2 18200 10304 18200 10304 0 _0744_
rlabel metal2 15176 5824 15176 5824 0 _0745_
rlabel metal2 20888 8400 20888 8400 0 _0746_
rlabel metal2 15176 4928 15176 4928 0 _0747_
rlabel metal2 21784 4592 21784 4592 0 _0748_
rlabel metal2 22792 6384 22792 6384 0 _0749_
rlabel metal3 17248 7224 17248 7224 0 _0750_
rlabel metal2 21336 7896 21336 7896 0 _0751_
rlabel metal2 24136 8736 24136 8736 0 _0752_
rlabel metal2 24304 8232 24304 8232 0 _0753_
rlabel metal2 13664 9016 13664 9016 0 _0754_
rlabel metal2 23128 8512 23128 8512 0 _0755_
rlabel metal2 24024 8512 24024 8512 0 _0756_
rlabel metal3 26236 8344 26236 8344 0 _0757_
rlabel metal2 28616 6440 28616 6440 0 _0758_
rlabel metal2 40264 4704 40264 4704 0 _0759_
rlabel metal2 43736 4816 43736 4816 0 _0760_
rlabel metal2 43064 3528 43064 3528 0 _0761_
rlabel metal2 41160 3584 41160 3584 0 _0762_
rlabel metal3 42672 5208 42672 5208 0 _0763_
rlabel metal2 46760 5936 46760 5936 0 _0764_
rlabel metal3 50176 11368 50176 11368 0 _0765_
rlabel metal2 50008 12208 50008 12208 0 _0766_
rlabel metal2 51464 7896 51464 7896 0 _0767_
rlabel metal2 49896 17248 49896 17248 0 _0768_
rlabel metal2 51464 17080 51464 17080 0 _0769_
rlabel metal2 52920 16352 52920 16352 0 _0770_
rlabel metal2 49000 16576 49000 16576 0 _0771_
rlabel metal2 49896 16576 49896 16576 0 _0772_
rlabel metal2 49112 16016 49112 16016 0 _0773_
rlabel metal2 43512 16464 43512 16464 0 _0774_
rlabel metal2 25424 5208 25424 5208 0 _0775_
rlabel metal3 45752 16072 45752 16072 0 _0776_
rlabel metal3 40376 16856 40376 16856 0 _0777_
rlabel metal2 42280 16408 42280 16408 0 _0778_
rlabel metal2 42336 15288 42336 15288 0 _0779_
rlabel metal2 43288 16240 43288 16240 0 _0780_
rlabel metal2 44184 16240 44184 16240 0 _0781_
rlabel metal2 52472 15680 52472 15680 0 _0782_
rlabel metal2 54376 9408 54376 9408 0 _0783_
rlabel metal2 53144 8120 53144 8120 0 _0784_
rlabel metal3 52416 9800 52416 9800 0 _0785_
rlabel metal2 52920 9240 52920 9240 0 _0786_
rlabel metal2 50232 8848 50232 8848 0 _0787_
rlabel metal2 49560 9016 49560 9016 0 _0788_
rlabel metal3 21952 11592 21952 11592 0 _0789_
rlabel metal2 19768 11424 19768 11424 0 _0790_
rlabel metal2 54936 10304 54936 10304 0 _0791_
rlabel metal2 55944 10248 55944 10248 0 _0792_
rlabel metal2 34888 25088 34888 25088 0 _0793_
rlabel metal2 49896 14784 49896 14784 0 _0794_
rlabel metal2 50792 13496 50792 13496 0 _0795_
rlabel metal2 45864 4648 45864 4648 0 _0796_
rlabel metal2 43736 5880 43736 5880 0 _0797_
rlabel metal3 47880 3304 47880 3304 0 _0798_
rlabel metal2 37800 5432 37800 5432 0 _0799_
rlabel metal3 39928 4312 39928 4312 0 _0800_
rlabel metal2 38192 3752 38192 3752 0 _0801_
rlabel metal3 40096 5768 40096 5768 0 _0802_
rlabel metal2 35560 6664 35560 6664 0 _0803_
rlabel metal3 34608 6664 34608 6664 0 _0804_
rlabel metal3 33880 6776 33880 6776 0 _0805_
rlabel metal2 38696 6328 38696 6328 0 _0806_
rlabel metal2 27944 10360 27944 10360 0 _0807_
rlabel metal2 17864 12208 17864 12208 0 _0808_
rlabel metal2 27944 8680 27944 8680 0 _0809_
rlabel metal2 28392 7728 28392 7728 0 _0810_
rlabel metal2 38808 6832 38808 6832 0 _0811_
rlabel metal2 37464 7672 37464 7672 0 _0812_
rlabel metal2 38920 8624 38920 8624 0 _0813_
rlabel metal2 23016 9408 23016 9408 0 _0814_
rlabel metal3 17248 10472 17248 10472 0 _0815_
rlabel metal3 24360 8232 24360 8232 0 _0816_
rlabel metal2 22232 8316 22232 8316 0 _0817_
rlabel metal2 22456 8736 22456 8736 0 _0818_
rlabel metal2 25928 8960 25928 8960 0 _0819_
rlabel metal3 21560 10584 21560 10584 0 _0820_
rlabel metal2 24360 10248 24360 10248 0 _0821_
rlabel metal2 19656 10416 19656 10416 0 _0822_
rlabel metal2 25368 11368 25368 11368 0 _0823_
rlabel metal2 38696 8512 38696 8512 0 _0824_
rlabel metal2 39928 9016 39928 9016 0 _0825_
rlabel metal2 39816 6384 39816 6384 0 _0826_
rlabel metal2 43624 7056 43624 7056 0 _0827_
rlabel metal2 45752 6776 45752 6776 0 _0828_
rlabel metal2 54936 14000 54936 14000 0 _0829_
rlabel metal2 53088 16184 53088 16184 0 _0830_
rlabel metal2 54824 15232 54824 15232 0 _0831_
rlabel metal3 43176 15176 43176 15176 0 _0832_
rlabel metal2 43456 15176 43456 15176 0 _0833_
rlabel metal3 47432 17808 47432 17808 0 _0834_
rlabel metal2 50344 21392 50344 21392 0 _0835_
rlabel metal2 54712 17192 54712 17192 0 _0836_
rlabel metal2 46536 16352 46536 16352 0 _0837_
rlabel metal2 23464 11312 23464 11312 0 _0838_
rlabel metal2 25256 10248 25256 10248 0 _0839_
rlabel metal2 25592 11480 25592 11480 0 _0840_
rlabel metal2 45752 18200 45752 18200 0 _0841_
rlabel metal2 53144 17192 53144 17192 0 _0842_
rlabel metal2 54376 16800 54376 16800 0 _0843_
rlabel metal2 55720 16800 55720 16800 0 _0844_
rlabel metal2 56952 16072 56952 16072 0 _0845_
rlabel metal2 55608 17528 55608 17528 0 _0846_
rlabel metal3 52976 18424 52976 18424 0 _0847_
rlabel metal3 50316 18424 50316 18424 0 _0848_
rlabel metal2 56056 18368 56056 18368 0 _0849_
rlabel metal2 56728 16576 56728 16576 0 _0850_
rlabel metal2 56112 15400 56112 15400 0 _0851_
rlabel metal2 54712 14000 54712 14000 0 _0852_
rlabel metal2 55440 12376 55440 12376 0 _0853_
rlabel metal2 54936 8512 54936 8512 0 _0854_
rlabel metal2 55496 8288 55496 8288 0 _0855_
rlabel metal2 54824 10528 54824 10528 0 _0856_
rlabel metal2 55160 9296 55160 9296 0 _0857_
rlabel metal2 22904 11200 22904 11200 0 _0858_
rlabel metal3 20664 11368 20664 11368 0 _0859_
rlabel metal3 13608 34776 13608 34776 0 _0860_
rlabel metal2 22568 11592 22568 11592 0 _0861_
rlabel metal2 18200 11648 18200 11648 0 _0862_
rlabel metal2 19768 17528 19768 17528 0 _0863_
rlabel metal2 27552 24696 27552 24696 0 _0864_
rlabel metal2 19880 19432 19880 19432 0 _0865_
rlabel metal2 56840 12152 56840 12152 0 _0866_
rlabel metal2 55496 9296 55496 9296 0 _0867_
rlabel metal3 56728 8792 56728 8792 0 _0868_
rlabel metal2 58072 11144 58072 11144 0 _0869_
rlabel metal2 52080 13048 52080 13048 0 _0870_
rlabel metal3 53928 14504 53928 14504 0 _0871_
rlabel metal2 55664 16072 55664 16072 0 _0872_
rlabel metal2 55160 14728 55160 14728 0 _0873_
rlabel metal2 56056 16240 56056 16240 0 _0874_
rlabel metal2 55048 19264 55048 19264 0 _0875_
rlabel metal2 55552 17864 55552 17864 0 _0876_
rlabel metal2 56280 21560 56280 21560 0 _0877_
rlabel metal2 52472 27776 52472 27776 0 _0878_
rlabel metal2 53928 27608 53928 27608 0 _0879_
rlabel metal3 42952 10248 42952 10248 0 _0880_
rlabel metal2 41160 5768 41160 5768 0 _0881_
rlabel metal2 38248 6776 38248 6776 0 _0882_
rlabel metal2 41496 17808 41496 17808 0 _0883_
rlabel metal3 43232 18424 43232 18424 0 _0884_
rlabel metal2 35392 6888 35392 6888 0 _0885_
rlabel metal2 36288 6888 36288 6888 0 _0886_
rlabel metal2 40264 12320 40264 12320 0 _0887_
rlabel metal3 32760 15848 32760 15848 0 _0888_
rlabel metal2 39928 13216 39928 13216 0 _0889_
rlabel metal2 40152 12712 40152 12712 0 _0890_
rlabel metal2 38920 7224 38920 7224 0 _0891_
rlabel metal2 40152 8064 40152 8064 0 _0892_
rlabel metal2 40936 11088 40936 11088 0 _0893_
rlabel metal2 35112 10080 35112 10080 0 _0894_
rlabel metal2 33656 9128 33656 9128 0 _0895_
rlabel metal2 23016 12432 23016 12432 0 _0896_
rlabel metal2 19096 18200 19096 18200 0 _0897_
rlabel metal2 31752 9128 31752 9128 0 _0898_
rlabel metal2 31192 9688 31192 9688 0 _0899_
rlabel metal2 34888 9968 34888 9968 0 _0900_
rlabel metal2 35784 11312 35784 11312 0 _0901_
rlabel metal2 36568 9016 36568 9016 0 _0902_
rlabel metal2 38136 8960 38136 8960 0 _0903_
rlabel metal2 37128 10528 37128 10528 0 _0904_
rlabel metal2 31920 12376 31920 12376 0 _0905_
rlabel metal2 28224 10472 28224 10472 0 _0906_
rlabel metal2 27608 15848 27608 15848 0 _0907_
rlabel metal2 32088 11480 32088 11480 0 _0908_
rlabel metal2 32816 12376 32816 12376 0 _0909_
rlabel metal2 33488 11480 33488 11480 0 _0910_
rlabel metal3 35168 10696 35168 10696 0 _0911_
rlabel metal2 41272 11648 41272 11648 0 _0912_
rlabel metal2 42952 17696 42952 17696 0 _0913_
rlabel metal2 41832 19152 41832 19152 0 _0914_
rlabel metal3 56056 26992 56056 26992 0 _0915_
rlabel metal2 56784 26936 56784 26936 0 _0916_
rlabel metal2 56056 17080 56056 17080 0 _0917_
rlabel metal2 57064 16352 57064 16352 0 _0918_
rlabel metal2 57176 24808 57176 24808 0 _0919_
rlabel metal2 54488 17696 54488 17696 0 _0920_
rlabel metal2 53536 26936 53536 26936 0 _0921_
rlabel metal2 45192 22736 45192 22736 0 _0922_
rlabel metal3 36400 23240 36400 23240 0 _0923_
rlabel metal2 45864 24864 45864 24864 0 _0924_
rlabel metal2 46032 24472 46032 24472 0 _0925_
rlabel metal2 46424 24640 46424 24640 0 _0926_
rlabel metal2 44856 18312 44856 18312 0 _0927_
rlabel metal2 45752 23688 45752 23688 0 _0928_
rlabel metal2 46984 25760 46984 25760 0 _0929_
rlabel metal2 54040 26040 54040 26040 0 _0930_
rlabel metal2 51576 24808 51576 24808 0 _0931_
rlabel metal2 48104 22456 48104 22456 0 _0932_
rlabel metal2 51576 23464 51576 23464 0 _0933_
rlabel metal2 49784 24080 49784 24080 0 _0934_
rlabel metal3 50260 23688 50260 23688 0 _0935_
rlabel metal3 51408 24808 51408 24808 0 _0936_
rlabel metal2 52584 24304 52584 24304 0 _0937_
rlabel metal2 51072 24696 51072 24696 0 _0938_
rlabel via2 53144 24696 53144 24696 0 _0939_
rlabel metal3 56224 26152 56224 26152 0 _0940_
rlabel metal2 57624 25032 57624 25032 0 _0941_
rlabel metal2 57960 16576 57960 16576 0 _0942_
rlabel metal2 57232 12264 57232 12264 0 _0943_
rlabel metal3 20608 15848 20608 15848 0 _0944_
rlabel metal2 18872 18480 18872 18480 0 _0945_
rlabel metal3 13048 29064 13048 29064 0 _0946_
rlabel metal2 20440 18704 20440 18704 0 _0947_
rlabel metal2 19488 20552 19488 20552 0 _0948_
rlabel metal2 56728 13048 56728 13048 0 _0949_
rlabel metal2 57624 13048 57624 13048 0 _0950_
rlabel metal2 57288 34552 57288 34552 0 _0951_
rlabel metal2 52584 28056 52584 28056 0 _0952_
rlabel metal2 57176 27496 57176 27496 0 _0953_
rlabel metal2 57288 29904 57288 29904 0 _0954_
rlabel metal2 56056 13496 56056 13496 0 _0955_
rlabel metal2 57624 14840 57624 14840 0 _0956_
rlabel metal2 54768 18088 54768 18088 0 _0957_
rlabel metal2 56168 25088 56168 25088 0 _0958_
rlabel metal3 55496 25480 55496 25480 0 _0959_
rlabel metal2 54040 30548 54040 30548 0 _0960_
rlabel metal3 53760 25256 53760 25256 0 _0961_
rlabel metal2 53704 26152 53704 26152 0 _0962_
rlabel metal3 53704 32536 53704 32536 0 _0963_
rlabel metal3 46648 25592 46648 25592 0 _0964_
rlabel metal2 44464 24696 44464 24696 0 _0965_
rlabel metal2 45528 25144 45528 25144 0 _0966_
rlabel metal2 44520 25760 44520 25760 0 _0967_
rlabel metal2 44856 31864 44856 31864 0 _0968_
rlabel metal2 39368 25872 39368 25872 0 _0969_
rlabel metal2 39760 26488 39760 26488 0 _0970_
rlabel metal2 39480 25536 39480 25536 0 _0971_
rlabel metal2 35000 25928 35000 25928 0 _0972_
rlabel metal3 41272 23128 41272 23128 0 _0973_
rlabel metal3 40768 26264 40768 26264 0 _0974_
rlabel metal2 41832 25592 41832 25592 0 _0975_
rlabel metal2 54040 32368 54040 32368 0 _0976_
rlabel metal2 54936 32928 54936 32928 0 _0977_
rlabel metal2 54264 34216 54264 34216 0 _0978_
rlabel metal2 52248 28168 52248 28168 0 _0979_
rlabel metal2 51184 33208 51184 33208 0 _0980_
rlabel metal2 42392 20832 42392 20832 0 _0981_
rlabel metal2 43848 19208 43848 19208 0 _0982_
rlabel metal2 46592 19992 46592 19992 0 _0983_
rlabel metal2 43960 20440 43960 20440 0 _0984_
rlabel metal2 46480 28504 46480 28504 0 _0985_
rlabel metal2 34664 17192 34664 17192 0 _0986_
rlabel metal3 40768 14504 40768 14504 0 _0987_
rlabel metal2 39648 12264 39648 12264 0 _0988_
rlabel metal2 40936 11872 40936 11872 0 _0989_
rlabel metal2 41160 13328 41160 13328 0 _0990_
rlabel metal2 34384 15288 34384 15288 0 _0991_
rlabel metal2 34552 15148 34552 15148 0 _0992_
rlabel metal2 35672 16072 35672 16072 0 _0993_
rlabel metal3 35168 14280 35168 14280 0 _0994_
rlabel metal2 36456 14112 36456 14112 0 _0995_
rlabel metal2 36456 11144 36456 11144 0 _0996_
rlabel metal2 36904 11088 36904 11088 0 _0997_
rlabel metal2 36344 12096 36344 12096 0 _0998_
rlabel metal2 22120 13440 22120 13440 0 _0999_
rlabel metal2 32424 13160 32424 13160 0 _1000_
rlabel metal2 32536 13272 32536 13272 0 _1001_
rlabel metal2 33880 12096 33880 12096 0 _1002_
rlabel metal2 33656 13328 33656 13328 0 _1003_
rlabel metal2 33992 12768 33992 12768 0 _1004_
rlabel metal2 29848 11480 29848 11480 0 _1005_
rlabel metal2 30296 11928 30296 11928 0 _1006_
rlabel metal2 31920 11368 31920 11368 0 _1007_
rlabel metal2 29624 10528 29624 10528 0 _1008_
rlabel metal2 31080 11760 31080 11760 0 _1009_
rlabel metal2 26376 11144 26376 11144 0 _1010_
rlabel metal2 27440 15400 27440 15400 0 _1011_
rlabel metal3 33040 12936 33040 12936 0 _1012_
rlabel metal2 37688 12544 37688 12544 0 _1013_
rlabel metal2 41384 13272 41384 13272 0 _1014_
rlabel metal2 42952 19936 42952 19936 0 _1015_
rlabel metal2 43792 21672 43792 21672 0 _1016_
rlabel metal2 45304 29008 45304 29008 0 _1017_
rlabel metal2 44968 29064 44968 29064 0 _1018_
rlabel metal2 45752 29848 45752 29848 0 _1019_
rlabel metal3 50904 33208 50904 33208 0 _1020_
rlabel metal3 53984 34104 53984 34104 0 _1021_
rlabel metal2 56056 31836 56056 31836 0 _1022_
rlabel metal2 55832 32760 55832 32760 0 _1023_
rlabel metal2 56616 34496 56616 34496 0 _1024_
rlabel metal2 20104 34104 20104 34104 0 _1025_
rlabel metal3 14616 34104 14616 34104 0 _1026_
rlabel metal2 21224 33712 21224 33712 0 _1027_
rlabel metal2 20328 34832 20328 34832 0 _1028_
rlabel metal2 50792 31528 50792 31528 0 _1029_
rlabel metal2 57624 34104 57624 34104 0 _1030_
rlabel metal2 56112 32760 56112 32760 0 _1031_
rlabel metal2 52808 35616 52808 35616 0 _1032_
rlabel metal2 54712 34664 54712 34664 0 _1033_
rlabel metal3 55888 35672 55888 35672 0 _1034_
rlabel metal2 52808 36176 52808 36176 0 _1035_
rlabel metal2 50792 33824 50792 33824 0 _1036_
rlabel metal2 50120 33824 50120 33824 0 _1037_
rlabel metal2 50568 34608 50568 34608 0 _1038_
rlabel metal2 53256 32816 53256 32816 0 _1039_
rlabel metal2 53704 33320 53704 33320 0 _1040_
rlabel metal2 48888 34048 48888 34048 0 _1041_
rlabel metal2 38808 32816 38808 32816 0 _1042_
rlabel metal3 44576 32760 44576 32760 0 _1043_
rlabel metal2 43960 25592 43960 25592 0 _1044_
rlabel metal2 40152 31472 40152 31472 0 _1045_
rlabel metal3 13384 26936 13384 26936 0 _1046_
rlabel metal3 25144 26264 25144 26264 0 _1047_
rlabel metal3 35392 26488 35392 26488 0 _1048_
rlabel metal3 37352 25256 37352 25256 0 _1049_
rlabel metal3 37464 25368 37464 25368 0 _1050_
rlabel metal2 36400 26040 36400 26040 0 _1051_
rlabel metal3 39704 31640 39704 31640 0 _1052_
rlabel metal3 42840 31752 42840 31752 0 _1053_
rlabel metal2 46032 33208 46032 33208 0 _1054_
rlabel metal3 45136 33320 45136 33320 0 _1055_
rlabel metal2 43624 29792 43624 29792 0 _1056_
rlabel metal2 42952 29792 42952 29792 0 _1057_
rlabel metal2 43736 29400 43736 29400 0 _1058_
rlabel metal2 41720 32704 41720 32704 0 _1059_
rlabel metal2 40824 26684 40824 26684 0 _1060_
rlabel metal2 39984 26152 39984 26152 0 _1061_
rlabel metal2 40264 31640 40264 31640 0 _1062_
rlabel metal2 41272 20832 41272 20832 0 _1063_
rlabel metal2 44184 21112 44184 21112 0 _1064_
rlabel metal2 41496 20944 41496 20944 0 _1065_
rlabel metal2 39480 20720 39480 20720 0 _1066_
rlabel metal2 40376 14000 40376 14000 0 _1067_
rlabel metal2 41720 13832 41720 13832 0 _1068_
rlabel metal2 40824 15568 40824 15568 0 _1069_
rlabel metal3 35168 17640 35168 17640 0 _1070_
rlabel metal2 24248 17416 24248 17416 0 _1071_
rlabel metal2 35560 17864 35560 17864 0 _1072_
rlabel metal2 34496 20104 34496 20104 0 _1073_
rlabel metal2 36960 12264 36960 12264 0 _1074_
rlabel metal2 37352 13048 37352 13048 0 _1075_
rlabel metal2 34664 19152 34664 19152 0 _1076_
rlabel metal3 30352 15848 30352 15848 0 _1077_
rlabel metal2 25984 11256 25984 11256 0 _1078_
rlabel metal2 26544 15288 26544 15288 0 _1079_
rlabel metal2 26824 14504 26824 14504 0 _1080_
rlabel metal2 29456 12936 29456 12936 0 _1081_
rlabel metal2 23240 11312 23240 11312 0 _1082_
rlabel metal2 30520 13104 30520 13104 0 _1083_
rlabel metal3 24416 13944 24416 13944 0 _1084_
rlabel metal2 28616 14000 28616 14000 0 _1085_
rlabel metal3 28672 15288 28672 15288 0 _1086_
rlabel metal3 30072 16072 30072 16072 0 _1087_
rlabel metal2 31080 18200 31080 18200 0 _1088_
rlabel metal2 32536 13832 32536 13832 0 _1089_
rlabel metal2 34496 13608 34496 13608 0 _1090_
rlabel metal2 34440 18032 34440 18032 0 _1091_
rlabel metal2 33656 17360 33656 17360 0 _1092_
rlabel metal2 32200 18536 32200 18536 0 _1093_
rlabel metal3 32760 18424 32760 18424 0 _1094_
rlabel metal2 31528 18928 31528 18928 0 _1095_
rlabel metal3 34272 19992 34272 19992 0 _1096_
rlabel metal2 36344 20888 36344 20888 0 _1097_
rlabel metal2 37352 20328 37352 20328 0 _1098_
rlabel metal2 36568 29008 36568 29008 0 _1099_
rlabel metal2 22232 27328 22232 27328 0 _1100_
rlabel metal2 35672 29232 35672 29232 0 _1101_
rlabel metal3 40040 30128 40040 30128 0 _1102_
rlabel metal2 41272 31864 41272 31864 0 _1103_
rlabel metal2 47544 33712 47544 33712 0 _1104_
rlabel metal2 50176 33320 50176 33320 0 _1105_
rlabel metal2 52920 35784 52920 35784 0 _1106_
rlabel metal2 51688 36064 51688 36064 0 _1107_
rlabel metal2 21336 34664 21336 34664 0 _1108_
rlabel metal3 10024 34160 10024 34160 0 _1109_
rlabel metal3 50736 34776 50736 34776 0 _1110_
rlabel metal2 51912 34496 51912 34496 0 _1111_
rlabel metal2 21672 35280 21672 35280 0 _1112_
rlabel metal2 22624 16632 22624 16632 0 _1113_
rlabel metal2 53368 35112 53368 35112 0 _1114_
rlabel metal2 52136 36288 52136 36288 0 _1115_
rlabel metal3 48272 34104 48272 34104 0 _1116_
rlabel metal2 49280 34216 49280 34216 0 _1117_
rlabel metal2 49784 33712 49784 33712 0 _1118_
rlabel metal2 49448 33936 49448 33936 0 _1119_
rlabel metal3 40936 32536 40936 32536 0 _1120_
rlabel metal2 41160 32480 41160 32480 0 _1121_
rlabel metal2 40936 32480 40936 32480 0 _1122_
rlabel metal2 41048 32424 41048 32424 0 _1123_
rlabel metal2 41608 32928 41608 32928 0 _1124_
rlabel metal2 44688 31752 44688 31752 0 _1125_
rlabel metal2 43848 33600 43848 33600 0 _1126_
rlabel metal2 36008 31696 36008 31696 0 _1127_
rlabel metal3 37520 32648 37520 32648 0 _1128_
rlabel metal2 38808 32200 38808 32200 0 _1129_
rlabel metal2 34216 24500 34216 24500 0 _1130_
rlabel metal2 33992 26152 33992 26152 0 _1131_
rlabel metal2 33880 28896 33880 28896 0 _1132_
rlabel metal2 26432 19208 26432 19208 0 _1133_
rlabel metal3 33544 29624 33544 29624 0 _1134_
rlabel metal2 33656 29288 33656 29288 0 _1135_
rlabel metal3 22680 22344 22680 22344 0 _1136_
rlabel metal2 21392 26824 21392 26824 0 _1137_
rlabel metal2 33432 28952 33432 28952 0 _1138_
rlabel metal3 34440 31752 34440 31752 0 _1139_
rlabel metal2 39480 32200 39480 32200 0 _1140_
rlabel metal2 38248 33712 38248 33712 0 _1141_
rlabel metal3 36344 29288 36344 29288 0 _1142_
rlabel metal2 35560 29848 35560 29848 0 _1143_
rlabel metal3 34832 31080 34832 31080 0 _1144_
rlabel metal3 36568 25704 36568 25704 0 _1145_
rlabel metal2 36344 26824 36344 26824 0 _1146_
rlabel metal2 36064 30856 36064 30856 0 _1147_
rlabel metal3 37296 20776 37296 20776 0 _1148_
rlabel metal2 37240 21560 37240 21560 0 _1149_
rlabel metal2 30520 21112 30520 21112 0 _1150_
rlabel metal2 33096 19600 33096 19600 0 _1151_
rlabel metal2 32872 19432 32872 19432 0 _1152_
rlabel metal2 33880 19264 33880 19264 0 _1153_
rlabel metal2 29960 19656 29960 19656 0 _1154_
rlabel metal2 25816 18312 25816 18312 0 _1155_
rlabel metal2 33768 18424 33768 18424 0 _1156_
rlabel metal3 31360 19096 31360 19096 0 _1157_
rlabel metal2 30072 16184 30072 16184 0 _1158_
rlabel metal2 31528 17640 31528 17640 0 _1159_
rlabel metal2 30632 18256 30632 18256 0 _1160_
rlabel metal2 28280 14896 28280 14896 0 _1161_
rlabel metal2 28280 15848 28280 15848 0 _1162_
rlabel metal3 24304 14504 24304 14504 0 _1163_
rlabel metal3 23968 12152 23968 12152 0 _1164_
rlabel metal3 23856 13720 23856 13720 0 _1165_
rlabel metal3 24976 14280 24976 14280 0 _1166_
rlabel metal2 26040 15624 26040 15624 0 _1167_
rlabel metal2 27608 16128 27608 16128 0 _1168_
rlabel metal2 27384 17248 27384 17248 0 _1169_
rlabel metal2 29232 12936 29232 12936 0 _1170_
rlabel metal3 30128 12712 30128 12712 0 _1171_
rlabel metal2 30688 17528 30688 17528 0 _1172_
rlabel metal2 32312 16408 32312 16408 0 _1173_
rlabel metal2 29624 17528 29624 17528 0 _1174_
rlabel metal2 30128 17752 30128 17752 0 _1175_
rlabel metal3 28560 17640 28560 17640 0 _1176_
rlabel metal2 28392 18368 28392 18368 0 _1177_
rlabel metal3 28784 19208 28784 19208 0 _1178_
rlabel metal3 28560 19992 28560 19992 0 _1179_
rlabel metal3 28392 25704 28392 25704 0 _1180_
rlabel metal2 12880 28504 12880 28504 0 _1181_
rlabel metal2 23016 28672 23016 28672 0 _1182_
rlabel metal2 14504 28616 14504 28616 0 _1183_
rlabel metal2 25256 26544 25256 26544 0 _1184_
rlabel metal2 23352 28840 23352 28840 0 _1185_
rlabel metal2 25928 28840 25928 28840 0 _1186_
rlabel metal2 31864 31024 31864 31024 0 _1187_
rlabel metal2 39144 33712 39144 33712 0 _1188_
rlabel metal3 39872 34104 39872 34104 0 _1189_
rlabel metal2 36904 34048 36904 34048 0 _1190_
rlabel metal2 24472 35336 24472 35336 0 _1191_
rlabel metal2 22568 34944 22568 34944 0 _1192_
rlabel metal2 21784 34608 21784 34608 0 _1193_
rlabel metal2 21952 35448 21952 35448 0 _1194_
rlabel metal2 25928 35168 25928 35168 0 _1195_
rlabel metal2 24248 34496 24248 34496 0 _1196_
rlabel metal2 26712 20048 26712 20048 0 _1197_
rlabel metal2 33768 34944 33768 34944 0 _1198_
rlabel metal2 36568 34496 36568 34496 0 _1199_
rlabel metal2 32984 34496 32984 34496 0 _1200_
rlabel metal2 39032 34048 39032 34048 0 _1201_
rlabel metal3 36512 33208 36512 33208 0 _1202_
rlabel metal2 35560 33600 35560 33600 0 _1203_
rlabel metal2 35448 33488 35448 33488 0 _1204_
rlabel metal2 23968 24920 23968 24920 0 _1205_
rlabel metal3 30016 30184 30016 30184 0 _1206_
rlabel metal2 31752 30968 31752 30968 0 _1207_
rlabel metal2 32704 30856 32704 30856 0 _1208_
rlabel metal2 33208 31416 33208 31416 0 _1209_
rlabel metal2 32312 31976 32312 31976 0 _1210_
rlabel metal3 38808 32536 38808 32536 0 _1211_
rlabel metal2 32648 33152 32648 33152 0 _1212_
rlabel metal3 25200 28392 25200 28392 0 _1213_
rlabel metal2 25480 28504 25480 28504 0 _1214_
rlabel metal3 24416 29960 24416 29960 0 _1215_
rlabel metal2 25816 29008 25816 29008 0 _1216_
rlabel metal2 24584 30352 24584 30352 0 _1217_
rlabel metal2 30464 20216 30464 20216 0 _1218_
rlabel metal2 28056 21784 28056 21784 0 _1219_
rlabel metal2 23800 21056 23800 21056 0 _1220_
rlabel metal2 29904 18648 29904 18648 0 _1221_
rlabel metal2 22904 19264 22904 19264 0 _1222_
rlabel metal2 30744 18144 30744 18144 0 _1223_
rlabel metal2 20664 17976 20664 17976 0 _1224_
rlabel metal2 28392 16576 28392 16576 0 _1225_
rlabel metal2 21784 16744 21784 16744 0 _1226_
rlabel metal2 27272 15624 27272 15624 0 _1227_
rlabel metal2 21448 15344 21448 15344 0 _1228_
rlabel metal2 23240 13944 23240 13944 0 _1229_
rlabel metal3 23072 13832 23072 13832 0 _1230_
rlabel metal2 21560 15148 21560 15148 0 _1231_
rlabel metal3 22008 17080 22008 17080 0 _1232_
rlabel metal2 25928 14672 25928 14672 0 _1233_
rlabel metal2 25368 16296 25368 16296 0 _1234_
rlabel metal3 25144 16072 25144 16072 0 _1235_
rlabel metal3 25256 16856 25256 16856 0 _1236_
rlabel metal2 25592 15932 25592 15932 0 _1237_
rlabel metal2 23464 16856 23464 16856 0 _1238_
rlabel metal2 22680 16912 22680 16912 0 _1239_
rlabel via2 21336 17640 21336 17640 0 _1240_
rlabel metal2 22792 18928 22792 18928 0 _1241_
rlabel metal3 20328 21784 20328 21784 0 _1242_
rlabel metal2 20272 30072 20272 30072 0 _1243_
rlabel metal3 21000 22344 21000 22344 0 _1244_
rlabel metal2 18592 30296 18592 30296 0 _1245_
rlabel metal2 19320 29736 19320 29736 0 _1246_
rlabel metal3 21784 29400 21784 29400 0 _1247_
rlabel metal2 26600 30856 26600 30856 0 _1248_
rlabel metal2 33432 32032 33432 32032 0 _1249_
rlabel metal2 26712 31080 26712 31080 0 _1250_
rlabel metal2 33152 30184 33152 30184 0 _1251_
rlabel metal2 34776 31416 34776 31416 0 _1252_
rlabel metal2 27720 31808 27720 31808 0 _1253_
rlabel metal2 26152 31080 26152 31080 0 _1254_
rlabel metal3 28728 32536 28728 32536 0 _1255_
rlabel metal2 34048 33432 34048 33432 0 _1256_
rlabel metal3 33208 33992 33208 33992 0 _1257_
rlabel metal2 26040 34048 26040 34048 0 _1258_
rlabel metal2 24024 33992 24024 33992 0 _1259_
rlabel metal2 12600 33544 12600 33544 0 _1260_
rlabel metal2 14952 30128 14952 30128 0 _1261_
rlabel metal2 34664 33264 34664 33264 0 _1262_
rlabel metal3 29848 33936 29848 33936 0 _1263_
rlabel metal2 22456 33600 22456 33600 0 _1264_
rlabel metal2 32704 32536 32704 32536 0 _1265_
rlabel metal3 32032 32536 32032 32536 0 _1266_
rlabel metal3 26096 32648 26096 32648 0 _1267_
rlabel metal2 23464 20496 23464 20496 0 _1268_
rlabel metal2 23352 20664 23352 20664 0 _1269_
rlabel metal2 21952 15512 21952 15512 0 _1270_
rlabel metal2 20888 18032 20888 18032 0 _1271_
rlabel metal2 21448 19600 21448 19600 0 _1272_
rlabel metal2 21896 21504 21896 21504 0 _1273_
rlabel metal2 22680 20328 22680 20328 0 _1274_
rlabel metal3 23688 15288 23688 15288 0 _1275_
rlabel metal2 25984 18424 25984 18424 0 _1276_
rlabel metal2 24808 18480 24808 18480 0 _1277_
rlabel metal2 24584 17136 24584 17136 0 _1278_
rlabel metal2 26320 18424 26320 18424 0 _1279_
rlabel metal2 25256 17696 25256 17696 0 _1280_
rlabel metal2 23688 15680 23688 15680 0 _1281_
rlabel metal3 21840 14280 21840 14280 0 _1282_
rlabel metal2 20608 16072 20608 16072 0 _1283_
rlabel metal2 21784 16128 21784 16128 0 _1284_
rlabel metal2 24360 19992 24360 19992 0 _1285_
rlabel metal2 25368 12712 25368 12712 0 _1286_
rlabel metal2 24920 13216 24920 13216 0 _1287_
rlabel metal2 22344 18928 22344 18928 0 _1288_
rlabel metal2 21784 21952 21784 21952 0 _1289_
rlabel metal2 19768 28896 19768 28896 0 _1290_
rlabel metal2 19152 31192 19152 31192 0 _1291_
rlabel metal2 19712 30408 19712 30408 0 _1292_
rlabel metal3 20552 31192 20552 31192 0 _1293_
rlabel metal2 26376 32200 26376 32200 0 _1294_
rlabel metal2 25928 32144 25928 32144 0 _1295_
rlabel metal2 21560 31808 21560 31808 0 _1296_
rlabel metal2 21224 28672 21224 28672 0 _1297_
rlabel metal2 21616 29624 21616 29624 0 _1298_
rlabel metal2 32088 29848 32088 29848 0 _1299_
rlabel metal2 23688 29792 23688 29792 0 _1300_
rlabel metal2 24080 30408 24080 30408 0 _1301_
rlabel metal2 23352 30408 23352 30408 0 _1302_
rlabel metal2 23016 30968 23016 30968 0 _1303_
rlabel metal2 24024 31024 24024 31024 0 _1304_
rlabel metal2 23912 31416 23912 31416 0 _1305_
rlabel metal2 23128 32088 23128 32088 0 _1306_
rlabel metal2 23240 33040 23240 33040 0 _1307_
rlabel metal2 24920 33656 24920 33656 0 _1308_
rlabel metal2 24136 33656 24136 33656 0 _1309_
rlabel metal2 7616 33096 7616 33096 0 _1310_
rlabel metal2 13888 28616 13888 28616 0 _1311_
rlabel metal3 7112 15288 7112 15288 0 _1312_
rlabel metal2 7224 16352 7224 16352 0 _1313_
rlabel metal3 4144 14504 4144 14504 0 _1314_
rlabel metal3 6272 14616 6272 14616 0 _1315_
rlabel metal2 6328 16184 6328 16184 0 _1316_
rlabel metal2 5880 14392 5880 14392 0 _1317_
rlabel metal2 9016 15512 9016 15512 0 _1318_
rlabel metal2 8120 13272 8120 13272 0 _1319_
rlabel metal2 8736 12824 8736 12824 0 _1320_
rlabel metal2 6832 12152 6832 12152 0 _1321_
rlabel metal2 7560 12208 7560 12208 0 _1322_
rlabel metal2 6216 8736 6216 8736 0 _1323_
rlabel metal2 2856 7784 2856 7784 0 _1324_
rlabel metal2 2296 9576 2296 9576 0 _1325_
rlabel metal3 7056 7336 7056 7336 0 _1326_
rlabel metal3 6608 7448 6608 7448 0 _1327_
rlabel metal2 4648 6664 4648 6664 0 _1328_
rlabel metal2 4760 4816 4760 4816 0 _1329_
rlabel metal2 9128 6160 9128 6160 0 _1330_
rlabel metal2 5096 5488 5096 5488 0 _1331_
rlabel metal2 4984 5936 4984 5936 0 _1332_
rlabel metal2 6664 5208 6664 5208 0 _1333_
rlabel metal2 8120 4648 8120 4648 0 _1334_
rlabel metal2 13552 11256 13552 11256 0 _1335_
rlabel metal2 9912 4816 9912 4816 0 _1336_
rlabel metal2 10248 4592 10248 4592 0 _1337_
rlabel metal2 12152 4144 12152 4144 0 _1338_
rlabel metal3 23296 2408 23296 2408 0 _1339_
rlabel metal3 11704 4312 11704 4312 0 _1340_
rlabel metal2 13272 4200 13272 4200 0 _1341_
rlabel metal2 13720 4592 13720 4592 0 _1342_
rlabel metal2 12712 4592 12712 4592 0 _1343_
rlabel metal2 15400 7784 15400 7784 0 _1344_
rlabel metal2 14056 5824 14056 5824 0 _1345_
rlabel metal3 12992 5880 12992 5880 0 _1346_
rlabel metal3 15624 8064 15624 8064 0 _1347_
rlabel metal2 13496 6776 13496 6776 0 _1348_
rlabel metal3 11648 9912 11648 9912 0 _1349_
rlabel metal3 13440 8008 13440 8008 0 _1350_
rlabel metal3 14000 8120 14000 8120 0 _1351_
rlabel metal2 15176 9296 15176 9296 0 _1352_
rlabel metal2 15904 9688 15904 9688 0 _1353_
rlabel metal2 9016 16408 9016 16408 0 _1354_
rlabel metal2 7000 16856 7000 16856 0 _1355_
rlabel metal3 47152 20664 47152 20664 0 _1356_
rlabel metal3 22232 9408 22232 9408 0 a\[0\]\[0\]
rlabel metal2 19656 9576 19656 9576 0 a\[0\]\[1\]
rlabel metal3 21056 16184 21056 16184 0 a\[0\]\[2\]
rlabel metal2 22456 12488 22456 12488 0 a\[0\]\[3\]
rlabel metal2 18760 11256 18760 11256 0 a\[0\]\[4\]
rlabel metal2 21448 13664 21448 13664 0 a\[0\]\[5\]
rlabel metal2 23352 16912 23352 16912 0 a\[0\]\[6\]
rlabel metal2 25368 15680 25368 15680 0 a\[0\]\[7\]
rlabel metal2 4648 18480 4648 18480 0 a\[1\]\[0\]
rlabel metal3 8176 24584 8176 24584 0 a\[1\]\[1\]
rlabel metal2 8568 27020 8568 27020 0 a\[1\]\[2\]
rlabel metal2 8120 22904 8120 22904 0 a\[1\]\[3\]
rlabel metal2 7672 28896 7672 28896 0 a\[1\]\[4\]
rlabel metal2 8344 31780 8344 31780 0 a\[1\]\[5\]
rlabel metal2 6664 30856 6664 30856 0 a\[1\]\[6\]
rlabel metal3 11872 31528 11872 31528 0 a\[1\]\[7\]
rlabel metal3 40768 16968 40768 16968 0 b\[0\]\[0\]
rlabel metal3 42672 15512 42672 15512 0 b\[0\]\[1\]
rlabel metal2 43176 17416 43176 17416 0 b\[0\]\[2\]
rlabel metal2 46872 18312 46872 18312 0 b\[0\]\[3\]
rlabel metal2 46536 24080 46536 24080 0 b\[0\]\[4\]
rlabel metal2 50288 25256 50288 25256 0 b\[0\]\[5\]
rlabel metal2 14280 27664 14280 27664 0 b\[0\]\[6\]
rlabel metal2 13608 29288 13608 29288 0 b\[0\]\[7\]
rlabel metal3 4984 20888 4984 20888 0 b\[1\]\[0\]
rlabel metal3 6552 25592 6552 25592 0 b\[1\]\[1\]
rlabel metal3 6104 26376 6104 26376 0 b\[1\]\[2\]
rlabel metal2 4648 22792 4648 22792 0 b\[1\]\[3\]
rlabel metal2 4760 29064 4760 29064 0 b\[1\]\[4\]
rlabel metal2 4648 33376 4648 33376 0 b\[1\]\[5\]
rlabel metal3 6888 31864 6888 31864 0 b\[1\]\[6\]
rlabel metal3 10416 32424 10416 32424 0 b\[1\]\[7\]
rlabel metal3 8288 27832 8288 27832 0 bflip
rlabel metal2 47880 21112 47880 21112 0 c\[0\]\[0\]
rlabel metal3 21000 21392 21000 21392 0 c\[0\]\[1\]
rlabel metal2 19096 18984 19096 18984 0 c\[0\]\[2\]
rlabel metal2 19544 20944 19544 20944 0 c\[0\]\[3\]
rlabel metal2 20272 23016 20272 23016 0 c\[0\]\[4\]
rlabel metal2 22456 21560 22456 21560 0 c\[0\]\[5\]
rlabel metal2 24584 26152 24584 26152 0 c\[0\]\[6\]
rlabel metal2 15512 24808 15512 24808 0 c\[0\]\[7\]
rlabel metal2 56616 35560 56616 35560 0 clk
rlabel metal2 26488 23184 26488 23184 0 clknet_0_clk
rlabel metal3 2464 16856 2464 16856 0 clknet_1_0__leaf_clk
rlabel metal2 4200 36064 4200 36064 0 clknet_1_1__leaf_clk
rlabel metal3 11144 15176 11144 15176 0 delta_t\[0\]
rlabel metal3 6048 15400 6048 15400 0 delta_t\[1\]
rlabel metal2 5768 12432 5768 12432 0 delta_t\[2\]
rlabel metal2 5656 10472 5656 10472 0 delta_t\[3\]
rlabel metal2 4648 9800 4648 9800 0 delta_t\[4\]
rlabel metal2 15848 5488 15848 5488 0 delta_t\[5\]
rlabel metal2 18648 8456 18648 8456 0 delta_t\[6\]
rlabel metal2 12544 6664 12544 6664 0 delta_t\[7\]
rlabel metal2 15680 8904 15680 8904 0 delta_t\[8\]
rlabel metal3 14336 9016 14336 9016 0 delta_t\[9\]
rlabel metal2 2968 4984 2968 4984 0 net1
rlabel metal2 2800 23688 2800 23688 0 net10
rlabel metal2 42392 5040 42392 5040 0 net100
rlabel metal3 16800 16968 16800 16968 0 net11
rlabel metal2 4536 28112 4536 28112 0 net12
rlabel metal2 3528 33992 3528 33992 0 net13
rlabel metal2 5712 29960 5712 29960 0 net14
rlabel metal2 3752 29400 3752 29400 0 net15
rlabel metal3 16800 21672 16800 21672 0 net16
rlabel metal3 1792 16744 1792 16744 0 net17
rlabel metal2 2072 13832 2072 13832 0 net18
rlabel metal2 8120 28728 8120 28728 0 net19
rlabel metal2 7672 18032 7672 18032 0 net2
rlabel metal2 10360 29232 10360 29232 0 net20
rlabel metal2 9856 28392 9856 28392 0 net21
rlabel metal2 5152 27944 5152 27944 0 net22
rlabel metal2 2072 26040 2072 26040 0 net23
rlabel metal2 30296 3136 30296 3136 0 net24
rlabel metal3 15400 8736 15400 8736 0 net25
rlabel metal2 29512 4256 29512 4256 0 net26
rlabel metal2 15848 3808 15848 3808 0 net27
rlabel metal2 17752 4648 17752 4648 0 net28
rlabel metal2 55048 36624 55048 36624 0 net29
rlabel metal3 28728 2744 28728 2744 0 net3
rlabel metal2 53592 36120 53592 36120 0 net30
rlabel metal2 46088 35280 46088 35280 0 net31
rlabel metal3 43512 36288 43512 36288 0 net32
rlabel metal2 47656 35560 47656 35560 0 net33
rlabel metal2 47824 36232 47824 36232 0 net34
rlabel metal2 42616 35560 42616 35560 0 net35
rlabel metal2 36456 35728 36456 35728 0 net36
rlabel metal3 21784 7952 21784 7952 0 net37
rlabel metal2 18200 35280 18200 35280 0 net38
rlabel metal3 16464 35560 16464 35560 0 net39
rlabel metal3 35616 2632 35616 2632 0 net4
rlabel metal2 14392 36512 14392 36512 0 net40
rlabel metal2 11816 35336 11816 35336 0 net41
rlabel metal2 8792 36624 8792 36624 0 net42
rlabel metal2 7112 35616 7112 35616 0 net43
rlabel metal3 5040 36568 5040 36568 0 net44
rlabel metal2 5656 35168 5656 35168 0 net45
rlabel metal2 37240 36512 37240 36512 0 net46
rlabel metal2 35784 35728 35784 35728 0 net47
rlabel metal2 32536 35616 32536 35616 0 net48
rlabel metal2 31304 35728 31304 35728 0 net49
rlabel metal2 16072 4088 16072 4088 0 net5
rlabel metal3 28392 35560 28392 35560 0 net50
rlabel metal2 21168 35560 21168 35560 0 net51
rlabel metal2 15624 34160 15624 34160 0 net52
rlabel metal2 19040 33432 19040 33432 0 net53
rlabel metal2 1848 10976 1848 10976 0 net54
rlabel metal2 9800 7448 9800 7448 0 net55
rlabel metal2 1904 15288 1904 15288 0 net56
rlabel metal2 16912 9800 16912 9800 0 net57
rlabel metal2 17752 14840 17752 14840 0 net58
rlabel metal2 16408 13160 16408 13160 0 net59
rlabel metal2 5488 28392 5488 28392 0 net6
rlabel metal2 5544 12488 5544 12488 0 net60
rlabel metal2 1848 21958 1848 21958 0 net61
rlabel metal2 2072 25200 2072 25200 0 net62
rlabel metal2 2296 20720 2296 20720 0 net63
rlabel metal2 5320 28224 5320 28224 0 net64
rlabel metal2 4648 31752 4648 31752 0 net65
rlabel metal2 4984 31360 4984 31360 0 net66
rlabel metal2 10248 29624 10248 29624 0 net67
rlabel metal3 10696 30184 10696 30184 0 net68
rlabel metal3 16632 20664 16632 20664 0 net69
rlabel metal2 2072 19264 2072 19264 0 net7
rlabel metal3 12712 27832 12712 27832 0 net70
rlabel metal2 2352 22120 2352 22120 0 net71
rlabel metal4 3752 17528 3752 17528 0 net72
rlabel metal2 37576 17808 37576 17808 0 net73
rlabel metal2 19656 21560 19656 21560 0 net74
rlabel metal2 20328 21896 20328 21896 0 net75
rlabel metal2 51800 31192 51800 31192 0 net76
rlabel metal2 22176 10472 22176 10472 0 net77
rlabel metal2 33096 5152 33096 5152 0 net78
rlabel metal2 32144 6552 32144 6552 0 net79
rlabel metal2 3304 24024 3304 24024 0 net8
rlabel metal2 22680 4816 22680 4816 0 net80
rlabel metal2 47936 32648 47936 32648 0 net81
rlabel metal2 54376 30856 54376 30856 0 net82
rlabel metal3 20384 7336 20384 7336 0 net83
rlabel metal2 45080 4200 45080 4200 0 net84
rlabel metal2 39032 6440 39032 6440 0 net85
rlabel metal2 41160 5040 41160 5040 0 net86
rlabel metal2 40376 5040 40376 5040 0 net87
rlabel metal2 26824 6384 26824 6384 0 net88
rlabel metal2 27608 5768 27608 5768 0 net89
rlabel metal2 2184 22792 2184 22792 0 net9
rlabel metal2 42392 17752 42392 17752 0 net90
rlabel metal3 43624 18648 43624 18648 0 net91
rlabel metal2 41944 5768 41944 5768 0 net92
rlabel metal3 35112 8344 35112 8344 0 net93
rlabel metal2 23072 3528 23072 3528 0 net94
rlabel metal2 39704 5320 39704 5320 0 net95
rlabel metal2 38136 6272 38136 6272 0 net96
rlabel metal3 41384 5880 41384 5880 0 net97
rlabel metal2 25256 6440 25256 6440 0 net98
rlabel metal2 41216 8456 41216 8456 0 net99
rlabel metal2 6776 15680 6776 15680 0 t_reg\[0\]
rlabel metal2 5768 16128 5768 16128 0 t_reg\[1\]
rlabel metal3 6440 12376 6440 12376 0 t_reg\[2\]
rlabel metal2 4648 8680 4648 8680 0 t_reg\[3\]
rlabel metal2 7224 4256 7224 4256 0 t_reg\[4\]
rlabel metal2 9352 3752 9352 3752 0 t_reg\[5\]
rlabel metal2 27888 3640 27888 3640 0 t_reg\[6\]
rlabel metal2 16968 4088 16968 4088 0 t_reg\[7\]
rlabel metal2 4816 6776 4816 6776 0 t_reg\[8\]
rlabel metal2 20440 9296 20440 9296 0 t_reg\[9\]
rlabel metal2 2968 3192 2968 3192 0 wb_clk_i
rlabel metal2 7896 2184 7896 2184 0 wb_rst_i
rlabel metal2 56952 1190 56952 1190 0 wbs_ack_o
rlabel metal2 47432 4256 47432 4256 0 wbs_adr_i[2]
rlabel metal2 52136 3416 52136 3416 0 wbs_adr_i[3]
rlabel metal2 17528 2086 17528 2086 0 wbs_cyc_i
rlabel metal2 3528 36064 3528 36064 0 wbs_dat_i[0]
rlabel metal3 854 19320 854 19320 0 wbs_dat_i[16]
rlabel metal2 1736 17920 1736 17920 0 wbs_dat_i[17]
rlabel metal2 2632 17360 2632 17360 0 wbs_dat_i[18]
rlabel metal2 1736 16408 1736 16408 0 wbs_dat_i[19]
rlabel metal2 11592 33936 11592 33936 0 wbs_dat_i[1]
rlabel metal3 910 14840 910 14840 0 wbs_dat_i[20]
rlabel metal2 2352 14392 2352 14392 0 wbs_dat_i[21]
rlabel metal2 1736 11648 1736 11648 0 wbs_dat_i[22]
rlabel metal3 854 11480 854 11480 0 wbs_dat_i[23]
rlabel metal3 8400 35504 8400 35504 0 wbs_dat_i[2]
rlabel metal2 1848 34384 1848 34384 0 wbs_dat_i[3]
rlabel metal2 1680 34104 1680 34104 0 wbs_dat_i[4]
rlabel metal2 6216 32648 6216 32648 0 wbs_dat_i[5]
rlabel metal2 5096 29848 5096 29848 0 wbs_dat_i[6]
rlabel metal3 2744 29960 2744 29960 0 wbs_dat_i[7]
rlabel metal2 1736 29176 1736 29176 0 wbs_dat_i[8]
rlabel metal2 2520 26600 2520 26600 0 wbs_dat_i[9]
rlabel metal3 32872 3528 32872 3528 0 wbs_sel_i[0]
rlabel metal2 32536 2184 32536 2184 0 wbs_sel_i[1]
rlabel metal2 37408 2520 37408 2520 0 wbs_sel_i[2]
rlabel metal2 10584 4032 10584 4032 0 wbs_stb_i
rlabel metal2 22456 1302 22456 1302 0 wbs_we_i
rlabel metal2 19320 37912 19320 37912 0 x_end[0]
rlabel metal2 17416 36736 17416 36736 0 x_end[1]
rlabel metal2 14840 37912 14840 37912 0 x_end[2]
rlabel metal2 12040 35560 12040 35560 0 x_end[3]
rlabel metal2 10696 36400 10696 36400 0 x_end[4]
rlabel metal2 8120 37408 8120 37408 0 x_end[5]
rlabel metal2 5824 33992 5824 33992 0 x_end[6]
rlabel metal2 2968 37506 2968 37506 0 x_end[7]
rlabel metal2 36568 37898 36568 37898 0 x_start[0]
rlabel metal2 35112 35168 35112 35168 0 x_start[1]
rlabel metal2 33768 36232 33768 36232 0 x_start[2]
rlabel metal2 30520 35448 30520 35448 0 x_start[3]
rlabel metal2 27496 36568 27496 36568 0 x_start[4]
rlabel metal2 25536 36568 25536 36568 0 x_start[5]
rlabel metal2 23184 36568 23184 36568 0 x_start[6]
rlabel metal2 21560 37912 21560 37912 0 x_start[7]
rlabel metal2 54488 37842 54488 37842 0 y[0]
rlabel metal3 53032 36456 53032 36456 0 y[1]
rlabel metal3 53536 36344 53536 36344 0 y[2]
rlabel metal3 50456 35616 50456 35616 0 y[3]
rlabel metal2 51352 31892 51352 31892 0 y[4]
rlabel metal2 47376 36344 47376 36344 0 y[5]
rlabel metal2 42280 36680 42280 36680 0 y[6]
rlabel metal2 41160 35448 41160 35448 0 y[7]
<< properties >>
string FIXED_BBOX 0 0 60000 40000
<< end >>
