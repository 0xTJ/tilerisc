magic
tech gf180mcuD
magscale 1 5
timestamp 1700139167
<< obsm1 >>
rect 500 500 43686 27388
<< metal2 >>
rect 1872 27588 1928 27988
rect 2222 27588 2278 27988
rect 2672 27588 2728 27988
rect 6722 27588 6778 27988
rect 7072 27588 7128 27988
rect 7272 27588 7328 27988
rect 7497 27588 7553 27988
rect 7722 27588 7778 27988
rect 8022 27588 8078 27988
rect 12122 27588 12178 27988
rect 12522 27588 12578 27988
rect 12872 27588 12928 27988
rect 15472 27588 15528 27988
rect 15972 27588 16028 27988
rect 16372 27588 16428 27988
rect 16672 27588 16728 27988
rect 18422 27588 18478 27988
rect 23284 27588 23340 27988
rect 26472 27588 26528 27988
rect 27322 27588 27378 27988
rect 28172 27588 28228 27988
rect 29622 27588 29678 27988
rect 31672 27588 31728 27988
rect 31872 27588 31928 27988
rect 32472 27588 32528 27988
rect 36522 27588 36578 27988
rect 36872 27588 36928 27988
rect 37072 27588 37128 27988
rect 37272 27588 37328 27988
rect 37472 27588 37528 27988
rect 37822 27588 37878 27988
rect 41922 27588 41978 27988
rect 42322 27588 42378 27988
rect 42672 27588 42728 27988
<< obsm2 >>
rect 500 27558 1842 27636
rect 1958 27558 2192 27636
rect 2308 27558 2642 27636
rect 2758 27558 6692 27636
rect 6808 27558 7042 27636
rect 7158 27558 7242 27636
rect 7358 27558 7467 27636
rect 7583 27558 7692 27636
rect 7808 27558 7992 27636
rect 8108 27558 12092 27636
rect 12208 27558 12492 27636
rect 12608 27558 12842 27636
rect 12958 27558 15442 27636
rect 15558 27558 15942 27636
rect 16058 27558 16342 27636
rect 16458 27558 16642 27636
rect 16758 27558 18392 27636
rect 18508 27558 23254 27636
rect 23370 27558 26442 27636
rect 26558 27558 27292 27636
rect 27408 27558 28142 27636
rect 28258 27558 29592 27636
rect 29708 27558 31642 27636
rect 31758 27558 31842 27636
rect 31958 27558 32442 27636
rect 32558 27558 36492 27636
rect 36608 27558 36842 27636
rect 36958 27558 37042 27636
rect 37158 27558 37242 27636
rect 37358 27558 37442 27636
rect 37558 27558 37792 27636
rect 37908 27558 41892 27636
rect 42008 27558 42292 27636
rect 42408 27558 42642 27636
rect 42758 27558 43686 27636
rect 500 500 43686 27558
<< obsm3 >>
rect 500 500 43686 27388
<< metal4 >>
rect 522 1568 822 26264
rect 922 1568 1222 26264
rect 42863 1568 43163 26264
rect 43263 1568 43563 26264
<< labels >>
rlabel metal2 s 26472 27588 26528 27988 6 A[0]
port 1 nsew signal input
rlabel metal2 s 27322 27588 27378 27988 6 A[1]
port 2 nsew signal input
rlabel metal2 s 28172 27588 28228 27988 6 A[2]
port 3 nsew signal input
rlabel metal2 s 15472 27588 15528 27988 6 A[3]
port 4 nsew signal input
rlabel metal2 s 15972 27588 16028 27988 6 A[4]
port 5 nsew signal input
rlabel metal2 s 16372 27588 16428 27988 6 A[5]
port 6 nsew signal input
rlabel metal2 s 16672 27588 16728 27988 6 A[6]
port 7 nsew signal input
rlabel metal2 s 18422 27588 18478 27988 6 CEN
port 8 nsew signal input
rlabel metal2 s 29622 27588 29678 27988 6 CLK
port 9 nsew signal input
rlabel metal2 s 42672 27588 42728 27988 6 D[0]
port 10 nsew signal input
rlabel metal2 s 37472 27588 37528 27988 6 D[1]
port 11 nsew signal input
rlabel metal2 s 36872 27588 36928 27988 6 D[2]
port 12 nsew signal input
rlabel metal2 s 31672 27588 31728 27988 6 D[3]
port 13 nsew signal input
rlabel metal2 s 12872 27588 12928 27988 6 D[4]
port 14 nsew signal input
rlabel metal2 s 7722 27588 7778 27988 6 D[5]
port 15 nsew signal input
rlabel metal2 s 7072 27588 7128 27988 6 D[6]
port 16 nsew signal input
rlabel metal2 s 1872 27588 1928 27988 6 D[7]
port 17 nsew signal input
rlabel metal2 s 23284 27588 23340 27988 6 GWEN
port 18 nsew signal input
rlabel metal2 s 41922 27588 41978 27988 6 Q[0]
port 19 nsew signal output
rlabel metal2 s 37822 27588 37878 27988 6 Q[1]
port 20 nsew signal output
rlabel metal2 s 36522 27588 36578 27988 6 Q[2]
port 21 nsew signal output
rlabel metal2 s 32472 27588 32528 27988 6 Q[3]
port 22 nsew signal output
rlabel metal2 s 12122 27588 12178 27988 6 Q[4]
port 23 nsew signal output
rlabel metal2 s 8022 27588 8078 27988 6 Q[5]
port 24 nsew signal output
rlabel metal2 s 6722 27588 6778 27988 6 Q[6]
port 25 nsew signal output
rlabel metal2 s 2672 27588 2728 27988 6 Q[7]
port 26 nsew signal output
rlabel metal4 s 522 1568 822 26264 6 VDD
port 27 nsew power bidirectional
rlabel metal4 s 42863 1568 43163 26264 6 VDD
port 27 nsew power bidirectional
rlabel metal4 s 922 1568 1222 26264 6 VSS
port 28 nsew ground bidirectional
rlabel metal4 s 43263 1568 43563 26264 6 VSS
port 28 nsew ground bidirectional
rlabel metal2 s 42322 27588 42378 27988 6 WEN[0]
port 29 nsew signal input
rlabel metal2 s 37272 27588 37328 27988 6 WEN[1]
port 30 nsew signal input
rlabel metal2 s 37072 27588 37128 27988 6 WEN[2]
port 31 nsew signal input
rlabel metal2 s 31872 27588 31928 27988 6 WEN[3]
port 32 nsew signal input
rlabel metal2 s 12522 27588 12578 27988 6 WEN[4]
port 33 nsew signal input
rlabel metal2 s 7497 27588 7553 27988 6 WEN[5]
port 34 nsew signal input
rlabel metal2 s 7272 27588 7328 27988 6 WEN[6]
port 35 nsew signal input
rlabel metal2 s 2222 27588 2278 27988 6 WEN[7]
port 36 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 44486 27988
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2445002
string GDS_FILE /home/thomas/Documents/Projects/tilerisc/openlane/gf180_ram_128x8_wrapper/runs/23_11_16_07_52/results/signoff/gf180_ram_128x8_wrapper.magic.gds
string GDS_START 2348322
<< end >>

