// This is the unpowered netlist.
module tinyrv (clk,
    mem_ld_en,
    mem_st_en,
    inst,
    mem_addr,
    mem_ld_dat,
    mem_ld_mask,
    mem_st_dat,
    mem_st_mask,
    pc,
    pc_next);
 input clk;
 output mem_ld_en;
 output mem_st_en;
 input [31:0] inst;
 output [31:0] mem_addr;
 input [31:0] mem_ld_dat;
 output [3:0] mem_ld_mask;
 output [31:0] mem_st_dat;
 output [3:0] mem_st_mask;
 input [31:0] pc;
 output [31:0] pc_next;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \reg_file.reg_storage[10][0] ;
 wire \reg_file.reg_storage[10][10] ;
 wire \reg_file.reg_storage[10][11] ;
 wire \reg_file.reg_storage[10][12] ;
 wire \reg_file.reg_storage[10][13] ;
 wire \reg_file.reg_storage[10][14] ;
 wire \reg_file.reg_storage[10][15] ;
 wire \reg_file.reg_storage[10][16] ;
 wire \reg_file.reg_storage[10][17] ;
 wire \reg_file.reg_storage[10][18] ;
 wire \reg_file.reg_storage[10][19] ;
 wire \reg_file.reg_storage[10][1] ;
 wire \reg_file.reg_storage[10][20] ;
 wire \reg_file.reg_storage[10][21] ;
 wire \reg_file.reg_storage[10][22] ;
 wire \reg_file.reg_storage[10][23] ;
 wire \reg_file.reg_storage[10][24] ;
 wire \reg_file.reg_storage[10][25] ;
 wire \reg_file.reg_storage[10][26] ;
 wire \reg_file.reg_storage[10][27] ;
 wire \reg_file.reg_storage[10][28] ;
 wire \reg_file.reg_storage[10][29] ;
 wire \reg_file.reg_storage[10][2] ;
 wire \reg_file.reg_storage[10][30] ;
 wire \reg_file.reg_storage[10][31] ;
 wire \reg_file.reg_storage[10][3] ;
 wire \reg_file.reg_storage[10][4] ;
 wire \reg_file.reg_storage[10][5] ;
 wire \reg_file.reg_storage[10][6] ;
 wire \reg_file.reg_storage[10][7] ;
 wire \reg_file.reg_storage[10][8] ;
 wire \reg_file.reg_storage[10][9] ;
 wire \reg_file.reg_storage[11][0] ;
 wire \reg_file.reg_storage[11][10] ;
 wire \reg_file.reg_storage[11][11] ;
 wire \reg_file.reg_storage[11][12] ;
 wire \reg_file.reg_storage[11][13] ;
 wire \reg_file.reg_storage[11][14] ;
 wire \reg_file.reg_storage[11][15] ;
 wire \reg_file.reg_storage[11][16] ;
 wire \reg_file.reg_storage[11][17] ;
 wire \reg_file.reg_storage[11][18] ;
 wire \reg_file.reg_storage[11][19] ;
 wire \reg_file.reg_storage[11][1] ;
 wire \reg_file.reg_storage[11][20] ;
 wire \reg_file.reg_storage[11][21] ;
 wire \reg_file.reg_storage[11][22] ;
 wire \reg_file.reg_storage[11][23] ;
 wire \reg_file.reg_storage[11][24] ;
 wire \reg_file.reg_storage[11][25] ;
 wire \reg_file.reg_storage[11][26] ;
 wire \reg_file.reg_storage[11][27] ;
 wire \reg_file.reg_storage[11][28] ;
 wire \reg_file.reg_storage[11][29] ;
 wire \reg_file.reg_storage[11][2] ;
 wire \reg_file.reg_storage[11][30] ;
 wire \reg_file.reg_storage[11][31] ;
 wire \reg_file.reg_storage[11][3] ;
 wire \reg_file.reg_storage[11][4] ;
 wire \reg_file.reg_storage[11][5] ;
 wire \reg_file.reg_storage[11][6] ;
 wire \reg_file.reg_storage[11][7] ;
 wire \reg_file.reg_storage[11][8] ;
 wire \reg_file.reg_storage[11][9] ;
 wire \reg_file.reg_storage[12][0] ;
 wire \reg_file.reg_storage[12][10] ;
 wire \reg_file.reg_storage[12][11] ;
 wire \reg_file.reg_storage[12][12] ;
 wire \reg_file.reg_storage[12][13] ;
 wire \reg_file.reg_storage[12][14] ;
 wire \reg_file.reg_storage[12][15] ;
 wire \reg_file.reg_storage[12][16] ;
 wire \reg_file.reg_storage[12][17] ;
 wire \reg_file.reg_storage[12][18] ;
 wire \reg_file.reg_storage[12][19] ;
 wire \reg_file.reg_storage[12][1] ;
 wire \reg_file.reg_storage[12][20] ;
 wire \reg_file.reg_storage[12][21] ;
 wire \reg_file.reg_storage[12][22] ;
 wire \reg_file.reg_storage[12][23] ;
 wire \reg_file.reg_storage[12][24] ;
 wire \reg_file.reg_storage[12][25] ;
 wire \reg_file.reg_storage[12][26] ;
 wire \reg_file.reg_storage[12][27] ;
 wire \reg_file.reg_storage[12][28] ;
 wire \reg_file.reg_storage[12][29] ;
 wire \reg_file.reg_storage[12][2] ;
 wire \reg_file.reg_storage[12][30] ;
 wire \reg_file.reg_storage[12][31] ;
 wire \reg_file.reg_storage[12][3] ;
 wire \reg_file.reg_storage[12][4] ;
 wire \reg_file.reg_storage[12][5] ;
 wire \reg_file.reg_storage[12][6] ;
 wire \reg_file.reg_storage[12][7] ;
 wire \reg_file.reg_storage[12][8] ;
 wire \reg_file.reg_storage[12][9] ;
 wire \reg_file.reg_storage[13][0] ;
 wire \reg_file.reg_storage[13][10] ;
 wire \reg_file.reg_storage[13][11] ;
 wire \reg_file.reg_storage[13][12] ;
 wire \reg_file.reg_storage[13][13] ;
 wire \reg_file.reg_storage[13][14] ;
 wire \reg_file.reg_storage[13][15] ;
 wire \reg_file.reg_storage[13][16] ;
 wire \reg_file.reg_storage[13][17] ;
 wire \reg_file.reg_storage[13][18] ;
 wire \reg_file.reg_storage[13][19] ;
 wire \reg_file.reg_storage[13][1] ;
 wire \reg_file.reg_storage[13][20] ;
 wire \reg_file.reg_storage[13][21] ;
 wire \reg_file.reg_storage[13][22] ;
 wire \reg_file.reg_storage[13][23] ;
 wire \reg_file.reg_storage[13][24] ;
 wire \reg_file.reg_storage[13][25] ;
 wire \reg_file.reg_storage[13][26] ;
 wire \reg_file.reg_storage[13][27] ;
 wire \reg_file.reg_storage[13][28] ;
 wire \reg_file.reg_storage[13][29] ;
 wire \reg_file.reg_storage[13][2] ;
 wire \reg_file.reg_storage[13][30] ;
 wire \reg_file.reg_storage[13][31] ;
 wire \reg_file.reg_storage[13][3] ;
 wire \reg_file.reg_storage[13][4] ;
 wire \reg_file.reg_storage[13][5] ;
 wire \reg_file.reg_storage[13][6] ;
 wire \reg_file.reg_storage[13][7] ;
 wire \reg_file.reg_storage[13][8] ;
 wire \reg_file.reg_storage[13][9] ;
 wire \reg_file.reg_storage[14][0] ;
 wire \reg_file.reg_storage[14][10] ;
 wire \reg_file.reg_storage[14][11] ;
 wire \reg_file.reg_storage[14][12] ;
 wire \reg_file.reg_storage[14][13] ;
 wire \reg_file.reg_storage[14][14] ;
 wire \reg_file.reg_storage[14][15] ;
 wire \reg_file.reg_storage[14][16] ;
 wire \reg_file.reg_storage[14][17] ;
 wire \reg_file.reg_storage[14][18] ;
 wire \reg_file.reg_storage[14][19] ;
 wire \reg_file.reg_storage[14][1] ;
 wire \reg_file.reg_storage[14][20] ;
 wire \reg_file.reg_storage[14][21] ;
 wire \reg_file.reg_storage[14][22] ;
 wire \reg_file.reg_storage[14][23] ;
 wire \reg_file.reg_storage[14][24] ;
 wire \reg_file.reg_storage[14][25] ;
 wire \reg_file.reg_storage[14][26] ;
 wire \reg_file.reg_storage[14][27] ;
 wire \reg_file.reg_storage[14][28] ;
 wire \reg_file.reg_storage[14][29] ;
 wire \reg_file.reg_storage[14][2] ;
 wire \reg_file.reg_storage[14][30] ;
 wire \reg_file.reg_storage[14][31] ;
 wire \reg_file.reg_storage[14][3] ;
 wire \reg_file.reg_storage[14][4] ;
 wire \reg_file.reg_storage[14][5] ;
 wire \reg_file.reg_storage[14][6] ;
 wire \reg_file.reg_storage[14][7] ;
 wire \reg_file.reg_storage[14][8] ;
 wire \reg_file.reg_storage[14][9] ;
 wire \reg_file.reg_storage[15][0] ;
 wire \reg_file.reg_storage[15][10] ;
 wire \reg_file.reg_storage[15][11] ;
 wire \reg_file.reg_storage[15][12] ;
 wire \reg_file.reg_storage[15][13] ;
 wire \reg_file.reg_storage[15][14] ;
 wire \reg_file.reg_storage[15][15] ;
 wire \reg_file.reg_storage[15][16] ;
 wire \reg_file.reg_storage[15][17] ;
 wire \reg_file.reg_storage[15][18] ;
 wire \reg_file.reg_storage[15][19] ;
 wire \reg_file.reg_storage[15][1] ;
 wire \reg_file.reg_storage[15][20] ;
 wire \reg_file.reg_storage[15][21] ;
 wire \reg_file.reg_storage[15][22] ;
 wire \reg_file.reg_storage[15][23] ;
 wire \reg_file.reg_storage[15][24] ;
 wire \reg_file.reg_storage[15][25] ;
 wire \reg_file.reg_storage[15][26] ;
 wire \reg_file.reg_storage[15][27] ;
 wire \reg_file.reg_storage[15][28] ;
 wire \reg_file.reg_storage[15][29] ;
 wire \reg_file.reg_storage[15][2] ;
 wire \reg_file.reg_storage[15][30] ;
 wire \reg_file.reg_storage[15][31] ;
 wire \reg_file.reg_storage[15][3] ;
 wire \reg_file.reg_storage[15][4] ;
 wire \reg_file.reg_storage[15][5] ;
 wire \reg_file.reg_storage[15][6] ;
 wire \reg_file.reg_storage[15][7] ;
 wire \reg_file.reg_storage[15][8] ;
 wire \reg_file.reg_storage[15][9] ;
 wire \reg_file.reg_storage[1][0] ;
 wire \reg_file.reg_storage[1][10] ;
 wire \reg_file.reg_storage[1][11] ;
 wire \reg_file.reg_storage[1][12] ;
 wire \reg_file.reg_storage[1][13] ;
 wire \reg_file.reg_storage[1][14] ;
 wire \reg_file.reg_storage[1][15] ;
 wire \reg_file.reg_storage[1][16] ;
 wire \reg_file.reg_storage[1][17] ;
 wire \reg_file.reg_storage[1][18] ;
 wire \reg_file.reg_storage[1][19] ;
 wire \reg_file.reg_storage[1][1] ;
 wire \reg_file.reg_storage[1][20] ;
 wire \reg_file.reg_storage[1][21] ;
 wire \reg_file.reg_storage[1][22] ;
 wire \reg_file.reg_storage[1][23] ;
 wire \reg_file.reg_storage[1][24] ;
 wire \reg_file.reg_storage[1][25] ;
 wire \reg_file.reg_storage[1][26] ;
 wire \reg_file.reg_storage[1][27] ;
 wire \reg_file.reg_storage[1][28] ;
 wire \reg_file.reg_storage[1][29] ;
 wire \reg_file.reg_storage[1][2] ;
 wire \reg_file.reg_storage[1][30] ;
 wire \reg_file.reg_storage[1][31] ;
 wire \reg_file.reg_storage[1][3] ;
 wire \reg_file.reg_storage[1][4] ;
 wire \reg_file.reg_storage[1][5] ;
 wire \reg_file.reg_storage[1][6] ;
 wire \reg_file.reg_storage[1][7] ;
 wire \reg_file.reg_storage[1][8] ;
 wire \reg_file.reg_storage[1][9] ;
 wire \reg_file.reg_storage[2][0] ;
 wire \reg_file.reg_storage[2][10] ;
 wire \reg_file.reg_storage[2][11] ;
 wire \reg_file.reg_storage[2][12] ;
 wire \reg_file.reg_storage[2][13] ;
 wire \reg_file.reg_storage[2][14] ;
 wire \reg_file.reg_storage[2][15] ;
 wire \reg_file.reg_storage[2][16] ;
 wire \reg_file.reg_storage[2][17] ;
 wire \reg_file.reg_storage[2][18] ;
 wire \reg_file.reg_storage[2][19] ;
 wire \reg_file.reg_storage[2][1] ;
 wire \reg_file.reg_storage[2][20] ;
 wire \reg_file.reg_storage[2][21] ;
 wire \reg_file.reg_storage[2][22] ;
 wire \reg_file.reg_storage[2][23] ;
 wire \reg_file.reg_storage[2][24] ;
 wire \reg_file.reg_storage[2][25] ;
 wire \reg_file.reg_storage[2][26] ;
 wire \reg_file.reg_storage[2][27] ;
 wire \reg_file.reg_storage[2][28] ;
 wire \reg_file.reg_storage[2][29] ;
 wire \reg_file.reg_storage[2][2] ;
 wire \reg_file.reg_storage[2][30] ;
 wire \reg_file.reg_storage[2][31] ;
 wire \reg_file.reg_storage[2][3] ;
 wire \reg_file.reg_storage[2][4] ;
 wire \reg_file.reg_storage[2][5] ;
 wire \reg_file.reg_storage[2][6] ;
 wire \reg_file.reg_storage[2][7] ;
 wire \reg_file.reg_storage[2][8] ;
 wire \reg_file.reg_storage[2][9] ;
 wire \reg_file.reg_storage[3][0] ;
 wire \reg_file.reg_storage[3][10] ;
 wire \reg_file.reg_storage[3][11] ;
 wire \reg_file.reg_storage[3][12] ;
 wire \reg_file.reg_storage[3][13] ;
 wire \reg_file.reg_storage[3][14] ;
 wire \reg_file.reg_storage[3][15] ;
 wire \reg_file.reg_storage[3][16] ;
 wire \reg_file.reg_storage[3][17] ;
 wire \reg_file.reg_storage[3][18] ;
 wire \reg_file.reg_storage[3][19] ;
 wire \reg_file.reg_storage[3][1] ;
 wire \reg_file.reg_storage[3][20] ;
 wire \reg_file.reg_storage[3][21] ;
 wire \reg_file.reg_storage[3][22] ;
 wire \reg_file.reg_storage[3][23] ;
 wire \reg_file.reg_storage[3][24] ;
 wire \reg_file.reg_storage[3][25] ;
 wire \reg_file.reg_storage[3][26] ;
 wire \reg_file.reg_storage[3][27] ;
 wire \reg_file.reg_storage[3][28] ;
 wire \reg_file.reg_storage[3][29] ;
 wire \reg_file.reg_storage[3][2] ;
 wire \reg_file.reg_storage[3][30] ;
 wire \reg_file.reg_storage[3][31] ;
 wire \reg_file.reg_storage[3][3] ;
 wire \reg_file.reg_storage[3][4] ;
 wire \reg_file.reg_storage[3][5] ;
 wire \reg_file.reg_storage[3][6] ;
 wire \reg_file.reg_storage[3][7] ;
 wire \reg_file.reg_storage[3][8] ;
 wire \reg_file.reg_storage[3][9] ;
 wire \reg_file.reg_storage[4][0] ;
 wire \reg_file.reg_storage[4][10] ;
 wire \reg_file.reg_storage[4][11] ;
 wire \reg_file.reg_storage[4][12] ;
 wire \reg_file.reg_storage[4][13] ;
 wire \reg_file.reg_storage[4][14] ;
 wire \reg_file.reg_storage[4][15] ;
 wire \reg_file.reg_storage[4][16] ;
 wire \reg_file.reg_storage[4][17] ;
 wire \reg_file.reg_storage[4][18] ;
 wire \reg_file.reg_storage[4][19] ;
 wire \reg_file.reg_storage[4][1] ;
 wire \reg_file.reg_storage[4][20] ;
 wire \reg_file.reg_storage[4][21] ;
 wire \reg_file.reg_storage[4][22] ;
 wire \reg_file.reg_storage[4][23] ;
 wire \reg_file.reg_storage[4][24] ;
 wire \reg_file.reg_storage[4][25] ;
 wire \reg_file.reg_storage[4][26] ;
 wire \reg_file.reg_storage[4][27] ;
 wire \reg_file.reg_storage[4][28] ;
 wire \reg_file.reg_storage[4][29] ;
 wire \reg_file.reg_storage[4][2] ;
 wire \reg_file.reg_storage[4][30] ;
 wire \reg_file.reg_storage[4][31] ;
 wire \reg_file.reg_storage[4][3] ;
 wire \reg_file.reg_storage[4][4] ;
 wire \reg_file.reg_storage[4][5] ;
 wire \reg_file.reg_storage[4][6] ;
 wire \reg_file.reg_storage[4][7] ;
 wire \reg_file.reg_storage[4][8] ;
 wire \reg_file.reg_storage[4][9] ;
 wire \reg_file.reg_storage[5][0] ;
 wire \reg_file.reg_storage[5][10] ;
 wire \reg_file.reg_storage[5][11] ;
 wire \reg_file.reg_storage[5][12] ;
 wire \reg_file.reg_storage[5][13] ;
 wire \reg_file.reg_storage[5][14] ;
 wire \reg_file.reg_storage[5][15] ;
 wire \reg_file.reg_storage[5][16] ;
 wire \reg_file.reg_storage[5][17] ;
 wire \reg_file.reg_storage[5][18] ;
 wire \reg_file.reg_storage[5][19] ;
 wire \reg_file.reg_storage[5][1] ;
 wire \reg_file.reg_storage[5][20] ;
 wire \reg_file.reg_storage[5][21] ;
 wire \reg_file.reg_storage[5][22] ;
 wire \reg_file.reg_storage[5][23] ;
 wire \reg_file.reg_storage[5][24] ;
 wire \reg_file.reg_storage[5][25] ;
 wire \reg_file.reg_storage[5][26] ;
 wire \reg_file.reg_storage[5][27] ;
 wire \reg_file.reg_storage[5][28] ;
 wire \reg_file.reg_storage[5][29] ;
 wire \reg_file.reg_storage[5][2] ;
 wire \reg_file.reg_storage[5][30] ;
 wire \reg_file.reg_storage[5][31] ;
 wire \reg_file.reg_storage[5][3] ;
 wire \reg_file.reg_storage[5][4] ;
 wire \reg_file.reg_storage[5][5] ;
 wire \reg_file.reg_storage[5][6] ;
 wire \reg_file.reg_storage[5][7] ;
 wire \reg_file.reg_storage[5][8] ;
 wire \reg_file.reg_storage[5][9] ;
 wire \reg_file.reg_storage[6][0] ;
 wire \reg_file.reg_storage[6][10] ;
 wire \reg_file.reg_storage[6][11] ;
 wire \reg_file.reg_storage[6][12] ;
 wire \reg_file.reg_storage[6][13] ;
 wire \reg_file.reg_storage[6][14] ;
 wire \reg_file.reg_storage[6][15] ;
 wire \reg_file.reg_storage[6][16] ;
 wire \reg_file.reg_storage[6][17] ;
 wire \reg_file.reg_storage[6][18] ;
 wire \reg_file.reg_storage[6][19] ;
 wire \reg_file.reg_storage[6][1] ;
 wire \reg_file.reg_storage[6][20] ;
 wire \reg_file.reg_storage[6][21] ;
 wire \reg_file.reg_storage[6][22] ;
 wire \reg_file.reg_storage[6][23] ;
 wire \reg_file.reg_storage[6][24] ;
 wire \reg_file.reg_storage[6][25] ;
 wire \reg_file.reg_storage[6][26] ;
 wire \reg_file.reg_storage[6][27] ;
 wire \reg_file.reg_storage[6][28] ;
 wire \reg_file.reg_storage[6][29] ;
 wire \reg_file.reg_storage[6][2] ;
 wire \reg_file.reg_storage[6][30] ;
 wire \reg_file.reg_storage[6][31] ;
 wire \reg_file.reg_storage[6][3] ;
 wire \reg_file.reg_storage[6][4] ;
 wire \reg_file.reg_storage[6][5] ;
 wire \reg_file.reg_storage[6][6] ;
 wire \reg_file.reg_storage[6][7] ;
 wire \reg_file.reg_storage[6][8] ;
 wire \reg_file.reg_storage[6][9] ;
 wire \reg_file.reg_storage[7][0] ;
 wire \reg_file.reg_storage[7][10] ;
 wire \reg_file.reg_storage[7][11] ;
 wire \reg_file.reg_storage[7][12] ;
 wire \reg_file.reg_storage[7][13] ;
 wire \reg_file.reg_storage[7][14] ;
 wire \reg_file.reg_storage[7][15] ;
 wire \reg_file.reg_storage[7][16] ;
 wire \reg_file.reg_storage[7][17] ;
 wire \reg_file.reg_storage[7][18] ;
 wire \reg_file.reg_storage[7][19] ;
 wire \reg_file.reg_storage[7][1] ;
 wire \reg_file.reg_storage[7][20] ;
 wire \reg_file.reg_storage[7][21] ;
 wire \reg_file.reg_storage[7][22] ;
 wire \reg_file.reg_storage[7][23] ;
 wire \reg_file.reg_storage[7][24] ;
 wire \reg_file.reg_storage[7][25] ;
 wire \reg_file.reg_storage[7][26] ;
 wire \reg_file.reg_storage[7][27] ;
 wire \reg_file.reg_storage[7][28] ;
 wire \reg_file.reg_storage[7][29] ;
 wire \reg_file.reg_storage[7][2] ;
 wire \reg_file.reg_storage[7][30] ;
 wire \reg_file.reg_storage[7][31] ;
 wire \reg_file.reg_storage[7][3] ;
 wire \reg_file.reg_storage[7][4] ;
 wire \reg_file.reg_storage[7][5] ;
 wire \reg_file.reg_storage[7][6] ;
 wire \reg_file.reg_storage[7][7] ;
 wire \reg_file.reg_storage[7][8] ;
 wire \reg_file.reg_storage[7][9] ;
 wire \reg_file.reg_storage[8][0] ;
 wire \reg_file.reg_storage[8][10] ;
 wire \reg_file.reg_storage[8][11] ;
 wire \reg_file.reg_storage[8][12] ;
 wire \reg_file.reg_storage[8][13] ;
 wire \reg_file.reg_storage[8][14] ;
 wire \reg_file.reg_storage[8][15] ;
 wire \reg_file.reg_storage[8][16] ;
 wire \reg_file.reg_storage[8][17] ;
 wire \reg_file.reg_storage[8][18] ;
 wire \reg_file.reg_storage[8][19] ;
 wire \reg_file.reg_storage[8][1] ;
 wire \reg_file.reg_storage[8][20] ;
 wire \reg_file.reg_storage[8][21] ;
 wire \reg_file.reg_storage[8][22] ;
 wire \reg_file.reg_storage[8][23] ;
 wire \reg_file.reg_storage[8][24] ;
 wire \reg_file.reg_storage[8][25] ;
 wire \reg_file.reg_storage[8][26] ;
 wire \reg_file.reg_storage[8][27] ;
 wire \reg_file.reg_storage[8][28] ;
 wire \reg_file.reg_storage[8][29] ;
 wire \reg_file.reg_storage[8][2] ;
 wire \reg_file.reg_storage[8][30] ;
 wire \reg_file.reg_storage[8][31] ;
 wire \reg_file.reg_storage[8][3] ;
 wire \reg_file.reg_storage[8][4] ;
 wire \reg_file.reg_storage[8][5] ;
 wire \reg_file.reg_storage[8][6] ;
 wire \reg_file.reg_storage[8][7] ;
 wire \reg_file.reg_storage[8][8] ;
 wire \reg_file.reg_storage[8][9] ;
 wire \reg_file.reg_storage[9][0] ;
 wire \reg_file.reg_storage[9][10] ;
 wire \reg_file.reg_storage[9][11] ;
 wire \reg_file.reg_storage[9][12] ;
 wire \reg_file.reg_storage[9][13] ;
 wire \reg_file.reg_storage[9][14] ;
 wire \reg_file.reg_storage[9][15] ;
 wire \reg_file.reg_storage[9][16] ;
 wire \reg_file.reg_storage[9][17] ;
 wire \reg_file.reg_storage[9][18] ;
 wire \reg_file.reg_storage[9][19] ;
 wire \reg_file.reg_storage[9][1] ;
 wire \reg_file.reg_storage[9][20] ;
 wire \reg_file.reg_storage[9][21] ;
 wire \reg_file.reg_storage[9][22] ;
 wire \reg_file.reg_storage[9][23] ;
 wire \reg_file.reg_storage[9][24] ;
 wire \reg_file.reg_storage[9][25] ;
 wire \reg_file.reg_storage[9][26] ;
 wire \reg_file.reg_storage[9][27] ;
 wire \reg_file.reg_storage[9][28] ;
 wire \reg_file.reg_storage[9][29] ;
 wire \reg_file.reg_storage[9][2] ;
 wire \reg_file.reg_storage[9][30] ;
 wire \reg_file.reg_storage[9][31] ;
 wire \reg_file.reg_storage[9][3] ;
 wire \reg_file.reg_storage[9][4] ;
 wire \reg_file.reg_storage[9][5] ;
 wire \reg_file.reg_storage[9][6] ;
 wire \reg_file.reg_storage[9][7] ;
 wire \reg_file.reg_storage[9][8] ;
 wire \reg_file.reg_storage[9][9] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A3 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__I (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__I (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__I (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__I (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I0 (.I(\reg_file.reg_storage[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I1 (.I(\reg_file.reg_storage[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I2 (.I(\reg_file.reg_storage[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I3 (.I(\reg_file.reg_storage[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__S0 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__S1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__I (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__S (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__S (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__I0 (.I(\reg_file.reg_storage[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__I1 (.I(\reg_file.reg_storage[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__I2 (.I(\reg_file.reg_storage[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__I3 (.I(\reg_file.reg_storage[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__S0 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__S1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I0 (.I(\reg_file.reg_storage[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I1 (.I(\reg_file.reg_storage[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I2 (.I(\reg_file.reg_storage[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I3 (.I(\reg_file.reg_storage[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__S0 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__S1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__S0 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__S1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__I (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__I0 (.I(\reg_file.reg_storage[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__S1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__S (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__S (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__S1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__I3 (.I(\reg_file.reg_storage[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__S1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__S (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__S (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__S (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__S0 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__S0 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__C (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__I (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__I1 (.I(\reg_file.reg_storage[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__I3 (.I(\reg_file.reg_storage[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__S0 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__S (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__S1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__I (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__S0 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__S0 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__S1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__S (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__S (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__S (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__S1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__C (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__I (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__I (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__I (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__S0 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__S (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__S0 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__S0 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__I (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__S0 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__S1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__I (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__I (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__I (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__I0 (.I(\reg_file.reg_storage[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__S0 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__S1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__S (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__S (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__I (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__S0 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__S1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__S0 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__S1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__S0 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__S1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__S0 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__S1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__S (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__S (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__S0 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__S1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__S0 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__S1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__S0 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__S1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__I (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A3 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__I (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__I (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__I (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A3 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__I (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A3 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__I (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__I0 (.I(\reg_file.reg_storage[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__I1 (.I(\reg_file.reg_storage[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__I2 (.I(\reg_file.reg_storage[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__I3 (.I(\reg_file.reg_storage[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__S0 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__S1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__I (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__S (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__I (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__S (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__I (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__I0 (.I(\reg_file.reg_storage[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__I1 (.I(\reg_file.reg_storage[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__I2 (.I(\reg_file.reg_storage[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__I3 (.I(\reg_file.reg_storage[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__S0 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__S1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__I0 (.I(\reg_file.reg_storage[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__I1 (.I(\reg_file.reg_storage[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__I2 (.I(\reg_file.reg_storage[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__I3 (.I(\reg_file.reg_storage[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__S0 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__S1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__S0 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__S1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A3 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__I (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__I (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__B (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A2 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A3 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__I (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__I (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__B2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__I (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__I (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__I (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__I (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__B (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__I (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__I (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__I (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__B2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__I (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__I (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__B (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__I (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__I (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__B2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__I (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__I (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__I (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__I (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__S0 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__S1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__I (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__I (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__I (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__I (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__I (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__B (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__I (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__I (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__I (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__S0 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__S1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__S0 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__S1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__I (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__I (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__S0 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__S1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__I (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__I (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__I (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__I (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__I (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__S0 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__S1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__I (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__I (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__I (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__B (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__I (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__I (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__S0 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__S1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__S0 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__S1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__I (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__S0 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__S1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__I (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__S0 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__S1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__S (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__S (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__I (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__S0 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__S1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__S0 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__S1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__S0 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__S1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__B (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__I (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__I (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__I (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__I (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__I (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__I3 (.I(\reg_file.reg_storage[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__S0 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__S1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__I (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A2 (.I(\reg_file.reg_storage[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__B (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__I (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__I (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__I0 (.I(\reg_file.reg_storage[12][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__S0 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__S1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__S0 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__S1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__S0 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__S1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__I (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__I (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__I0 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I0 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__S (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__I (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__I (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__I (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__S0 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__I (.I(\reg_file.reg_storage[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__I (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__I (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__B (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__I (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__I2 (.I(\reg_file.reg_storage[14][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__I3 (.I(\reg_file.reg_storage[15][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__S0 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__S1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__S0 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__S1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__B1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__B2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__I (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A2 (.I(\reg_file.reg_storage[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__I (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__I (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__S0 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__S1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__S0 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__S1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__S0 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__S1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__B (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__B (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__B1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__B2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__S1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__I (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__S (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__I (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__S (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__S1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__I1 (.I(\reg_file.reg_storage[9][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__S1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__S0 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__S1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A3 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A1 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__I (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__S0 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__S1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__I (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__I (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__I (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__B (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__S0 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__S1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__S0 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__S1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__I (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__I2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__S0 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__S1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__I (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__I0 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__I0 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__S (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__S (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__I (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__S0 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__S1 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__B (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__I (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__I0 (.I(\reg_file.reg_storage[12][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__I1 (.I(\reg_file.reg_storage[13][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__S0 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__S1 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__S0 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__S1 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__I0 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__I3 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__S0 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__S1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__S0 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__S1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__B (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__S0 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__S1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__S0 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__S1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__I0 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__I3 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__S0 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__S1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__I3 (.I(\reg_file.reg_storage[7][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__S0 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__S1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__B (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__I (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__S0 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__S1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__I0 (.I(\reg_file.reg_storage[8][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__I1 (.I(\reg_file.reg_storage[9][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__I2 (.I(\reg_file.reg_storage[10][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__I3 (.I(\reg_file.reg_storage[11][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__S0 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__S1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__I2 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__S0 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__S1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A2 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__I (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__I3 (.I(\reg_file.reg_storage[7][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__S0 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__S1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__B (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__I1 (.I(\reg_file.reg_storage[13][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__S0 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__S1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__I0 (.I(\reg_file.reg_storage[8][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__I1 (.I(\reg_file.reg_storage[9][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__I3 (.I(\reg_file.reg_storage[11][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__S0 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__S1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__S0 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__S1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__S (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__I (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__I3 (.I(\reg_file.reg_storage[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__S0 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__S1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__S (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__S (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__I1 (.I(\reg_file.reg_storage[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__S0 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__S1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__S0 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__S1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__I0 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__I2 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__I3 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__S0 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__S1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__B1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__B2 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__I (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__I (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__I3 (.I(\reg_file.reg_storage[7][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__S0 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__S1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__S (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__S (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I0 (.I(\reg_file.reg_storage[12][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I1 (.I(\reg_file.reg_storage[13][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I2 (.I(\reg_file.reg_storage[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__S0 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__S1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__S0 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__S1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__I3 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__S0 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__S1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A3 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__I3 (.I(\reg_file.reg_storage[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__S0 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__S1 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__B (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__I1 (.I(\reg_file.reg_storage[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__S0 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__S1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__S0 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__S1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__I3 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__S0 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__S1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A2 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A1 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__I3 (.I(\reg_file.reg_storage[7][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__S0 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__S1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__B (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I0 (.I(\reg_file.reg_storage[12][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I1 (.I(\reg_file.reg_storage[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I2 (.I(\reg_file.reg_storage[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__S0 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__S1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__S0 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__S1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__I0 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__I3 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__S0 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__S1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__I (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__S (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__S (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__I (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__I0 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__I (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__I (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__I0 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__I1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__S (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__I (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__I (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__I (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__I (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A1 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__I (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__I (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__S0 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__S1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__S (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__I0 (.I(\reg_file.reg_storage[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__S (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__S0 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__S1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__S0 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__S1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__S0 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__S1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A3 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__I (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__S0 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__S1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A1 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__B (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__S0 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__S1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__S0 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__S1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__S0 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__S1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__S0 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__S1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__I (.I(\reg_file.reg_storage[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__B (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__S0 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__S1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__S0 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__S1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__I0 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__I2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__I3 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__S0 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__S1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__S0 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__S1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__B (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__S0 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__S1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__S0 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__S1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__S0 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__S1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__S (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__I (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__S0 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__S1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__S (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__S (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__S0 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__S1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__S0 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__S1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__S0 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__S1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__I (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__S0 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__S1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A1 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__B (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__S0 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__S1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__S0 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__S1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__S0 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__S1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A2 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__S0 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__S1 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__S (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__S (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__S0 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__S1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__S0 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__S1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__S0 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__S1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__A3 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__I (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__S0 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__S1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__S (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__S (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__S0 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__S1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__S0 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__S1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__S0 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__S1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__I (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__I (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__S (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__I0 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__I0 (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__I1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__I (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__I (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__S0 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__S1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__S (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__S (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__S0 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__S1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__S0 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__S1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__S0 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__S1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__I (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__I (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__I (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__S1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__B (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__A2 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__S1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__I0 (.I(\reg_file.reg_storage[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__S1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__S0 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__S1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__I (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__I (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__S0 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__S1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__S (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__S (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__S0 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__S1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__S0 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__S1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__S0 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__S1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__I (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__S0 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__S1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__S (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__S (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__S0 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__S1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__S0 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__S1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__S0 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__S1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__I (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__I (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__I (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__S0 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__S (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__S0 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__I3 (.I(\reg_file.reg_storage[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__S0 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__S0 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__S1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__I (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__S0 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__S1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__B (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__S0 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__S1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__I1 (.I(\reg_file.reg_storage[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__I3 (.I(\reg_file.reg_storage[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__S0 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__S1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__I2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__S0 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__S1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__S0 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__S1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__S0 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__S1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__I0 (.I(\reg_file.reg_storage[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__S0 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__S1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__I0 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__S0 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__S1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A2 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__I (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__C (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__B (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__I (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A4 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__I1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__I (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__I (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__I (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__I (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__I (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__I (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__I3 (.I(\reg_file.reg_storage[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__S0 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__S1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__S (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__S (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__I (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__I1 (.I(\reg_file.reg_storage[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__S0 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__S1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__S0 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__S1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__I3 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__S1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__I (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__I (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__I0 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__I (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__I3 (.I(\reg_file.reg_storage[7][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__S0 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__S1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__I (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__S (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__S (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__I0 (.I(\reg_file.reg_storage[12][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__I1 (.I(\reg_file.reg_storage[13][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__I2 (.I(\reg_file.reg_storage[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__S0 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__S1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__S0 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__S1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__I3 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__S1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__C (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__I (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__I1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__I (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A3 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A4 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__I (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__I3 (.I(\reg_file.reg_storage[7][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__S0 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__S1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__I (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__I (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__I (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__I (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__B (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A1 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__I0 (.I(\reg_file.reg_storage[12][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__I1 (.I(\reg_file.reg_storage[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__I2 (.I(\reg_file.reg_storage[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__S0 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__S1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__S0 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__S1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__S0 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__S1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A3 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__I3 (.I(\reg_file.reg_storage[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__S0 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__S1 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__S (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__S (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__I1 (.I(\reg_file.reg_storage[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__S0 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__S1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__S0 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__S1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__I2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__I3 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__S0 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__S1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__I (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__I (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__I3 (.I(\reg_file.reg_storage[7][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__S0 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__S1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__I (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__S0 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__S1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__I0 (.I(\reg_file.reg_storage[8][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__I1 (.I(\reg_file.reg_storage[9][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__I2 (.I(\reg_file.reg_storage[10][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__I3 (.I(\reg_file.reg_storage[11][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__S0 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__S1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__S0 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__S1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A2 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__I (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__I3 (.I(\reg_file.reg_storage[7][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__S0 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__S1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__I1 (.I(\reg_file.reg_storage[13][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__S0 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__S1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__I0 (.I(\reg_file.reg_storage[8][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__I1 (.I(\reg_file.reg_storage[9][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__I3 (.I(\reg_file.reg_storage[11][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__S0 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__S1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__S0 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__S1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__S0 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__S1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__S0 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__S1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__S0 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__S1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__I1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__S0 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__S1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__S0 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__S1 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__I0 (.I(\reg_file.reg_storage[12][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__I1 (.I(\reg_file.reg_storage[13][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__S0 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__S1 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__S0 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__S1 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__S0 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__S1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A2 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__I0 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__S (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__I (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__I (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__I (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__I (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__S0 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__S1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__I (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__S0 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__S1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A2 (.I(\reg_file.reg_storage[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__B2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__I0 (.I(\reg_file.reg_storage[12][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__S0 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__S1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__I3 (.I(\reg_file.reg_storage[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__S0 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__S1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__S0 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__S1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A1 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__I0 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__I0 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__S0 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__S1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__S (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__S0 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__S0 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__S0 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__S1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A2 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A2 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__I0 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__I1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__S0 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__S (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__S0 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__S0 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__S0 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__S1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A3 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A2 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A3 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A3 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__B (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__I (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__S0 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__S1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__I (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__S (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__I0 (.I(\reg_file.reg_storage[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__S (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__S0 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__S1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__S0 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__S1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__I (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__I (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__S0 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__S1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A2 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I0 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__I (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__I (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__I (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__I (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__I (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__I1 (.I(\reg_file.reg_storage[9][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__S0 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__S1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__I (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__S (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__S (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__I (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__I (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__S0 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__S1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__S0 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__S1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__S0 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__S1 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A3 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A2 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__I (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__S0 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__S1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__S (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__I0 (.I(\reg_file.reg_storage[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__S (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__I2 (.I(\reg_file.reg_storage[14][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__I3 (.I(\reg_file.reg_storage[15][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__S0 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__S1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__S0 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__S1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__S0 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__S1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A3 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__B (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__S0 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__S1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__S (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__S (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__S0 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__S1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__I (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__S0 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__S1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__S0 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__S1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A2 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A3 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__I (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__S0 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__S (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__S0 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__S1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__S0 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__S1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__S0 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__S1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__I (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__I (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__S0 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__S1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__S (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__S (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__S0 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__S0 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__S0 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__S1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__S0 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__S1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__S (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__I0 (.I(\reg_file.reg_storage[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__S (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__S0 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__S1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__S0 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__S1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__S0 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__S1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A2 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__I (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__I1 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__S (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__I (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__S1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__S (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__S (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__S1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__S1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__S0 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__S1 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A2 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__C (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__S0 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__S1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__S (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__I0 (.I(\reg_file.reg_storage[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__I1 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__S (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__S0 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__S1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__S0 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__S1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__S0 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__S1 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__S0 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__S1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__S (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__S (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__S0 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__S1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__S0 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__S1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__S0 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__S1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A2 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__I (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__S0 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__S1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__S (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__S (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__S0 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__S1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__S0 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__S1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__S0 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__S1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A2 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A2 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__S0 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__S1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__S (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__S (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__S0 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__S1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__S0 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__S1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__S0 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__S1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A4 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A2 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A2 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__I0 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__I1 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__I (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A2 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A2 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A2 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A3 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__I (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A2 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A2 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__B2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__B2 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__B (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A2 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A3 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A3 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__B1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__B2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__I (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__I (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A2 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__I0 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__I1 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__B1 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__B2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__B (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__I (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__I (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__I (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__I (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A1 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__B (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__I0 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__I1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A2 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A2 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A3 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__I (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__S (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__S (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__I1 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__S (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__C (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A1 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__I (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A1 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A2 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A3 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__S (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__C (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A2 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A1 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__I (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__I (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__I (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__I (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__I (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__I (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__I (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__I (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__I (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__S (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__I (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__S (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A2 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A2 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__I (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__I (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A1 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__I (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__C (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A3 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__I (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__I (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__I (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__I (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__S (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__I (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__I (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__I (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__B (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A2 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__I (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__I (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__B (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__I (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A1 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__B2 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A1 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__I (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__I (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A3 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__B1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__B3 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__S (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A1 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__I (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__I (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A2 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__I (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__S (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__I1 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__I (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__B (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A1 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__B (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A1 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__S (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__B (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__B1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__B2 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A1 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__B (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__I (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A3 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A4 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A3 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A2 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__B (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__I (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__B (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__I (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__I (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__I (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__I (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A2 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__I (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__S (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A2 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A2 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__I (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A2 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__B (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__B (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A3 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__I (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__I0 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__I1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__S (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A2 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A1 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__C (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__S (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__I0 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A1 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A2 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A1 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A2 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__B (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__B (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A2 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__I (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__I (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A2 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A2 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__I (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__I (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__A1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__I0 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__S (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__A2 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__I (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A2 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__I (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A2 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__A1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__A2 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A2 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__B (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__C (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A1 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__B (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__I (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__I0 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__I (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__B1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A1 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__B2 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__I (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__I (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A2 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__S (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A1 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A2 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__I (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__I (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__B (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__I (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__C (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__I (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__I (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__I (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A2 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__S (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A1 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__B1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A2 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__I (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A1 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A2 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A1 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__I (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__I (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__I (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A1 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__B (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A1 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A2 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A2 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A2 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A2 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A2 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__I (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__B (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__B (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__B2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__I (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__B1 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__B2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A1 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__I (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A1 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A1 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A2 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__I (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__B (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A2 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A2 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A2 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A1 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__B (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A1 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A3 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A1 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__B1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A2 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__B (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A1 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__B (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__I (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__I (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__C2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A2 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A1 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__B (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A2 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A2 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A1 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A2 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__S (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__A2 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A2 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__A1 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__B1 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__B2 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__I (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A2 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__I (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__I (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__I0 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__I1 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__I (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__B (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A1 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A2 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__A2 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__B (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__B (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__I (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__I (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A1 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__A2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__I0 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__I1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__S (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__I0 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__I1 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__B (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__B1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__I (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__I (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__B (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__I0 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__A1 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__A2 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__I0 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__I1 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A3 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__B1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__B2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__C (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__A1 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__A2 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__I (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__I (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__A2 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__B (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__A2 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__I (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__I (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__I (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__I (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__A2 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__I0 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__I1 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__S (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__S (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__A2 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__A1 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__I (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A2 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A2 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__A2 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A2 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__A2 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A1 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__C1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__I (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A2 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__B2 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A1 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__A2 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A1 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__I (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A2 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__S (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__I0 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__I1 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A2 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__A1 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__I (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__A2 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__A1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__A2 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A2 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A2 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A1 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__A1 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__B1 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A2 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__B1 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__A2 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A2 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__A2 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__A2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__A2 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A1 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A1 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A2 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__I0 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__I1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__S (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A3 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__I (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__A1 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__A2 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A1 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__A1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A1 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A2 (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A3 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__A2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__B (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__A2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__B1 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__B2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__A1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__I (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A1 (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__A1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__I0 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__S (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A2 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A2 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__A2 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__B1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A2 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__B (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__B (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__I (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__A2 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A1 (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A2 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A2 (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__A1 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A2 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__B1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__A2 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__B (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__B (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A2 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__A2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__I (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__A1 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__A2 (.I(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A1 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A2 (.I(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A1 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A2 (.I(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A2 (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A1 (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__A1 (.I(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A1 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A1 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A1 (.I(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__A1 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A2 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A2 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__I0 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__I1 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A1 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A2 (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__I (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A2 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__B (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__I (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A1 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__S (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__C (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__A2 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A2 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A1 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A1 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__A1 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__A1 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__I (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__A1 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__A1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__A2 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A2 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__A2 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A2 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A1 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A2 (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__A1 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A1 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A1 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__A1 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__B (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A3 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__B (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__C (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__A1 (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__A2 (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__B (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__A2 (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A2 (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__B (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__B1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__B (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__C (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A2 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A1 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A2 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__B (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__A2 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__B1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__B2 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__I (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__I (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A2 (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A3 (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__I (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A1 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A2 (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__A1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__I (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A3 (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A1 (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A1 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__A1 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__A1 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__A1 (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A1 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A1 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A1 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A1 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A1 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A1 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A1 (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A1 (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A1 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__I (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A1 (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A1 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A1 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A3 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A2 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A1 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A1 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A1 (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A1 (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__B2 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__A1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__B2 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__B2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A1 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__B2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__A1 (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__B2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__B2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A1 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__B2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__B2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A1 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A3 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A1 (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A2 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__B (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__A1 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A1 (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7181__B (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__B (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__I (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A1 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__I (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__I (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__A2 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__A1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A1 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A2 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__A2 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__B2 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__A1 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A2 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__B2 (.I(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A2 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__A1 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__I (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__A2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__B2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A1 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A2 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A3 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__A2 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__B2 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__B2 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__A2 (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__A2 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A2 (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__A2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__B2 (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__A2 (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__A2 (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A2 (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__B1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__B2 (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__A2 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A2 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__I (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A3 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A2 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A3 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A1 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__B1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__B2 (.I(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7313__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__A2 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__A2 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__A2 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__A2 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7338__A2 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__A2 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A1 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__I (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__A2 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__A2 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A2 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A2 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A2 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__A2 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A2 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__A2 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__A2 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__A2 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A2 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__A2 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__A2 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__A2 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__A2 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A2 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7394__A2 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__A2 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__A2 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7401__A2 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7402__B1 (.I(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A1 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__A2 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__A2 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__A2 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__A2 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A2 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__A2 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__I (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__A2 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__A2 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__A2 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__A2 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__A2 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__A2 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A2 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__A2 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7453__A1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__A2 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__A2 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__I (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__A2 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__A2 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__A2 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__A2 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__A2 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__A1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__A2 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7500__I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A1 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A2 (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__A2 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__I (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7532__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__A2 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__B1 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7537__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__A2 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__B1 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__A2 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__A3 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__A2 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A2 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7562__A2 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7562__A4 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__A2 (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__A2 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__B (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__I (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A1 (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A2 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7583__I (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__I1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__A2 (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__I (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__A2 (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__B1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__B2 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__C (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__I (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A1 (.I(\reg_file.reg_storage[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__A2 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A3 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__A1 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__I (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__I (.I(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__I2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__I3 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__A1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__B1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__C (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__A1 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__I (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__I (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__A2 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__A1 (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__I (.I(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__A1 (.I(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__B1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__B2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A2 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__B1 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__B2 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__C (.I(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__I (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7639__I (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7641__S (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__I2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__I3 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__A2 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__B1 (.I(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7652__I (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__I (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__S (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__A1 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__A2 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__B (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__I2 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__I3 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__A1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__A1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__B1 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__B2 (.I(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__I (.I(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__A2 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A1 (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__I2 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__I3 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__I (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A1 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A2 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__B1 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__I (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__S (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__I2 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__I3 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__A1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7683__I (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7684__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7684__A2 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__A2 (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__B1 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__B2 (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__I (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A2 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7690__A1 (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7693__I1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__A2 (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A1 (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__B1 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__B2 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A2 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__I (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__S (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__I (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7707__B (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A1 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__A2 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__B1 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__A1 (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__A2 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__A1 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__A2 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__I (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__S (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__I1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__B (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A2 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__B2 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__C (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__A1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__B1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__B2 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__I (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A2 (.I(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A1 (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__A1 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__I (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A1 (.I(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A1 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__A2 (.I(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A1 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__B (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__A1 (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__A2 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__I (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__S (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__I1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7751__B (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A1 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A1 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__B1 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__B2 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__C (.I(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A1 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A2 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__I (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__S (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A1 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__I (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__A1 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__B1 (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__B2 (.I(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__I (.I(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__I (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__S (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A1 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A2 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__B1 (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__B2 (.I(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__I (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__S (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__I (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7796__I1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__B (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__A2 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__B (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__A1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__B2 (.I(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__I (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7806__A2 (.I(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A1 (.I(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A2 (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__A2 (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A1 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__A2 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__A1 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__A2 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__B (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__I (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__S (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__A1 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__A2 (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__I (.I(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A2 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__B2 (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__I (.I(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A2 (.I(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A1 (.I(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A2 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__A4 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A1 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A2 (.I(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__B2 (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__I (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__A2 (.I(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__A1 (.I(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__A1 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A2 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__A1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__B2 (.I(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__I (.I(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__A2 (.I(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A1 (.I(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__I (.I(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__A4 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__B2 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__A1 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__B2 (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__I (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A2 (.I(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__A1 (.I(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A4 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__A2 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__B2 (.I(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__A2 (.I(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A1 (.I(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A4 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__A1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__B1 (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__B2 (.I(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__A2 (.I(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A1 (.I(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A2 (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__A4 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__B (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__B1 (.I(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__B2 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__A2 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__A1 (.I(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A4 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__B (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__A2 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A2 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__B1 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__B2 (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__A2 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__A1 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__I (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__I (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__I (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__B2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__A1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__B2 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__C (.I(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__I (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A2 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__B2 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__B2 (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__C (.I(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__A2 (.I(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A1 (.I(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__I (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A2 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__A1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__B2 (.I(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__C (.I(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A2 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__B1 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__B2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__A1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__B2 (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__C (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__I (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__A2 (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__I (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__I (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__A1 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A2 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__C (.I(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__I (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A2 (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A1 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__A2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__B2 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__C (.I(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__I (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__A2 (.I(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__A2 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__A1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__C (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__I (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A2 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A2 (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__B1 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__B2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__A1 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__B2 (.I(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__C (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__I (.I(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__A2 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__A1 (.I(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__A2 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__A1 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__I (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7974__A3 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A1 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A3 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__I (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__A2 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__I (.I(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__S (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__S (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__A2 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__S (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__A2 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__S (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__S (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__A2 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__A2 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__S (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__S (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__S (.I(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8008__S (.I(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__I (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__A2 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__A1 (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__A2 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__S (.I(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__A2 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A1 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A2 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A2 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__A2 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__A2 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__A2 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__I (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__A2 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8024__A2 (.I(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__A2 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__A2 (.I(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8027__A2 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A1 (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A2 (.I(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8029__A2 (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A2 (.I(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__A2 (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__A1 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__A1 (.I(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8038__A2 (.I(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__A2 (.I(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A1 (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__A2 (.I(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__A1 (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__A2 (.I(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__A1 (.I(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__A1 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__A1 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A3 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__I (.I(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A1 (.I(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A2 (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__A2 (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A1 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A2 (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__A1 (.I(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__A2 (.I(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__I (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__I (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__I (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__I (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A2 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__I (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__I (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__S (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__S (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__A2 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__S (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A2 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__I (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__S (.I(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__S (.I(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__I (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__A2 (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__A2 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__S (.I(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__S (.I(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__S (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__S (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__I (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__A2 (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__A1 (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__S (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__A2 (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A1 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__A2 (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__I (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__A2 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__I (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__A2 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A2 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__A2 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__A2 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__A2 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__A1 (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__A2 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A2 (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__A2 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__A1 (.I(\reg_file.reg_storage[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__A2 (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__A2 (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__A1 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__A2 (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__A2 (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__A1 (.I(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__A2 (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A2 (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__A1 (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A1 (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A1 (.I(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__A1 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A1 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A2 (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__A1 (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__A2 (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__A1 (.I(\reg_file.reg_storage[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A1 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A1 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A2 (.I(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__I (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__I (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__A2 (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__I (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__S (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__S (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A2 (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__S (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__A2 (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__I (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__S (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__S (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__I (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__A2 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__A2 (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__S (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__S (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__S (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__S (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__I (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__A2 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A1 (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A2 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__S (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A2 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__A1 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__A2 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__A2 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A2 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__I (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__A2 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__I (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A1 (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__A2 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A2 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__A1 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__A1 (.I(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__A1 (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__A1 (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A1 (.I(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A1 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__A1 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__I (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8220__I (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A1 (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A2 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__I (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__I (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__A1 (.I(\reg_file.reg_storage[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__A2 (.I(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__I (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__A1 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__A2 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__I (.I(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__I (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__A2 (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__A2 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__I (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__I (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__I0 (.I(\reg_file.reg_storage[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__S (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__I (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__I1 (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__S (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__I (.I(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8246__A2 (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A2 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__I (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__S (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__I (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__A2 (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A2 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__I (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8256__I (.I(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__S (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__I (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__S (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__I (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__I (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8264__I (.I(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__A2 (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__A2 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__I (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8268__S (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__I (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__S (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__I (.I(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__S (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__I (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__S (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__I (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__I (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__A2 (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A2 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__S (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8287__I (.I(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__A2 (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__A2 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8291__I (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__A2 (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8294__A2 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__I (.I(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__I (.I(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__A2 (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8299__A2 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__I (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__I (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A2 (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__A2 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A2 (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__A2 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__I (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__A2 (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__A2 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__A2 (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__A2 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A1 (.I(\reg_file.reg_storage[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A2 (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8320__A2 (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__I (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__I (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__A1 (.I(\reg_file.reg_storage[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A1 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A2 (.I(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__I (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__A1 (.I(\reg_file.reg_storage[7][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__A2 (.I(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__I (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__I (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8332__A1 (.I(\reg_file.reg_storage[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A1 (.I(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A2 (.I(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__I (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__I (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__A1 (.I(\reg_file.reg_storage[7][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__I (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__I (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__I (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__I (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8347__I (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__I (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__A1 (.I(\reg_file.reg_storage[7][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__I (.I(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__I (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A1 (.I(\reg_file.reg_storage[7][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A1 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A1 (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A2 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8357__I (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__I (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__A1 (.I(\reg_file.reg_storage[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A1 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__A1 (.I(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__I (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__I (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8368__A2 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__A2 (.I(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__I (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__S (.I(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__I1 (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__S (.I(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__A2 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__A2 (.I(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__S (.I(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__A2 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__A2 (.I(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__I (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__S (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__S (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__I (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A2 (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8389__A2 (.I(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__S (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__S (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__S (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__S (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8398__I (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__A2 (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__A2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__S (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__A2 (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A1 (.I(\reg_file.reg_storage[14][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A2 (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__A2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__I (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__A2 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__A2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__I (.I(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__A2 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__A2 (.I(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8413__A2 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8414__A2 (.I(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__A2 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__A2 (.I(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__A2 (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8418__A2 (.I(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8419__A2 (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A2 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__A1 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__A1 (.I(\reg_file.reg_storage[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__I (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8427__A1 (.I(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__A1 (.I(\reg_file.reg_storage[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__A1 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__A1 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__A2 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__I (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__I (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__A1 (.I(\reg_file.reg_storage[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__A1 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__I (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__I (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__A2 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A2 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__I (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8454__S (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__I1 (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__S (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__A2 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__A2 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__S (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__A2 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__A2 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__I (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__S (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__S (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__I (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8470__A2 (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__A2 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__S (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__S (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__S (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8478__S (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__I (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A2 (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A2 (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__S (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A2 (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__A2 (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__A2 (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A2 (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__I (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A2 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A2 (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__I (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__A2 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A2 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A2 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A2 (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A2 (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A2 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__A1 (.I(\reg_file.reg_storage[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A1 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A1 (.I(\reg_file.reg_storage[13][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__I (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__A1 (.I(\reg_file.reg_storage[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__A1 (.I(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A1 (.I(\reg_file.reg_storage[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__A1 (.I(\reg_file.reg_storage[13][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__A1 (.I(\reg_file.reg_storage[13][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A1 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__A1 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__I (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__I (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__A1 (.I(\reg_file.reg_storage[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__I (.I(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__I (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8535__A2 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__A2 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__I (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__S (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__I1 (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__S (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__A2 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__A2 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__S (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__A2 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__A2 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8549__I (.I(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8550__S (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__S (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__I (.I(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A2 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__A2 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__S (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__S (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__S (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__S (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__I (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__A2 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__A2 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__S (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__A2 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__A2 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__A2 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__A2 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__I (.I(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__A2 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__A2 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__I (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__A2 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__A2 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__A2 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__A2 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__A2 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__A2 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__A2 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A2 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__A1 (.I(\reg_file.reg_storage[12][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__A2 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__A2 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__A1 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__A1 (.I(\reg_file.reg_storage[12][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__I (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__A1 (.I(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__A1 (.I(\reg_file.reg_storage[12][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__A1 (.I(\reg_file.reg_storage[12][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__A1 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__I (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__A1 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__A1 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__A2 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__I (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8611__I (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8612__A1 (.I(\reg_file.reg_storage[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__I (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__I (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__I (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__I (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__I (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__A1 (.I(\reg_file.reg_storage[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__A2 (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__I (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__I (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__I (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__S (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8628__I (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__S (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__I (.I(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8633__A2 (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8634__I (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8635__S (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8637__I (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__A1 (.I(\reg_file.reg_storage[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8639__A2 (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8640__I (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__I (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__S (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__I (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__S (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__I (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__I (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__A2 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__A2 (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__I (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__S (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8654__I (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__S (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8657__I (.I(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__S (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__I (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__S (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__I (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8664__I (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__A2 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8666__A2 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__S (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8670__I (.I(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8671__A2 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8672__A2 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__I (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8674__A2 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8675__A2 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8676__I (.I(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__I (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8679__A2 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8680__I (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8681__I (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8683__A2 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8685__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8686__A2 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8688__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8689__A2 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8691__A2 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__A2 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8694__A2 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8696__I (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8703__I (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8704__A2 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8706__I (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8708__A2 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__I (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8711__A2 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8713__I (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8714__A2 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8716__I (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8717__A1 (.I(\reg_file.reg_storage[8][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8719__I (.I(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__A1 (.I(\reg_file.reg_storage[8][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__A1 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__A2 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8726__A1 (.I(\reg_file.reg_storage[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__A1 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__I (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8730__I (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__I (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8732__I (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8733__A2 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8734__A2 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8735__I (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8736__I (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8737__S (.I(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__I0 (.I(\reg_file.reg_storage[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__S (.I(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8741__A2 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8742__A2 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8743__S (.I(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8745__A2 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__A2 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8747__I (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8748__S (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8750__S (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8752__I (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8753__A2 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8754__A2 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8755__S (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8757__S (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8759__S (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8761__S (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8763__I (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8764__A2 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8765__A2 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8766__S (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8768__A2 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8769__A2 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8770__A2 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8771__A2 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8772__I (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8773__A2 (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8774__A2 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8775__I (.I(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8776__A2 (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8777__A2 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__A2 (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__A2 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8780__A2 (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__A2 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8783__A2 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8784__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8785__A2 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8800__A1 (.I(\reg_file.reg_storage[11][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8802__A1 (.I(\reg_file.reg_storage[11][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8804__A1 (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8804__A2 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8808__A1 (.I(\reg_file.reg_storage[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8810__A1 (.I(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__I (.I(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8812__I (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8813__I (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8814__I (.I(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8815__A2 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8816__A2 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8817__I (.I(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8818__I (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8819__S (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8821__S (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8823__A2 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__A2 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8825__S (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8827__A2 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8828__A2 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8829__I (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8830__S (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8832__S (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8834__I (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8835__A2 (.I(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8836__A2 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8837__S (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8839__S (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8841__S (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8843__S (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8845__I (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8846__A2 (.I(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__A2 (.I(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8848__S (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8850__A2 (.I(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8851__A2 (.I(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8852__A2 (.I(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8853__A2 (.I(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8854__I (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8855__A2 (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8856__A2 (.I(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8857__I (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8858__A2 (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8859__A2 (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8860__A2 (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8861__A2 (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8862__A2 (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8863__A2 (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8864__A2 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8865__A2 (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8866__A2 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8867__A2 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8873__A2 (.I(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8876__A2 (.I(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8878__A2 (.I(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8880__A2 (.I(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8884__A1 (.I(\reg_file.reg_storage[10][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8886__A1 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8886__A2 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8887__I (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8889__I (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8890__A1 (.I(\reg_file.reg_storage[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8892__A1 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8893__I (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8894__I (.I(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8895__I (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8896__I (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8897__A2 (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8898__A2 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8899__I (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8900__I (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8901__S (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8903__I0 (.I(\reg_file.reg_storage[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8903__S (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8905__A2 (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8906__A2 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8907__S (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8909__A2 (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8910__A2 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8911__I (.I(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8912__S (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8914__S (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8916__I (.I(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8917__A2 (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8918__A2 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8919__S (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8921__S (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8923__S (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8925__S (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8927__I (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8928__A2 (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8929__A2 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8930__S (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8932__A2 (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8933__A2 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8934__A2 (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8935__A2 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8936__I (.I(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8937__A1 (.I(\reg_file.reg_storage[9][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8937__A2 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8938__A2 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8939__I (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8940__A2 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8941__A2 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8942__A2 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8943__A2 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8944__A2 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8945__A2 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8946__A2 (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8947__A2 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8948__A2 (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8949__A2 (.I(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8954__I (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8964__A1 (.I(\reg_file.reg_storage[9][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8966__A1 (.I(\reg_file.reg_storage[9][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8968__A1 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8968__A2 (.I(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8970__I (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8972__A2 (.I(_4407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8973__A1 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8973__A2 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8974__A1 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8974__A3 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8978__A2 (.I(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8979__A2 (.I(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8981__I (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8982__S (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8984__I1 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8984__S (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8986__A2 (.I(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8987__A2 (.I(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8988__S (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8990__A2 (.I(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8991__A2 (.I(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8992__I (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8993__S (.I(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8995__S (.I(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8997__I (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8998__A2 (.I(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8999__A1 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8999__A2 (.I(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9000__A2 (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9001__A2 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9002__S (.I(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9004__I0 (.I(\reg_file.reg_storage[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9004__I1 (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9004__S (.I(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9006__S (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9009__A1 (.I(\reg_file.reg_storage[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9009__A2 (.I(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9010__A2 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9011__A1 (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9011__A2 (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9012__A2 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9013__A1 (.I(\reg_file.reg_storage[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9013__A2 (.I(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9014__A2 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9015__A1 (.I(\reg_file.reg_storage[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9015__A2 (.I(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9016__A2 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9018__A2 (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9019__A2 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9020__I (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9021__A2 (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9022__A2 (.I(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9023__A2 (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9024__A2 (.I(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9025__A2 (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9026__A1 (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9026__A2 (.I(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9028__A2 (.I(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9030__A2 (.I(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9033__A1 (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9033__A2 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__I (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9036__A1 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9038__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9040__A1 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9043__A1 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9045__A1 (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9045__A2 (.I(_4407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9047__A1 (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9047__A2 (.I(_4407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9049__A1 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9049__A2 (.I(_4407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9050__A1 (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9050__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9054__A1 (.I(\reg_file.reg_storage[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9054__A2 (.I(_4457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9055__A1 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9055__A2 (.I(_4456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9056__A1 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9058__I (.I(_4460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9059__I (.I(_4461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9061__A2 (.I(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9062__A2 (.I(_4462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9064__I (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9065__S (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9067__I1 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9067__S (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9069__A2 (.I(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9070__A2 (.I(_4462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9071__S (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9073__A2 (.I(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9074__A2 (.I(_4462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9075__I (.I(_4460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9076__S (.I(_4472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9078__S (.I(_4472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9080__I (.I(_4460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9081__A2 (.I(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9082__A1 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9082__A2 (.I(_4462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9083__S (.I(_4472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9085__S (.I(_4472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9087__I1 (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9087__S (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9089__S (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9091__I (.I(_4461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9092__A2 (.I(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9093__A2 (.I(_4481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9094__I1 (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9094__S (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9096__A2 (.I(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9097__A2 (.I(_4481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9098__A2 (.I(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9099__A2 (.I(_4481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9100__I (.I(_4460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9101__A2 (.I(_4486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9102__A2 (.I(_4481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9103__I (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9104__A2 (.I(_4486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9105__A2 (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9106__A2 (.I(_4486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9107__A2 (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9108__A2 (.I(_4486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9109__A1 (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9109__A2 (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9110__A2 (.I(_4461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9111__A2 (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9112__A2 (.I(_4461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9113__A2 (.I(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9114__A2 (.I(_4457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9115__A1 (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9115__A2 (.I(_4456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9116__A2 (.I(_4457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9117__A1 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9117__A2 (.I(_4456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9119__A2 (.I(_4496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9120__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9120__A2 (.I(_4456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9122__A2 (.I(_4496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9123__A1 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9123__A2 (.I(_4498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9124__A2 (.I(_4496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9125__A1 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9125__A2 (.I(_4498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9126__A2 (.I(_4496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9127__A1 (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9127__A2 (.I(_4498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9129__A1 (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9129__A2 (.I(_4498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9131__A1 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9131__A2 (.I(_4457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9132__A1 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9132__A2 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9136__A1 (.I(\reg_file.reg_storage[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9137__A1 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9138__A1 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9140__I (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9141__I (.I(_4511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9143__A2 (.I(_4513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9144__A2 (.I(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9146__I (.I(_4515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9147__S (.I(_4516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9149__I1 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9149__S (.I(_4516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9151__A2 (.I(_4513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9152__A2 (.I(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9153__S (.I(_4516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9155__A2 (.I(_4513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9156__A2 (.I(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9157__I (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9158__S (.I(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9160__S (.I(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9162__I (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9163__A2 (.I(_4525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9164__A1 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9164__A2 (.I(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9165__S (.I(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9167__S (.I(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9169__I1 (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9169__S (.I(_4515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9171__S (.I(_4515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9173__I (.I(_4511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9174__A2 (.I(_4525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9175__A2 (.I(_4531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9176__I1 (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9176__S (.I(_4515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9178__A2 (.I(_4525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9179__A2 (.I(_4531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9180__A1 (.I(\reg_file.reg_storage[15][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9180__A2 (.I(_4525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9181__A2 (.I(_4531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9182__I (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9183__A2 (.I(_4536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9184__A2 (.I(_4531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9185__I (.I(_4516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9186__A2 (.I(_4536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9187__A2 (.I(_4538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9188__A2 (.I(_4536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9189__A2 (.I(_4538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9190__A2 (.I(_4536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9191__A1 (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9191__A2 (.I(_4538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9192__A2 (.I(_4511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9193__A2 (.I(_4538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9194__A2 (.I(_4511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9195__A2 (.I(_4513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9197__A1 (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9199__A1 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9202__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9205__A1 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9207__A1 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9209__A1 (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9211__A1 (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9213__A1 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9224__CLK (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9231__CLK (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9252__CLK (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9281__CLK (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9287__CLK (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9294__CLK (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9309__CLK (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9330__CLK (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9383__CLK (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9534__CLK (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9539__CLK (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9569__CLK (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9573__CLK (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9599__CLK (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9610__CLK (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9626__CLK (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_clk_I (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_clk_I (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_clk_I (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_clk_I (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_clk_I (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_126_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_128_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_129_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_130_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_131_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_132_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_133_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_134_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_135_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_136_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clk_I (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clk_I (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clk_I (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clk_I (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clk_I (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clk_I (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clk_I (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clk_I (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clk_I (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clk_I (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clk_I (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clk_I (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clk_I (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clk_I (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clk_I (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clk_I (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(inst[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(inst[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(inst[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(inst[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(inst[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(inst[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(inst[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(inst[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(inst[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(inst[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(inst[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(inst[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(inst[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(inst[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(inst[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(inst[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(inst[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(inst[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(inst[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(inst[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(inst[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(inst[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(inst[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(inst[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(inst[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(mem_ld_dat[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(mem_ld_dat[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(mem_ld_dat[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(mem_ld_dat[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(mem_ld_dat[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(mem_ld_dat[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(mem_ld_dat[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(inst[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(mem_ld_dat[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(mem_ld_dat[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(mem_ld_dat[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(mem_ld_dat[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(mem_ld_dat[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(mem_ld_dat[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(mem_ld_dat[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(mem_ld_dat[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(mem_ld_dat[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(mem_ld_dat[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(inst[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(mem_ld_dat[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(mem_ld_dat[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(mem_ld_dat[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(mem_ld_dat[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(mem_ld_dat[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(mem_ld_dat[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(mem_ld_dat[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(mem_ld_dat[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(mem_ld_dat[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(mem_ld_dat[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(inst[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(mem_ld_dat[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(mem_ld_dat[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(mem_ld_dat[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(mem_ld_dat[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(mem_ld_dat[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(pc[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(pc[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(pc[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(pc[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(pc[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(inst[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(pc[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(pc[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(pc[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(pc[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(pc[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(pc[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(pc[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(pc[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(pc[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(pc[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(inst[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(pc[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(pc[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(pc[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(pc[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(pc[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(pc[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(pc[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(pc[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(pc[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(pc[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(inst[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(pc[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(pc[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(pc[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(pc[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(pc[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(pc[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(pc[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(inst[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_load_slew1_I (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output102_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output103_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output104_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output108_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output109_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output124_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output128_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output129_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output134_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output135_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output136_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output137_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output138_I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output139_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output140_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output141_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output142_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output143_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output144_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output145_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output149_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output152_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output153_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output154_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output155_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output156_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output157_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output158_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output159_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output160_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output161_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output162_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output163_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output164_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output166_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output175_I (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output180_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output185_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output186_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output188_I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output189_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output191_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output194_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output195_I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer16_I (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer17_I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer18_I (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer19_I (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer20_I (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer22_I (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer23_I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer25_I (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer27_I (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer28_I (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer30_I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer8_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer9_I (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_438 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4554_ (.I(net13),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4555_ (.I(_0480_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4556_ (.I(net14),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4557_ (.I(_0482_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4558_ (.A1(_0481_),
    .A2(_0483_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4559_ (.I(net15),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4560_ (.A1(_0485_),
    .A2(net16),
    .A3(net17),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4561_ (.A1(_0484_),
    .A2(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4562_ (.I(_0487_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4563_ (.I(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4564_ (.I(_0489_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4565_ (.I(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4566_ (.I(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4567_ (.I(_0492_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4568_ (.I(_0493_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4569_ (.I(net13),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4570_ (.I(_0495_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4571_ (.I(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4572_ (.I(net14),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4573_ (.I(_0498_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4574_ (.I(_0499_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4575_ (.I0(\reg_file.reg_storage[4][0] ),
    .I1(\reg_file.reg_storage[5][0] ),
    .I2(\reg_file.reg_storage[6][0] ),
    .I3(\reg_file.reg_storage[7][0] ),
    .S0(_0497_),
    .S1(_0500_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4576_ (.I(net13),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4577_ (.I(_0502_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4578_ (.I0(\reg_file.reg_storage[2][0] ),
    .I1(\reg_file.reg_storage[3][0] ),
    .S(_0503_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4579_ (.I0(\reg_file.reg_storage[1][0] ),
    .I1(_0504_),
    .S(_0500_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4580_ (.I0(\reg_file.reg_storage[12][0] ),
    .I1(\reg_file.reg_storage[13][0] ),
    .I2(\reg_file.reg_storage[14][0] ),
    .I3(\reg_file.reg_storage[15][0] ),
    .S0(_0497_),
    .S1(_0500_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4581_ (.I0(\reg_file.reg_storage[8][0] ),
    .I1(\reg_file.reg_storage[9][0] ),
    .I2(\reg_file.reg_storage[10][0] ),
    .I3(\reg_file.reg_storage[11][0] ),
    .S0(_0497_),
    .S1(_0500_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4582_ (.I(net15),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4583_ (.I(_0508_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4584_ (.I(net16),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4585_ (.I0(_0501_),
    .I1(_0505_),
    .I2(_0506_),
    .I3(_0507_),
    .S0(_0509_),
    .S1(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4586_ (.A1(_0494_),
    .A2(net231),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4587_ (.I(_0512_),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4588_ (.I(_0495_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4589_ (.I(_0482_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4590_ (.I0(\reg_file.reg_storage[8][1] ),
    .I1(\reg_file.reg_storage[9][1] ),
    .I2(\reg_file.reg_storage[10][1] ),
    .I3(\reg_file.reg_storage[11][1] ),
    .S0(_0513_),
    .S1(_0514_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4591_ (.I0(\reg_file.reg_storage[2][1] ),
    .I1(\reg_file.reg_storage[3][1] ),
    .S(_0502_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4592_ (.I0(\reg_file.reg_storage[1][1] ),
    .I1(_0516_),
    .S(_0514_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4593_ (.I(_0482_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4594_ (.I0(\reg_file.reg_storage[12][1] ),
    .I1(\reg_file.reg_storage[13][1] ),
    .I2(\reg_file.reg_storage[14][1] ),
    .I3(\reg_file.reg_storage[15][1] ),
    .S0(_0480_),
    .S1(_0518_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4595_ (.I0(\reg_file.reg_storage[4][1] ),
    .I1(\reg_file.reg_storage[5][1] ),
    .I2(\reg_file.reg_storage[6][1] ),
    .I3(\reg_file.reg_storage[7][1] ),
    .S0(_0480_),
    .S1(_0518_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4596_ (.I(net16),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4597_ (.I0(_0515_),
    .I1(_0517_),
    .I2(_0519_),
    .I3(_0520_),
    .S0(_0521_),
    .S1(_0485_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4598_ (.A1(_0487_),
    .A2(_0522_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4599_ (.I(_0523_),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4600_ (.I0(\reg_file.reg_storage[4][2] ),
    .I1(\reg_file.reg_storage[5][2] ),
    .I2(\reg_file.reg_storage[6][2] ),
    .I3(\reg_file.reg_storage[7][2] ),
    .S0(_0513_),
    .S1(_0514_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4601_ (.I0(\reg_file.reg_storage[2][2] ),
    .I1(\reg_file.reg_storage[3][2] ),
    .S(_0502_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4602_ (.I0(\reg_file.reg_storage[1][2] ),
    .I1(_0525_),
    .S(_0499_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4603_ (.I0(_0524_),
    .I1(_0526_),
    .S(_0509_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4604_ (.I(_0521_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4605_ (.I0(\reg_file.reg_storage[12][2] ),
    .I1(\reg_file.reg_storage[13][2] ),
    .I2(\reg_file.reg_storage[14][2] ),
    .I3(\reg_file.reg_storage[15][2] ),
    .S0(_0495_),
    .S1(net229),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4606_ (.I0(\reg_file.reg_storage[8][2] ),
    .I1(\reg_file.reg_storage[9][2] ),
    .I2(\reg_file.reg_storage[10][2] ),
    .I3(\reg_file.reg_storage[11][2] ),
    .S0(_0495_),
    .S1(net229),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4607_ (.I0(_0529_),
    .I1(_0530_),
    .S(_0508_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4608_ (.A1(_0528_),
    .A2(_0531_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4609_ (.A1(_0510_),
    .A2(_0527_),
    .B(_0532_),
    .C(_0487_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _4610_ (.I(_0533_),
    .ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4611_ (.I(_0513_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4612_ (.I(_0482_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4613_ (.I0(\reg_file.reg_storage[8][3] ),
    .I1(\reg_file.reg_storage[9][3] ),
    .I2(\reg_file.reg_storage[10][3] ),
    .I3(\reg_file.reg_storage[11][3] ),
    .S0(_0534_),
    .S1(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4614_ (.I0(\reg_file.reg_storage[2][3] ),
    .I1(\reg_file.reg_storage[3][3] ),
    .S(_0496_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4615_ (.I0(\reg_file.reg_storage[1][3] ),
    .I1(_0537_),
    .S(_0535_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4616_ (.I(_0498_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4617_ (.I0(\reg_file.reg_storage[12][3] ),
    .I1(\reg_file.reg_storage[13][3] ),
    .I2(\reg_file.reg_storage[14][3] ),
    .I3(\reg_file.reg_storage[15][3] ),
    .S0(_0481_),
    .S1(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4618_ (.I0(\reg_file.reg_storage[4][3] ),
    .I1(\reg_file.reg_storage[5][3] ),
    .I2(\reg_file.reg_storage[6][3] ),
    .I3(\reg_file.reg_storage[7][3] ),
    .S0(_0481_),
    .S1(_0535_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4619_ (.I(_0521_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4620_ (.I(_0485_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4621_ (.I0(_0536_),
    .I1(_0538_),
    .I2(_0540_),
    .I3(_0541_),
    .S0(_0542_),
    .S1(_0543_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4622_ (.A1(_0488_),
    .A2(_0544_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4623_ (.I(_0545_),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4624_ (.I0(\reg_file.reg_storage[8][4] ),
    .I1(\reg_file.reg_storage[9][4] ),
    .I2(\reg_file.reg_storage[10][4] ),
    .I3(\reg_file.reg_storage[11][4] ),
    .S0(_0496_),
    .S1(_0499_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4625_ (.I0(\reg_file.reg_storage[2][4] ),
    .I1(\reg_file.reg_storage[3][4] ),
    .S(_0502_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4626_ (.I0(\reg_file.reg_storage[1][4] ),
    .I1(_0547_),
    .S(_0499_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4627_ (.I0(_0546_),
    .I1(_0548_),
    .S(_0528_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4628_ (.I0(\reg_file.reg_storage[4][4] ),
    .I1(\reg_file.reg_storage[5][4] ),
    .I2(\reg_file.reg_storage[6][4] ),
    .I3(\reg_file.reg_storage[7][4] ),
    .S0(_0480_),
    .S1(_0518_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4629_ (.A1(_0510_),
    .A2(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4630_ (.I0(\reg_file.reg_storage[12][4] ),
    .I1(\reg_file.reg_storage[13][4] ),
    .I2(\reg_file.reg_storage[14][4] ),
    .I3(\reg_file.reg_storage[15][4] ),
    .S0(_0513_),
    .S1(_0514_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4631_ (.A1(_0528_),
    .A2(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4632_ (.A1(_0551_),
    .A2(_0553_),
    .B(_0543_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4633_ (.A1(_0543_),
    .A2(_0549_),
    .B(_0554_),
    .C(_0487_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _4634_ (.I(_0555_),
    .ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4635_ (.I(_0496_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4636_ (.I(_0483_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4637_ (.I0(\reg_file.reg_storage[8][5] ),
    .I1(\reg_file.reg_storage[9][5] ),
    .I2(\reg_file.reg_storage[10][5] ),
    .I3(\reg_file.reg_storage[11][5] ),
    .S0(_0556_),
    .S1(_0557_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4638_ (.I0(\reg_file.reg_storage[2][5] ),
    .I1(\reg_file.reg_storage[3][5] ),
    .S(_0503_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4639_ (.I0(\reg_file.reg_storage[1][5] ),
    .I1(_0559_),
    .S(_0557_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4640_ (.I0(\reg_file.reg_storage[12][5] ),
    .I1(\reg_file.reg_storage[13][5] ),
    .I2(\reg_file.reg_storage[14][5] ),
    .I3(\reg_file.reg_storage[15][5] ),
    .S0(_0556_),
    .S1(_0557_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4641_ (.I0(\reg_file.reg_storage[4][5] ),
    .I1(\reg_file.reg_storage[5][5] ),
    .I2(\reg_file.reg_storage[6][5] ),
    .I3(\reg_file.reg_storage[7][5] ),
    .S0(_0556_),
    .S1(_0557_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4642_ (.I(_0485_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4643_ (.I0(_0558_),
    .I1(_0560_),
    .I2(_0561_),
    .I3(_0562_),
    .S0(_0542_),
    .S1(_0563_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4644_ (.A1(_0494_),
    .A2(net221),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4645_ (.I(_0565_),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4646_ (.I(_0503_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4647_ (.I(_0483_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4648_ (.I0(\reg_file.reg_storage[8][6] ),
    .I1(\reg_file.reg_storage[9][6] ),
    .I2(\reg_file.reg_storage[10][6] ),
    .I3(\reg_file.reg_storage[11][6] ),
    .S0(_0566_),
    .S1(_0567_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4649_ (.I0(\reg_file.reg_storage[2][6] ),
    .I1(\reg_file.reg_storage[3][6] ),
    .S(_0534_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4650_ (.I(net14),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4651_ (.I0(\reg_file.reg_storage[1][6] ),
    .I1(_0569_),
    .S(_0570_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4652_ (.I(_0503_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4653_ (.I0(\reg_file.reg_storage[12][6] ),
    .I1(\reg_file.reg_storage[13][6] ),
    .I2(\reg_file.reg_storage[14][6] ),
    .I3(\reg_file.reg_storage[15][6] ),
    .S0(_0572_),
    .S1(_0570_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4654_ (.I0(\reg_file.reg_storage[4][6] ),
    .I1(\reg_file.reg_storage[5][6] ),
    .I2(\reg_file.reg_storage[6][6] ),
    .I3(\reg_file.reg_storage[7][6] ),
    .S0(_0572_),
    .S1(_0570_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4655_ (.I0(_0568_),
    .I1(_0571_),
    .I2(_0573_),
    .I3(_0574_),
    .S0(_0542_),
    .S1(_0563_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4656_ (.A1(_0494_),
    .A2(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4657_ (.I(_0576_),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4658_ (.I(_0481_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4659_ (.I(_0539_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4660_ (.I0(\reg_file.reg_storage[8][7] ),
    .I1(\reg_file.reg_storage[9][7] ),
    .I2(\reg_file.reg_storage[10][7] ),
    .I3(\reg_file.reg_storage[11][7] ),
    .S0(_0577_),
    .S1(_0578_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4661_ (.I0(\reg_file.reg_storage[2][7] ),
    .I1(\reg_file.reg_storage[3][7] ),
    .S(_0497_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4662_ (.I0(\reg_file.reg_storage[1][7] ),
    .I1(_0580_),
    .S(_0578_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4663_ (.I0(\reg_file.reg_storage[12][7] ),
    .I1(\reg_file.reg_storage[13][7] ),
    .I2(\reg_file.reg_storage[14][7] ),
    .I3(\reg_file.reg_storage[15][7] ),
    .S0(_0566_),
    .S1(_0567_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4664_ (.I0(\reg_file.reg_storage[4][7] ),
    .I1(\reg_file.reg_storage[5][7] ),
    .I2(\reg_file.reg_storage[6][7] ),
    .I3(\reg_file.reg_storage[7][7] ),
    .S0(_0566_),
    .S1(_0567_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4665_ (.I0(_0579_),
    .I1(_0581_),
    .I2(_0582_),
    .I3(_0583_),
    .S0(_0542_),
    .S1(_0563_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4666_ (.A1(_0493_),
    .A2(_0584_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4667_ (.I(_0585_),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4668_ (.I(net27),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4669_ (.I(_0586_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4670_ (.I(net28),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4671_ (.I(net29),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4672_ (.A1(net12),
    .A2(net1),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _4673_ (.A1(net26),
    .A2(net23),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4674_ (.A1(_0588_),
    .A2(_0589_),
    .A3(_0590_),
    .A4(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4675_ (.I(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4676_ (.A1(_0587_),
    .A2(_0593_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4677_ (.I(_0594_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4678_ (.I(_0595_),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4679_ (.I(net28),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4680_ (.I(_0596_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4681_ (.I(net27),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4682_ (.I(_0598_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4683_ (.I(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4684_ (.I(net29),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4685_ (.I(_0590_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4686_ (.I(_0591_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4687_ (.A1(_0601_),
    .A2(_0602_),
    .A3(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4688_ (.I(_0604_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4689_ (.A1(_0597_),
    .A2(_0600_),
    .A3(_0605_),
    .ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4690_ (.I(net65),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4691_ (.I(net26),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4692_ (.I(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4693_ (.I(_0588_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _4694_ (.A1(net12),
    .A2(net1),
    .A3(net23),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4695_ (.I(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4696_ (.A1(_0609_),
    .A2(_0587_),
    .A3(_0601_),
    .A4(_0611_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4697_ (.I(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4698_ (.I(_0589_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4699_ (.A1(_0614_),
    .A2(_0602_),
    .A3(_0603_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4700_ (.I(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4701_ (.A1(_0609_),
    .A2(_0587_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4702_ (.I(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _4703_ (.A1(_0608_),
    .A2(_0613_),
    .B1(_0616_),
    .B2(_0618_),
    .C(_0605_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4704_ (.I(_0619_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4705_ (.I(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4706_ (.A1(_0606_),
    .A2(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4707_ (.I(net8),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4708_ (.I(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4709_ (.I(net9),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4710_ (.I(net11),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4711_ (.I(net7),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4712_ (.I(_0627_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4713_ (.A1(net10),
    .A2(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4714_ (.A1(_0624_),
    .A2(_0625_),
    .A3(_0626_),
    .A4(_0629_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4715_ (.I(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4716_ (.I(net7),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4717_ (.I(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4718_ (.I(net8),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4719_ (.I(_0634_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4720_ (.I0(\reg_file.reg_storage[4][0] ),
    .I1(\reg_file.reg_storage[5][0] ),
    .I2(\reg_file.reg_storage[6][0] ),
    .I3(\reg_file.reg_storage[7][0] ),
    .S0(_0633_),
    .S1(_0635_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4721_ (.I(_0627_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4722_ (.I(_0637_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4723_ (.I0(\reg_file.reg_storage[2][0] ),
    .I1(\reg_file.reg_storage[3][0] ),
    .S(_0638_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4724_ (.I(net8),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4725_ (.I(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4726_ (.I(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4727_ (.I0(\reg_file.reg_storage[1][0] ),
    .I1(_0639_),
    .S(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4728_ (.I(_0632_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4729_ (.I(_0634_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4730_ (.I0(\reg_file.reg_storage[12][0] ),
    .I1(\reg_file.reg_storage[13][0] ),
    .I2(\reg_file.reg_storage[14][0] ),
    .I3(\reg_file.reg_storage[15][0] ),
    .S0(_0644_),
    .S1(_0645_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4731_ (.I0(\reg_file.reg_storage[8][0] ),
    .I1(\reg_file.reg_storage[9][0] ),
    .I2(\reg_file.reg_storage[10][0] ),
    .I3(\reg_file.reg_storage[11][0] ),
    .S0(_0644_),
    .S1(_0645_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4732_ (.I(_0625_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4733_ (.I(net10),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4734_ (.I0(_0636_),
    .I1(_0643_),
    .I2(_0646_),
    .I3(_0647_),
    .S0(_0648_),
    .S1(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4735_ (.A1(_0620_),
    .A2(_0631_),
    .A3(_0650_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4736_ (.A1(_0609_),
    .A2(_0604_),
    .B1(_0612_),
    .B2(_0607_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4737_ (.A1(_0598_),
    .A2(_0589_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _4738_ (.A1(_0607_),
    .A2(_0597_),
    .A3(_0611_),
    .A4(_0653_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4739_ (.A1(_0588_),
    .A2(_0598_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4740_ (.A1(_0614_),
    .A2(_0602_),
    .A3(_0603_),
    .A4(_0655_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4741_ (.A1(_0654_),
    .A2(_0656_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4742_ (.I(_0556_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4743_ (.I(_0658_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4744_ (.A1(_0652_),
    .A2(_0657_),
    .B(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4745_ (.A1(_0601_),
    .A2(_0590_),
    .A3(_0591_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _4746_ (.A1(_0588_),
    .A2(_0586_),
    .A3(_0601_),
    .A4(net230),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _4747_ (.I(_0607_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4748_ (.A1(net26),
    .A2(_0589_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _4749_ (.A1(_0596_),
    .A2(_0598_),
    .A3(_0610_),
    .A4(_0664_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4750_ (.A1(_0586_),
    .A2(_0661_),
    .B1(_0662_),
    .B2(_0663_),
    .C(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4751_ (.A1(_0599_),
    .A2(_0593_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4752_ (.A1(_0666_),
    .A2(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4753_ (.I(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4754_ (.I(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4755_ (.I(_0670_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4756_ (.I(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4757_ (.I(_0666_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4758_ (.I(_0667_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4759_ (.A1(_0489_),
    .A2(_0511_),
    .A3(_0673_),
    .A4(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _4760_ (.A1(_0622_),
    .A2(_0651_),
    .B1(_0660_),
    .B2(_0672_),
    .C(net216),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4761_ (.I(_0676_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4762_ (.A1(_0622_),
    .A2(_0651_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4763_ (.A1(_0666_),
    .A2(_0667_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4764_ (.I(_0679_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4765_ (.A1(_0663_),
    .A2(_0662_),
    .B(_0593_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4766_ (.I(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4767_ (.A1(_0654_),
    .A2(net215),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4768_ (.I(_0683_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4769_ (.I(_0572_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4770_ (.I(_0685_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4771_ (.I(_0686_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _4772_ (.I(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4773_ (.A1(_0682_),
    .A2(_0684_),
    .B(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4774_ (.I(_0488_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4775_ (.I(_0673_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4776_ (.I(_0674_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4777_ (.A1(_0690_),
    .A2(_0511_),
    .A3(_0691_),
    .A4(_0692_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4778_ (.A1(_0680_),
    .A2(_0689_),
    .B(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4779_ (.I(_0694_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4780_ (.A1(_0678_),
    .A2(_0695_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4781_ (.A1(_0677_),
    .A2(_0696_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4782_ (.A1(_0597_),
    .A2(_0599_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4783_ (.A1(_0614_),
    .A2(_0602_),
    .A3(_0603_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4784_ (.A1(_0698_),
    .A2(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4785_ (.I(_0700_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4786_ (.A1(net6),
    .A2(_0701_),
    .A3(_0691_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4787_ (.I(_0702_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4788_ (.I(_0703_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _4789_ (.I(net4),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4790_ (.A1(_0617_),
    .A2(_0615_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4791_ (.A1(_0597_),
    .A2(_0599_),
    .A3(_0611_),
    .A4(_0664_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _4792_ (.A1(_0600_),
    .A2(_0605_),
    .B1(_0613_),
    .B2(_0608_),
    .C(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4793_ (.I(_0698_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4794_ (.I(_0699_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4795_ (.A1(net5),
    .A2(_0709_),
    .A3(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4796_ (.I(net6),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4797_ (.A1(_0705_),
    .A2(_0706_),
    .A3(_0708_),
    .B1(_0711_),
    .B2(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4798_ (.I(net5),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4799_ (.I(_0673_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4800_ (.I(_0706_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4801_ (.A1(_0714_),
    .A2(_0715_),
    .B(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4802_ (.I(_0717_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4803_ (.A1(_0713_),
    .A2(_0718_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4804_ (.A1(_0704_),
    .A2(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4805_ (.I(_0713_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _4806_ (.I(net24),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4807_ (.A1(_0712_),
    .A2(_0709_),
    .A3(_0710_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _4808_ (.A1(_0722_),
    .A2(_0716_),
    .A3(_0708_),
    .B(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4809_ (.A1(_0703_),
    .A2(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4810_ (.A1(_0721_),
    .A2(_0718_),
    .A3(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4811_ (.I(net5),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4812_ (.I(_0700_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4813_ (.A1(_0727_),
    .A2(_0708_),
    .B(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4814_ (.A1(_0713_),
    .A2(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4815_ (.I(_0730_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4816_ (.A1(_0704_),
    .A2(_0731_),
    .B(_0724_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4817_ (.A1(_0720_),
    .A2(_0726_),
    .A3(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4818_ (.I(_0668_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4819_ (.I(_0734_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4820_ (.I(_0735_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4821_ (.I(net3),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4822_ (.A1(_0592_),
    .A2(_0662_),
    .A3(_0654_),
    .A4(_0656_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4823_ (.I(_0738_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4824_ (.I(net17),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4825_ (.A1(_0737_),
    .A2(_0728_),
    .B1(_0739_),
    .B2(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4826_ (.A1(_0555_),
    .A2(_0671_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4827_ (.A1(_0736_),
    .A2(_0741_),
    .B(_0742_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4828_ (.I(_0743_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4829_ (.I(_0744_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4830_ (.I(_0662_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4831_ (.A1(_0663_),
    .A2(_0746_),
    .B1(_0710_),
    .B2(_0709_),
    .C(_0661_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4832_ (.I(_0747_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4833_ (.I(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4834_ (.I(_0749_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4835_ (.A1(net77),
    .A2(_0750_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4836_ (.A1(_0747_),
    .A2(_0630_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4837_ (.I(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4838_ (.I(_0753_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4839_ (.I(_0627_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4840_ (.I(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4841_ (.I(_0756_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4842_ (.I(_0757_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4843_ (.I(_0640_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4844_ (.I(_0759_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4845_ (.I(_0760_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4846_ (.I0(\reg_file.reg_storage[4][20] ),
    .I1(\reg_file.reg_storage[5][20] ),
    .I2(\reg_file.reg_storage[6][20] ),
    .I3(\reg_file.reg_storage[7][20] ),
    .S0(_0758_),
    .S1(_0761_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4847_ (.I(_0623_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4848_ (.I(_0763_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4849_ (.I(_0764_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4850_ (.I(\reg_file.reg_storage[1][20] ),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4851_ (.I(_0756_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4852_ (.I(_0767_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4853_ (.A1(_0768_),
    .A2(\reg_file.reg_storage[3][20] ),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4854_ (.I(_0627_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4855_ (.I(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4856_ (.I(_0771_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4857_ (.I(_0772_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4858_ (.I(_0763_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4859_ (.I(_0774_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4860_ (.A1(_0773_),
    .A2(\reg_file.reg_storage[2][20] ),
    .B(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4861_ (.A1(_0765_),
    .A2(_0766_),
    .B1(_0769_),
    .B2(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4862_ (.I(_0632_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4863_ (.I(_0778_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4864_ (.I(_0779_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4865_ (.I(_0760_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4866_ (.I0(\reg_file.reg_storage[12][20] ),
    .I1(\reg_file.reg_storage[13][20] ),
    .I2(\reg_file.reg_storage[14][20] ),
    .I3(\reg_file.reg_storage[15][20] ),
    .S0(_0780_),
    .S1(_0781_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4867_ (.I0(\reg_file.reg_storage[8][20] ),
    .I1(\reg_file.reg_storage[9][20] ),
    .I2(\reg_file.reg_storage[10][20] ),
    .I3(\reg_file.reg_storage[11][20] ),
    .S0(_0758_),
    .S1(_0781_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4868_ (.I(_0625_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4869_ (.I(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4870_ (.I(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4871_ (.I(_0649_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4872_ (.I(_0787_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4873_ (.I0(_0762_),
    .I1(_0777_),
    .I2(_0782_),
    .I3(_0783_),
    .S0(_0786_),
    .S1(_0788_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4874_ (.A1(_0754_),
    .A2(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4875_ (.A1(_0751_),
    .A2(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4876_ (.I(_0668_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4877_ (.A1(_0792_),
    .A2(_0660_),
    .B(_0675_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4878_ (.I(_0793_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4879_ (.I(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4880_ (.I(_0795_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4881_ (.A1(_0791_),
    .A2(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4882_ (.I(_0748_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4883_ (.A1(net78),
    .A2(_0798_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4884_ (.I(_0753_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4885_ (.I(_0638_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4886_ (.I(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4887_ (.I(_0640_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4888_ (.I(_0803_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4889_ (.I0(\reg_file.reg_storage[4][21] ),
    .I1(\reg_file.reg_storage[5][21] ),
    .I2(\reg_file.reg_storage[6][21] ),
    .I3(\reg_file.reg_storage[7][21] ),
    .S0(_0802_),
    .S1(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4890_ (.I(_0624_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4891_ (.I(_0806_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4892_ (.I(\reg_file.reg_storage[1][21] ),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4893_ (.I(_0755_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4894_ (.I(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4895_ (.I(_0810_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4896_ (.A1(_0811_),
    .A2(\reg_file.reg_storage[3][21] ),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4897_ (.I(_0771_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4898_ (.I(_0763_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4899_ (.A1(_0813_),
    .A2(\reg_file.reg_storage[2][21] ),
    .B(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4900_ (.A1(_0807_),
    .A2(_0808_),
    .B1(_0812_),
    .B2(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4901_ (.I(_0801_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4902_ (.I(_0635_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4903_ (.I0(\reg_file.reg_storage[12][21] ),
    .I1(\reg_file.reg_storage[13][21] ),
    .I2(\reg_file.reg_storage[14][21] ),
    .I3(\reg_file.reg_storage[15][21] ),
    .S0(_0817_),
    .S1(_0818_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4904_ (.I0(\reg_file.reg_storage[8][21] ),
    .I1(\reg_file.reg_storage[9][21] ),
    .I2(\reg_file.reg_storage[10][21] ),
    .I3(\reg_file.reg_storage[11][21] ),
    .S0(_0817_),
    .S1(_0818_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4905_ (.I(_0648_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4906_ (.I(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4907_ (.I(net10),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4908_ (.I(_0823_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4909_ (.I(_0824_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4910_ (.I0(_0805_),
    .I1(_0816_),
    .I2(_0819_),
    .I3(_0820_),
    .S0(_0822_),
    .S1(_0825_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4911_ (.A1(_0800_),
    .A2(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4912_ (.A1(_0799_),
    .A2(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4913_ (.I(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4914_ (.I(_0695_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4915_ (.I(_0830_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4916_ (.A1(_0829_),
    .A2(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4917_ (.A1(_0797_),
    .A2(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4918_ (.A1(_0619_),
    .A2(_0631_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4919_ (.I(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4920_ (.I(_0641_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4921_ (.I(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4922_ (.I0(\reg_file.reg_storage[4][22] ),
    .I1(\reg_file.reg_storage[5][22] ),
    .I2(\reg_file.reg_storage[6][22] ),
    .I3(\reg_file.reg_storage[7][22] ),
    .S0(_0757_),
    .S1(_0837_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4923_ (.I(_0633_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4924_ (.I0(\reg_file.reg_storage[2][22] ),
    .I1(\reg_file.reg_storage[3][22] ),
    .S(_0839_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4925_ (.I0(\reg_file.reg_storage[1][22] ),
    .I1(_0840_),
    .S(_0837_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4926_ (.I(_0635_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4927_ (.I0(\reg_file.reg_storage[12][22] ),
    .I1(\reg_file.reg_storage[13][22] ),
    .I2(\reg_file.reg_storage[14][22] ),
    .I3(\reg_file.reg_storage[15][22] ),
    .S0(_0757_),
    .S1(_0842_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4928_ (.I0(\reg_file.reg_storage[8][22] ),
    .I1(\reg_file.reg_storage[9][22] ),
    .I2(\reg_file.reg_storage[10][22] ),
    .I3(\reg_file.reg_storage[11][22] ),
    .S0(_0757_),
    .S1(_0842_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4929_ (.I0(_0838_),
    .I1(_0841_),
    .I2(_0843_),
    .I3(_0844_),
    .S0(_0785_),
    .S1(_0825_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4930_ (.I(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4931_ (.A1(net79),
    .A2(_0798_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4932_ (.A1(_0835_),
    .A2(_0846_),
    .B(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4933_ (.I(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4934_ (.I(_0695_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4935_ (.I(_0850_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4936_ (.I(_0749_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4937_ (.A1(net80),
    .A2(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4938_ (.I(_0638_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4939_ (.I(_0854_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4940_ (.I(_0641_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4941_ (.I(_0856_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4942_ (.I0(\reg_file.reg_storage[4][23] ),
    .I1(\reg_file.reg_storage[5][23] ),
    .I2(\reg_file.reg_storage[6][23] ),
    .I3(\reg_file.reg_storage[7][23] ),
    .S0(_0855_),
    .S1(_0857_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4943_ (.I(\reg_file.reg_storage[1][23] ),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4944_ (.I(_0756_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4945_ (.I(_0860_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4946_ (.A1(_0861_),
    .A2(\reg_file.reg_storage[3][23] ),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4947_ (.I(_0771_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4948_ (.A1(_0863_),
    .A2(\reg_file.reg_storage[2][23] ),
    .B(_0764_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4949_ (.A1(_0775_),
    .A2(_0859_),
    .B1(_0862_),
    .B2(_0864_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4950_ (.I(_0854_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4951_ (.I(_0856_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4952_ (.I0(\reg_file.reg_storage[12][23] ),
    .I1(\reg_file.reg_storage[13][23] ),
    .I2(\reg_file.reg_storage[14][23] ),
    .I3(\reg_file.reg_storage[15][23] ),
    .S0(_0866_),
    .S1(_0867_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4953_ (.I0(\reg_file.reg_storage[8][23] ),
    .I1(\reg_file.reg_storage[9][23] ),
    .I2(\reg_file.reg_storage[10][23] ),
    .I3(\reg_file.reg_storage[11][23] ),
    .S0(_0866_),
    .S1(_0867_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4954_ (.I(_0821_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4955_ (.I(_0824_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4956_ (.I0(_0858_),
    .I1(_0865_),
    .I2(_0868_),
    .I3(_0869_),
    .S0(_0870_),
    .S1(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4957_ (.A1(_0800_),
    .A2(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4958_ (.A1(_0853_),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4959_ (.I(_0830_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4960_ (.A1(_0874_),
    .A2(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4961_ (.A1(_0849_),
    .A2(_0851_),
    .B(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4962_ (.I(_0483_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4963_ (.I(_0878_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _4964_ (.I(net31),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4965_ (.A1(_0880_),
    .A2(_0618_),
    .A3(_0616_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4966_ (.I0(_0879_),
    .I1(_0881_),
    .S(_0739_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4967_ (.I0(net145),
    .I1(_0882_),
    .S(_0679_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4968_ (.I(net226),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4969_ (.I(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4970_ (.I(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4971_ (.I0(_0833_),
    .I1(_0877_),
    .S(_0886_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4972_ (.I(_0748_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4973_ (.I(_0888_),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4974_ (.I(_0753_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4975_ (.I(_0890_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4976_ (.I(_0756_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4977_ (.I(_0842_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4978_ (.I0(\reg_file.reg_storage[4][17] ),
    .I1(\reg_file.reg_storage[5][17] ),
    .I2(\reg_file.reg_storage[6][17] ),
    .I3(\reg_file.reg_storage[7][17] ),
    .S0(_0892_),
    .S1(_0893_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4979_ (.I(\reg_file.reg_storage[1][17] ),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4980_ (.I(_0854_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4981_ (.I(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4982_ (.A1(_0897_),
    .A2(\reg_file.reg_storage[3][17] ),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4983_ (.I(_0774_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4984_ (.A1(_0773_),
    .A2(\reg_file.reg_storage[2][17] ),
    .B(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4985_ (.A1(_0765_),
    .A2(_0895_),
    .B1(_0898_),
    .B2(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4986_ (.I(_0759_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4987_ (.I(_0902_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4988_ (.I0(\reg_file.reg_storage[12][17] ),
    .I1(\reg_file.reg_storage[13][17] ),
    .I2(\reg_file.reg_storage[14][17] ),
    .I3(\reg_file.reg_storage[15][17] ),
    .S0(_0861_),
    .S1(_0903_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4989_ (.I0(\reg_file.reg_storage[8][17] ),
    .I1(\reg_file.reg_storage[9][17] ),
    .I2(\reg_file.reg_storage[10][17] ),
    .I3(\reg_file.reg_storage[11][17] ),
    .S0(_0861_),
    .S1(_0893_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4990_ (.I(_0784_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4991_ (.I0(_0894_),
    .I1(_0901_),
    .I2(_0904_),
    .I3(_0905_),
    .S0(_0906_),
    .S1(_0788_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4992_ (.A1(net73),
    .A2(_0889_),
    .B1(_0891_),
    .B2(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4993_ (.I(_0794_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4994_ (.I(_0909_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4995_ (.I(net72),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4996_ (.I(_0620_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4997_ (.I(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _4998_ (.I(_0823_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4999_ (.I(\reg_file.reg_storage[2][16] ),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5000_ (.A1(_0892_),
    .A2(\reg_file.reg_storage[3][16] ),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5001_ (.A1(_0897_),
    .A2(_0915_),
    .B(_0916_),
    .C(_0893_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5002_ (.A1(_0893_),
    .A2(\reg_file.reg_storage[1][16] ),
    .B(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5003_ (.I(_0755_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5004_ (.I(_0919_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5005_ (.I(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5006_ (.I(_0836_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5007_ (.I0(\reg_file.reg_storage[4][16] ),
    .I1(\reg_file.reg_storage[5][16] ),
    .I2(\reg_file.reg_storage[6][16] ),
    .I3(\reg_file.reg_storage[7][16] ),
    .S0(_0921_),
    .S1(_0922_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5008_ (.A1(_0906_),
    .A2(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5009_ (.A1(_0906_),
    .A2(_0918_),
    .B(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5010_ (.I0(\reg_file.reg_storage[8][16] ),
    .I1(\reg_file.reg_storage[9][16] ),
    .I2(\reg_file.reg_storage[10][16] ),
    .I3(\reg_file.reg_storage[11][16] ),
    .S0(_0780_),
    .S1(_0781_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5011_ (.A1(net9),
    .A2(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5012_ (.I0(\reg_file.reg_storage[12][16] ),
    .I1(\reg_file.reg_storage[13][16] ),
    .I2(\reg_file.reg_storage[14][16] ),
    .I3(\reg_file.reg_storage[15][16] ),
    .S0(_0780_),
    .S1(_0781_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5013_ (.I(_0787_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5014_ (.A1(_0906_),
    .A2(_0928_),
    .B(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5015_ (.A1(_0927_),
    .A2(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5016_ (.A1(_0914_),
    .A2(_0925_),
    .B(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5017_ (.A1(_0911_),
    .A2(_0913_),
    .B1(_0835_),
    .B2(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5018_ (.A1(_0933_),
    .A2(_0796_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5019_ (.A1(_0908_),
    .A2(_0910_),
    .B(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5020_ (.I(net74),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5021_ (.I(_0621_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5022_ (.I(_0631_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5023_ (.I0(\reg_file.reg_storage[4][18] ),
    .I1(\reg_file.reg_storage[5][18] ),
    .I2(\reg_file.reg_storage[6][18] ),
    .I3(\reg_file.reg_storage[7][18] ),
    .S0(_0810_),
    .S1(_0842_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5024_ (.I(_0628_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5025_ (.I0(\reg_file.reg_storage[2][18] ),
    .I1(\reg_file.reg_storage[3][18] ),
    .S(_0940_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5026_ (.I(_0856_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5027_ (.I0(\reg_file.reg_storage[1][18] ),
    .I1(_0941_),
    .S(_0942_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5028_ (.I0(\reg_file.reg_storage[12][18] ),
    .I1(\reg_file.reg_storage[13][18] ),
    .I2(\reg_file.reg_storage[14][18] ),
    .I3(\reg_file.reg_storage[15][18] ),
    .S0(_0810_),
    .S1(_0942_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5029_ (.I0(\reg_file.reg_storage[8][18] ),
    .I1(\reg_file.reg_storage[9][18] ),
    .I2(\reg_file.reg_storage[10][18] ),
    .I3(\reg_file.reg_storage[11][18] ),
    .S0(_0810_),
    .S1(_0942_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5030_ (.I(_0649_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5031_ (.I0(_0939_),
    .I1(_0943_),
    .I2(_0944_),
    .I3(_0945_),
    .S0(_0785_),
    .S1(_0946_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5032_ (.A1(_0912_),
    .A2(_0938_),
    .A3(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5033_ (.A1(_0936_),
    .A2(_0937_),
    .B(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _5034_ (.I(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5035_ (.I(_0850_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _5036_ (.I(net75),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5037_ (.I0(\reg_file.reg_storage[4][19] ),
    .I1(\reg_file.reg_storage[5][19] ),
    .I2(\reg_file.reg_storage[6][19] ),
    .I3(\reg_file.reg_storage[7][19] ),
    .S0(_0921_),
    .S1(_0922_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5038_ (.I(_0774_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5039_ (.I(\reg_file.reg_storage[1][19] ),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5040_ (.A1(_0768_),
    .A2(\reg_file.reg_storage[3][19] ),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5041_ (.I(_0772_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5042_ (.I(_0763_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5043_ (.A1(_0957_),
    .A2(\reg_file.reg_storage[2][19] ),
    .B(_0958_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5044_ (.A1(_0954_),
    .A2(_0955_),
    .B1(_0956_),
    .B2(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5045_ (.I(_0836_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5046_ (.I0(\reg_file.reg_storage[12][19] ),
    .I1(\reg_file.reg_storage[13][19] ),
    .I2(\reg_file.reg_storage[14][19] ),
    .I3(\reg_file.reg_storage[15][19] ),
    .S0(_0896_),
    .S1(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5047_ (.I0(\reg_file.reg_storage[8][19] ),
    .I1(\reg_file.reg_storage[9][19] ),
    .I2(\reg_file.reg_storage[10][19] ),
    .I3(\reg_file.reg_storage[11][19] ),
    .S0(_0921_),
    .S1(_0961_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5048_ (.I(_0784_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5049_ (.I(_0964_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5050_ (.I0(_0953_),
    .I1(_0960_),
    .I2(_0962_),
    .I3(_0963_),
    .S0(_0965_),
    .S1(_0929_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5051_ (.A1(_0754_),
    .A2(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5052_ (.A1(_0952_),
    .A2(_0913_),
    .B(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5053_ (.I(_0968_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5054_ (.I(_0830_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5055_ (.A1(_0969_),
    .A2(_0970_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5056_ (.A1(_0950_),
    .A2(_0951_),
    .B(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5057_ (.I(_0884_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5058_ (.I0(_0935_),
    .I1(_0972_),
    .S(_0973_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5059_ (.I(net32),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5060_ (.A1(_0975_),
    .A2(_0709_),
    .A3(_0710_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5061_ (.I0(_0509_),
    .I1(_0976_),
    .S(net236),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5062_ (.I(_0680_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5063_ (.I0(_0533_),
    .I1(_0977_),
    .S(_0978_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5064_ (.I(_0979_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5065_ (.I0(_0887_),
    .I1(_0974_),
    .S(_0980_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5066_ (.A1(net85),
    .A2(_0750_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5067_ (.I(_0759_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5068_ (.I(_0983_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5069_ (.I0(\reg_file.reg_storage[4][28] ),
    .I1(\reg_file.reg_storage[5][28] ),
    .I2(\reg_file.reg_storage[6][28] ),
    .I3(\reg_file.reg_storage[7][28] ),
    .S0(_0780_),
    .S1(_0984_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5070_ (.I(\reg_file.reg_storage[1][28] ),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5071_ (.A1(_0768_),
    .A2(\reg_file.reg_storage[3][28] ),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5072_ (.A1(_0957_),
    .A2(\reg_file.reg_storage[2][28] ),
    .B(_0807_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5073_ (.A1(_0954_),
    .A2(_0986_),
    .B1(_0987_),
    .B2(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5074_ (.I(_0779_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5075_ (.I0(\reg_file.reg_storage[12][28] ),
    .I1(\reg_file.reg_storage[13][28] ),
    .I2(\reg_file.reg_storage[14][28] ),
    .I3(\reg_file.reg_storage[15][28] ),
    .S0(_0990_),
    .S1(_0984_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5076_ (.I0(\reg_file.reg_storage[8][28] ),
    .I1(\reg_file.reg_storage[9][28] ),
    .I2(\reg_file.reg_storage[10][28] ),
    .I3(\reg_file.reg_storage[11][28] ),
    .S0(_0990_),
    .S1(_0984_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5077_ (.I0(_0985_),
    .I1(_0989_),
    .I2(_0991_),
    .I3(_0992_),
    .S0(_0786_),
    .S1(_0929_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5078_ (.A1(_0754_),
    .A2(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5079_ (.A1(_0982_),
    .A2(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5080_ (.I(_0995_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5081_ (.I(_0996_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5082_ (.A1(net86),
    .A2(_0889_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5083_ (.I(_0817_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5084_ (.I0(\reg_file.reg_storage[4][29] ),
    .I1(\reg_file.reg_storage[5][29] ),
    .I2(\reg_file.reg_storage[6][29] ),
    .I3(\reg_file.reg_storage[7][29] ),
    .S0(_0999_),
    .S1(_0903_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5085_ (.I(\reg_file.reg_storage[1][29] ),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5086_ (.A1(_0897_),
    .A2(\reg_file.reg_storage[3][29] ),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5087_ (.A1(_0773_),
    .A2(\reg_file.reg_storage[2][29] ),
    .B(_0899_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5088_ (.A1(_0765_),
    .A2(_1001_),
    .B1(_1002_),
    .B2(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5089_ (.I0(\reg_file.reg_storage[12][29] ),
    .I1(\reg_file.reg_storage[13][29] ),
    .I2(\reg_file.reg_storage[14][29] ),
    .I3(\reg_file.reg_storage[15][29] ),
    .S0(_0999_),
    .S1(_0903_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5090_ (.I0(\reg_file.reg_storage[8][29] ),
    .I1(\reg_file.reg_storage[9][29] ),
    .I2(\reg_file.reg_storage[10][29] ),
    .I3(\reg_file.reg_storage[11][29] ),
    .S0(_0999_),
    .S1(_0903_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5091_ (.I0(_1000_),
    .I1(_1004_),
    .I2(_1005_),
    .I3(_1006_),
    .S0(_0786_),
    .S1(_0788_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5092_ (.A1(_0891_),
    .A2(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5093_ (.A1(_0998_),
    .A2(_1008_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5094_ (.I(_1009_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5095_ (.A1(_1010_),
    .A2(_0875_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5096_ (.A1(_0997_),
    .A2(_0851_),
    .B(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5097_ (.A1(net89),
    .A2(_0750_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5098_ (.I(_0753_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5099_ (.I0(\reg_file.reg_storage[4][31] ),
    .I1(\reg_file.reg_storage[5][31] ),
    .I2(\reg_file.reg_storage[6][31] ),
    .I3(\reg_file.reg_storage[7][31] ),
    .S0(_0896_),
    .S1(_0961_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5100_ (.I(\reg_file.reg_storage[1][31] ),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5101_ (.A1(_0892_),
    .A2(\reg_file.reg_storage[3][31] ),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5102_ (.A1(_0957_),
    .A2(\reg_file.reg_storage[2][31] ),
    .B(_0958_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5103_ (.A1(_0954_),
    .A2(_1016_),
    .B1(_1017_),
    .B2(_1018_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5104_ (.I(_0633_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5105_ (.I(_1020_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5106_ (.I(_0836_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5107_ (.I0(\reg_file.reg_storage[12][31] ),
    .I1(\reg_file.reg_storage[13][31] ),
    .I2(\reg_file.reg_storage[14][31] ),
    .I3(\reg_file.reg_storage[15][31] ),
    .S0(_1021_),
    .S1(_1022_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5108_ (.I0(\reg_file.reg_storage[8][31] ),
    .I1(\reg_file.reg_storage[9][31] ),
    .I2(\reg_file.reg_storage[10][31] ),
    .I3(\reg_file.reg_storage[11][31] ),
    .S0(_0896_),
    .S1(_0961_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5109_ (.I(_0824_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5110_ (.I0(_1015_),
    .I1(_1019_),
    .I2(_1023_),
    .I3(_1024_),
    .S0(_0965_),
    .S1(_1025_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5111_ (.A1(_1014_),
    .A2(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5112_ (.A1(_1013_),
    .A2(_1027_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5113_ (.I(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5114_ (.I(_0909_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5115_ (.A1(net88),
    .A2(_0889_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5116_ (.I0(\reg_file.reg_storage[4][30] ),
    .I1(\reg_file.reg_storage[5][30] ),
    .I2(\reg_file.reg_storage[6][30] ),
    .I3(\reg_file.reg_storage[7][30] ),
    .S0(_0811_),
    .S1(_0761_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5117_ (.I(\reg_file.reg_storage[1][30] ),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5118_ (.A1(_0897_),
    .A2(\reg_file.reg_storage[3][30] ),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5119_ (.A1(_0773_),
    .A2(\reg_file.reg_storage[2][30] ),
    .B(_0775_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5120_ (.A1(_0765_),
    .A2(_1033_),
    .B1(_1034_),
    .B2(_1035_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5121_ (.I0(\reg_file.reg_storage[12][30] ),
    .I1(\reg_file.reg_storage[13][30] ),
    .I2(\reg_file.reg_storage[14][30] ),
    .I3(\reg_file.reg_storage[15][30] ),
    .S0(_0758_),
    .S1(_0761_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5122_ (.I0(\reg_file.reg_storage[8][30] ),
    .I1(\reg_file.reg_storage[9][30] ),
    .I2(\reg_file.reg_storage[10][30] ),
    .I3(\reg_file.reg_storage[11][30] ),
    .S0(_0811_),
    .S1(_0761_),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5123_ (.I0(_1032_),
    .I1(_1036_),
    .I2(_1037_),
    .I3(_1038_),
    .S0(_0786_),
    .S1(_0788_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5124_ (.A1(_0891_),
    .A2(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5125_ (.A1(_1031_),
    .A2(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5126_ (.I(_0795_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5127_ (.A1(_1041_),
    .A2(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5128_ (.A1(_1029_),
    .A2(_1030_),
    .B(_1043_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5129_ (.I0(_1012_),
    .I1(_1044_),
    .S(_0886_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5130_ (.I(net81),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5131_ (.I(_0983_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5132_ (.I0(\reg_file.reg_storage[4][24] ),
    .I1(\reg_file.reg_storage[5][24] ),
    .I2(\reg_file.reg_storage[6][24] ),
    .I3(\reg_file.reg_storage[7][24] ),
    .S0(_0767_),
    .S1(_1047_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5133_ (.I(_0778_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5134_ (.I0(\reg_file.reg_storage[2][24] ),
    .I1(\reg_file.reg_storage[3][24] ),
    .S(_1049_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5135_ (.I0(\reg_file.reg_storage[1][24] ),
    .I1(_1050_),
    .S(_1047_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5136_ (.I0(\reg_file.reg_storage[12][24] ),
    .I1(\reg_file.reg_storage[13][24] ),
    .I2(\reg_file.reg_storage[14][24] ),
    .I3(\reg_file.reg_storage[15][24] ),
    .S0(_0802_),
    .S1(_0804_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5137_ (.I0(\reg_file.reg_storage[8][24] ),
    .I1(\reg_file.reg_storage[9][24] ),
    .I2(\reg_file.reg_storage[10][24] ),
    .I3(\reg_file.reg_storage[11][24] ),
    .S0(_0767_),
    .S1(_1047_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5138_ (.I0(_1048_),
    .I1(_1051_),
    .I2(_1052_),
    .I3(_1053_),
    .S0(_0822_),
    .S1(_0871_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5139_ (.I(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5140_ (.A1(_1046_),
    .A2(_0937_),
    .B1(_0835_),
    .B2(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5141_ (.I(_1056_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5142_ (.I(_0794_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5143_ (.A1(_1057_),
    .A2(_1058_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5144_ (.A1(net82),
    .A2(_0852_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5145_ (.I(_0940_),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5146_ (.I(net8),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5147_ (.I(_1062_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5148_ (.I0(\reg_file.reg_storage[4][25] ),
    .I1(\reg_file.reg_storage[5][25] ),
    .I2(\reg_file.reg_storage[6][25] ),
    .I3(\reg_file.reg_storage[7][25] ),
    .S0(_1061_),
    .S1(_1063_),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5149_ (.I0(\reg_file.reg_storage[2][25] ),
    .I1(\reg_file.reg_storage[3][25] ),
    .S(_0920_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5150_ (.I0(\reg_file.reg_storage[1][25] ),
    .I1(_1065_),
    .S(_1063_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5151_ (.I0(\reg_file.reg_storage[12][25] ),
    .I1(\reg_file.reg_storage[13][25] ),
    .I2(\reg_file.reg_storage[14][25] ),
    .I3(\reg_file.reg_storage[15][25] ),
    .S0(_0855_),
    .S1(_0857_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5152_ (.I0(\reg_file.reg_storage[8][25] ),
    .I1(\reg_file.reg_storage[9][25] ),
    .I2(\reg_file.reg_storage[10][25] ),
    .I3(\reg_file.reg_storage[11][25] ),
    .S0(_0855_),
    .S1(_1063_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5153_ (.I0(_1064_),
    .I1(_1066_),
    .I2(_1067_),
    .I3(_1068_),
    .S0(_0870_),
    .S1(_1025_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5154_ (.A1(_0937_),
    .A2(_0938_),
    .A3(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5155_ (.A1(_1060_),
    .A2(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5156_ (.A1(_1071_),
    .A2(_0796_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5157_ (.A1(_1059_),
    .A2(_1072_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5158_ (.A1(net83),
    .A2(_0750_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5159_ (.I0(\reg_file.reg_storage[4][26] ),
    .I1(\reg_file.reg_storage[5][26] ),
    .I2(\reg_file.reg_storage[6][26] ),
    .I3(\reg_file.reg_storage[7][26] ),
    .S0(_0990_),
    .S1(_0984_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5160_ (.I(\reg_file.reg_storage[1][26] ),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5161_ (.A1(_0768_),
    .A2(\reg_file.reg_storage[3][26] ),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5162_ (.A1(_0957_),
    .A2(\reg_file.reg_storage[2][26] ),
    .B(_0958_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5163_ (.A1(_0954_),
    .A2(_1076_),
    .B1(_1077_),
    .B2(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5164_ (.I0(\reg_file.reg_storage[12][26] ),
    .I1(\reg_file.reg_storage[13][26] ),
    .I2(\reg_file.reg_storage[14][26] ),
    .I3(\reg_file.reg_storage[15][26] ),
    .S0(_0921_),
    .S1(_0922_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5165_ (.I0(\reg_file.reg_storage[8][26] ),
    .I1(\reg_file.reg_storage[9][26] ),
    .I2(\reg_file.reg_storage[10][26] ),
    .I3(\reg_file.reg_storage[11][26] ),
    .S0(_0990_),
    .S1(_0922_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5166_ (.I0(_1075_),
    .I1(_1079_),
    .I2(_1080_),
    .I3(_1081_),
    .S0(_0965_),
    .S1(_0929_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5167_ (.A1(_0754_),
    .A2(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5168_ (.A1(_1074_),
    .A2(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5169_ (.I(_1084_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5170_ (.I(_0795_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5171_ (.A1(_1085_),
    .A2(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5172_ (.I(net84),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5173_ (.I0(\reg_file.reg_storage[4][27] ),
    .I1(\reg_file.reg_storage[5][27] ),
    .I2(\reg_file.reg_storage[6][27] ),
    .I3(\reg_file.reg_storage[7][27] ),
    .S0(_1061_),
    .S1(_1063_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5174_ (.I(\reg_file.reg_storage[1][27] ),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5175_ (.A1(_0861_),
    .A2(\reg_file.reg_storage[3][27] ),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5176_ (.A1(_0863_),
    .A2(\reg_file.reg_storage[2][27] ),
    .B(_0764_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5177_ (.A1(_0899_),
    .A2(_1090_),
    .B1(_1091_),
    .B2(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5178_ (.I0(\reg_file.reg_storage[12][27] ),
    .I1(\reg_file.reg_storage[13][27] ),
    .I2(\reg_file.reg_storage[14][27] ),
    .I3(\reg_file.reg_storage[15][27] ),
    .S0(_0866_),
    .S1(_0857_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5179_ (.I0(\reg_file.reg_storage[8][27] ),
    .I1(\reg_file.reg_storage[9][27] ),
    .I2(\reg_file.reg_storage[10][27] ),
    .I3(\reg_file.reg_storage[11][27] ),
    .S0(_0855_),
    .S1(_0857_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5180_ (.I0(_1089_),
    .I1(_1093_),
    .I2(_1094_),
    .I3(_1095_),
    .S0(_0870_),
    .S1(_1025_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5181_ (.A1(_1014_),
    .A2(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5182_ (.A1(_1088_),
    .A2(_0913_),
    .B(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5183_ (.I(_1098_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5184_ (.A1(_1099_),
    .A2(_0875_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5185_ (.A1(_1087_),
    .A2(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5186_ (.I0(_1073_),
    .I1(_1101_),
    .S(_0886_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5187_ (.I(_0979_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5188_ (.I0(_1045_),
    .I1(_1102_),
    .S(_1103_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5189_ (.I(_0510_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _5190_ (.I(net2),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5191_ (.A1(_1106_),
    .A2(_0618_),
    .A3(_0616_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5192_ (.I0(_1105_),
    .I1(_1107_),
    .S(_0739_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5193_ (.I0(_0545_),
    .I1(_1108_),
    .S(_0679_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5194_ (.I(_1109_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5195_ (.I(_1110_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5196_ (.I0(_0981_),
    .I1(_1104_),
    .S(_1111_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5197_ (.I(_0720_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5198_ (.I(_0672_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5199_ (.I(_0978_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5200_ (.I(_1115_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5201_ (.A1(net159),
    .A2(_1116_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5202_ (.A1(_1114_),
    .A2(_1108_),
    .B(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5203_ (.I(_1118_),
    .Z(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5204_ (.I(_1119_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5205_ (.A1(net68),
    .A2(_0852_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5206_ (.I(_0854_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5207_ (.I(_0983_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5208_ (.I0(\reg_file.reg_storage[4][12] ),
    .I1(\reg_file.reg_storage[5][12] ),
    .I2(\reg_file.reg_storage[6][12] ),
    .I3(\reg_file.reg_storage[7][12] ),
    .S0(_1122_),
    .S1(_1123_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5209_ (.I0(\reg_file.reg_storage[2][12] ),
    .I1(\reg_file.reg_storage[3][12] ),
    .S(_0920_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5210_ (.I0(\reg_file.reg_storage[1][12] ),
    .I1(_1125_),
    .S(_1123_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5211_ (.I0(\reg_file.reg_storage[12][12] ),
    .I1(\reg_file.reg_storage[13][12] ),
    .I2(\reg_file.reg_storage[14][12] ),
    .I3(\reg_file.reg_storage[15][12] ),
    .S0(_0767_),
    .S1(_1047_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5212_ (.I0(\reg_file.reg_storage[8][12] ),
    .I1(\reg_file.reg_storage[9][12] ),
    .I2(\reg_file.reg_storage[10][12] ),
    .I3(\reg_file.reg_storage[11][12] ),
    .S0(_1122_),
    .S1(_1123_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5213_ (.I0(_1124_),
    .I1(_1126_),
    .I2(_1127_),
    .I3(_1128_),
    .S0(_0822_),
    .S1(_0871_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5214_ (.A1(_0912_),
    .A2(_0938_),
    .A3(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5215_ (.A1(_1121_),
    .A2(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5216_ (.I(_1131_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5217_ (.A1(_1132_),
    .A2(_1042_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5218_ (.I(net69),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5219_ (.I(_0635_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5220_ (.I0(\reg_file.reg_storage[4][13] ),
    .I1(\reg_file.reg_storage[5][13] ),
    .I2(\reg_file.reg_storage[6][13] ),
    .I3(\reg_file.reg_storage[7][13] ),
    .S0(_1049_),
    .S1(_1135_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5221_ (.I(\reg_file.reg_storage[1][13] ),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5222_ (.A1(_1061_),
    .A2(\reg_file.reg_storage[3][13] ),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5223_ (.A1(_0772_),
    .A2(\reg_file.reg_storage[2][13] ),
    .B(_0806_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5224_ (.A1(_0764_),
    .A2(_1137_),
    .B1(_1138_),
    .B2(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5225_ (.I(_0642_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5226_ (.I0(\reg_file.reg_storage[12][13] ),
    .I1(\reg_file.reg_storage[13][13] ),
    .I2(\reg_file.reg_storage[14][13] ),
    .I3(\reg_file.reg_storage[15][13] ),
    .S0(_1049_),
    .S1(_1141_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5227_ (.I0(\reg_file.reg_storage[8][13] ),
    .I1(\reg_file.reg_storage[9][13] ),
    .I2(\reg_file.reg_storage[10][13] ),
    .I3(\reg_file.reg_storage[11][13] ),
    .S0(_1049_),
    .S1(_1141_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5228_ (.I0(_1136_),
    .I1(_1140_),
    .I2(_1142_),
    .I3(_1143_),
    .S0(_0964_),
    .S1(_0946_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5229_ (.A1(_0890_),
    .A2(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5230_ (.A1(_1134_),
    .A2(_0912_),
    .B(_1145_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5231_ (.I(_1146_),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5232_ (.I(_0830_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5233_ (.A1(_1147_),
    .A2(_1148_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5234_ (.A1(_1133_),
    .A2(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5235_ (.A1(net70),
    .A2(_0852_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5236_ (.I0(\reg_file.reg_storage[4][14] ),
    .I1(\reg_file.reg_storage[5][14] ),
    .I2(\reg_file.reg_storage[6][14] ),
    .I3(\reg_file.reg_storage[7][14] ),
    .S0(_1021_),
    .S1(_1022_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5237_ (.I(\reg_file.reg_storage[1][14] ),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5238_ (.A1(_0892_),
    .A2(\reg_file.reg_storage[3][14] ),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5239_ (.A1(_0863_),
    .A2(\reg_file.reg_storage[2][14] ),
    .B(_0958_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5240_ (.A1(_0899_),
    .A2(_1153_),
    .B1(_1154_),
    .B2(_1155_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5241_ (.I0(\reg_file.reg_storage[12][14] ),
    .I1(\reg_file.reg_storage[13][14] ),
    .I2(\reg_file.reg_storage[14][14] ),
    .I3(\reg_file.reg_storage[15][14] ),
    .S0(_1021_),
    .S1(_1022_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5242_ (.I0(\reg_file.reg_storage[8][14] ),
    .I1(\reg_file.reg_storage[9][14] ),
    .I2(\reg_file.reg_storage[10][14] ),
    .I3(\reg_file.reg_storage[11][14] ),
    .S0(_1021_),
    .S1(_1022_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5243_ (.I0(_1152_),
    .I1(_1156_),
    .I2(_1157_),
    .I3(_1158_),
    .S0(_0965_),
    .S1(_1025_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5244_ (.A1(_1014_),
    .A2(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5245_ (.A1(_1151_),
    .A2(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5246_ (.I(_1161_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5247_ (.I(_0795_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5248_ (.A1(_1162_),
    .A2(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _5249_ (.I(net71),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5250_ (.I0(\reg_file.reg_storage[4][15] ),
    .I1(\reg_file.reg_storage[5][15] ),
    .I2(\reg_file.reg_storage[6][15] ),
    .I3(\reg_file.reg_storage[7][15] ),
    .S0(_0802_),
    .S1(_0804_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5251_ (.I(\reg_file.reg_storage[1][15] ),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5252_ (.A1(_0811_),
    .A2(\reg_file.reg_storage[3][15] ),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5253_ (.A1(_0813_),
    .A2(\reg_file.reg_storage[2][15] ),
    .B(_0814_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5254_ (.A1(_0807_),
    .A2(_1167_),
    .B1(_1168_),
    .B2(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5255_ (.I0(\reg_file.reg_storage[12][15] ),
    .I1(\reg_file.reg_storage[13][15] ),
    .I2(\reg_file.reg_storage[14][15] ),
    .I3(\reg_file.reg_storage[15][15] ),
    .S0(_0817_),
    .S1(_0818_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5256_ (.I0(\reg_file.reg_storage[8][15] ),
    .I1(\reg_file.reg_storage[9][15] ),
    .I2(\reg_file.reg_storage[10][15] ),
    .I3(\reg_file.reg_storage[11][15] ),
    .S0(_0802_),
    .S1(_0804_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5257_ (.I0(_1166_),
    .I1(_1170_),
    .I2(_1171_),
    .I3(_1172_),
    .S0(_0822_),
    .S1(_0825_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5258_ (.A1(_0800_),
    .A2(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5259_ (.A1(_1165_),
    .A2(_0937_),
    .B(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5260_ (.A1(_1175_),
    .A2(_1148_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5261_ (.A1(_1164_),
    .A2(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5262_ (.I(_0885_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5263_ (.I0(_1150_),
    .I1(_1177_),
    .S(_1178_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5264_ (.I(_0882_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5265_ (.A1(_0490_),
    .A2(net218),
    .A3(_0715_),
    .A4(_0692_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5266_ (.A1(_0978_),
    .A2(_1180_),
    .B(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5267_ (.I(_1182_),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5268_ (.I0(\reg_file.reg_storage[4][11] ),
    .I1(\reg_file.reg_storage[5][11] ),
    .I2(\reg_file.reg_storage[6][11] ),
    .I3(\reg_file.reg_storage[7][11] ),
    .S0(_0779_),
    .S1(_0942_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5269_ (.I0(\reg_file.reg_storage[2][11] ),
    .I1(\reg_file.reg_storage[3][11] ),
    .S(_0801_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5270_ (.I0(\reg_file.reg_storage[1][11] ),
    .I1(_1185_),
    .S(_1135_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5271_ (.I0(\reg_file.reg_storage[12][11] ),
    .I1(\reg_file.reg_storage[13][11] ),
    .I2(\reg_file.reg_storage[14][11] ),
    .I3(\reg_file.reg_storage[15][11] ),
    .S0(_0920_),
    .S1(_1135_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5272_ (.I0(\reg_file.reg_storage[8][11] ),
    .I1(\reg_file.reg_storage[9][11] ),
    .I2(\reg_file.reg_storage[10][11] ),
    .I3(\reg_file.reg_storage[11][11] ),
    .S0(_0779_),
    .S1(_1135_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5273_ (.I0(_1184_),
    .I1(_1186_),
    .I2(_1187_),
    .I3(_1188_),
    .S0(_0964_),
    .S1(_0946_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5274_ (.I(_1189_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5275_ (.A1(net67),
    .A2(_0888_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5276_ (.A1(_0835_),
    .A2(_1190_),
    .B(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5277_ (.I(_1192_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5278_ (.I(_1193_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5279_ (.A1(net66),
    .A2(_0888_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5280_ (.I0(\reg_file.reg_storage[4][10] ),
    .I1(\reg_file.reg_storage[5][10] ),
    .I2(\reg_file.reg_storage[6][10] ),
    .I3(\reg_file.reg_storage[7][10] ),
    .S0(_0839_),
    .S1(_0902_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5281_ (.I(\reg_file.reg_storage[1][10] ),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5282_ (.A1(_1061_),
    .A2(\reg_file.reg_storage[3][10] ),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5283_ (.A1(_0772_),
    .A2(\reg_file.reg_storage[2][10] ),
    .B(_0806_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5284_ (.A1(_0814_),
    .A2(_1197_),
    .B1(_1198_),
    .B2(_1199_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5285_ (.I0(\reg_file.reg_storage[12][10] ),
    .I1(\reg_file.reg_storage[13][10] ),
    .I2(\reg_file.reg_storage[14][10] ),
    .I3(\reg_file.reg_storage[15][10] ),
    .S0(_0839_),
    .S1(_0760_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5286_ (.I0(\reg_file.reg_storage[8][10] ),
    .I1(\reg_file.reg_storage[9][10] ),
    .I2(\reg_file.reg_storage[10][10] ),
    .I3(\reg_file.reg_storage[11][10] ),
    .S0(_0839_),
    .S1(_0760_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5287_ (.I0(_1196_),
    .I1(_1200_),
    .I2(_1201_),
    .I3(_1202_),
    .S0(_0821_),
    .S1(_0787_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5288_ (.A1(_0890_),
    .A2(_1203_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5289_ (.A1(_1195_),
    .A2(_1204_),
    .A3(_0970_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5290_ (.A1(_1194_),
    .A2(_0951_),
    .B(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5291_ (.A1(net96),
    .A2(_0749_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5292_ (.I0(\reg_file.reg_storage[4][9] ),
    .I1(\reg_file.reg_storage[5][9] ),
    .I2(\reg_file.reg_storage[6][9] ),
    .I3(\reg_file.reg_storage[7][9] ),
    .S0(_0919_),
    .S1(_0856_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5293_ (.I0(\reg_file.reg_storage[2][9] ),
    .I1(\reg_file.reg_storage[3][9] ),
    .S(_0638_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5294_ (.I0(\reg_file.reg_storage[1][9] ),
    .I1(_1209_),
    .S(_0803_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5295_ (.I0(\reg_file.reg_storage[12][9] ),
    .I1(\reg_file.reg_storage[13][9] ),
    .I2(\reg_file.reg_storage[14][9] ),
    .I3(\reg_file.reg_storage[15][9] ),
    .S0(_0778_),
    .S1(_0803_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5296_ (.I0(\reg_file.reg_storage[8][9] ),
    .I1(\reg_file.reg_storage[9][9] ),
    .I2(\reg_file.reg_storage[10][9] ),
    .I3(\reg_file.reg_storage[11][9] ),
    .S0(_0778_),
    .S1(_0803_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5297_ (.I0(_1208_),
    .I1(_1210_),
    .I2(_1211_),
    .I3(_1212_),
    .S0(_0784_),
    .S1(_0824_),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5298_ (.A1(_0621_),
    .A2(_0938_),
    .A3(_1213_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5299_ (.A1(_1207_),
    .A2(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5300_ (.I(_1215_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5301_ (.I(_1216_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5302_ (.I(_0834_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5303_ (.I0(\reg_file.reg_storage[4][8] ),
    .I1(\reg_file.reg_storage[5][8] ),
    .I2(\reg_file.reg_storage[6][8] ),
    .I3(\reg_file.reg_storage[7][8] ),
    .S0(_0940_),
    .S1(_1062_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5304_ (.I0(\reg_file.reg_storage[2][8] ),
    .I1(\reg_file.reg_storage[3][8] ),
    .S(_0919_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5305_ (.I0(\reg_file.reg_storage[1][8] ),
    .I1(_1220_),
    .S(_1062_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5306_ (.I0(\reg_file.reg_storage[12][8] ),
    .I1(\reg_file.reg_storage[13][8] ),
    .I2(\reg_file.reg_storage[14][8] ),
    .I3(\reg_file.reg_storage[15][8] ),
    .S0(_0801_),
    .S1(_0983_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5307_ (.I0(\reg_file.reg_storage[8][8] ),
    .I1(\reg_file.reg_storage[9][8] ),
    .I2(\reg_file.reg_storage[10][8] ),
    .I3(\reg_file.reg_storage[11][8] ),
    .S0(_0940_),
    .S1(_1062_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5308_ (.I0(_1219_),
    .I1(_1221_),
    .I2(_1222_),
    .I3(_1223_),
    .S0(_0821_),
    .S1(_0787_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5309_ (.I(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5310_ (.A1(net95),
    .A2(_0749_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5311_ (.A1(_1218_),
    .A2(_1225_),
    .B(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5312_ (.I(_1227_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5313_ (.A1(_1228_),
    .A2(_1058_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5314_ (.A1(_1217_),
    .A2(_1086_),
    .B(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5315_ (.A1(_1183_),
    .A2(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5316_ (.A1(_1183_),
    .A2(_1206_),
    .B(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5317_ (.I0(_1179_),
    .I1(_1232_),
    .S(_1103_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5318_ (.A1(_1120_),
    .A2(_1233_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5319_ (.I(_0543_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _5320_ (.I(net32),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5321_ (.A1(_1236_),
    .A2(_0618_),
    .A3(_0616_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5322_ (.I0(_1235_),
    .I1(_1237_),
    .S(_0738_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5323_ (.I0(net156),
    .I1(_1238_),
    .S(_0679_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5324_ (.I(_1239_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5325_ (.I(_1240_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5326_ (.I(_1183_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5327_ (.I0(\reg_file.reg_storage[4][7] ),
    .I1(\reg_file.reg_storage[5][7] ),
    .I2(\reg_file.reg_storage[6][7] ),
    .I3(\reg_file.reg_storage[7][7] ),
    .S0(_0633_),
    .S1(_0642_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5328_ (.I0(\reg_file.reg_storage[2][7] ),
    .I1(\reg_file.reg_storage[3][7] ),
    .S(_0755_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5329_ (.I0(\reg_file.reg_storage[1][7] ),
    .I1(_1244_),
    .S(_0642_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5330_ (.I0(\reg_file.reg_storage[12][7] ),
    .I1(\reg_file.reg_storage[13][7] ),
    .I2(\reg_file.reg_storage[14][7] ),
    .I3(\reg_file.reg_storage[15][7] ),
    .S0(_0644_),
    .S1(_0645_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5331_ (.I0(\reg_file.reg_storage[8][7] ),
    .I1(\reg_file.reg_storage[9][7] ),
    .I2(\reg_file.reg_storage[10][7] ),
    .I3(\reg_file.reg_storage[11][7] ),
    .S0(_0644_),
    .S1(_0645_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5332_ (.I0(_1243_),
    .I1(_1245_),
    .I2(_1246_),
    .I3(_1247_),
    .S0(_0648_),
    .S1(_0649_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5333_ (.I(_1248_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5334_ (.A1(net94),
    .A2(_0748_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5335_ (.A1(_1218_),
    .A2(_1249_),
    .B(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5336_ (.I(_1251_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5337_ (.I(_0831_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5338_ (.A1(net93),
    .A2(_0798_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5339_ (.I0(\reg_file.reg_storage[4][6] ),
    .I1(\reg_file.reg_storage[5][6] ),
    .I2(\reg_file.reg_storage[6][6] ),
    .I3(\reg_file.reg_storage[7][6] ),
    .S0(_0860_),
    .S1(_0818_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5340_ (.I(\reg_file.reg_storage[1][6] ),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5341_ (.A1(\reg_file.reg_storage[3][6] ),
    .A2(_0758_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5342_ (.A1(\reg_file.reg_storage[2][6] ),
    .A2(_0813_),
    .B(_0774_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5343_ (.A1(_1256_),
    .A2(_0807_),
    .B1(_1257_),
    .B2(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5344_ (.I0(\reg_file.reg_storage[12][6] ),
    .I1(\reg_file.reg_storage[13][6] ),
    .I2(\reg_file.reg_storage[14][6] ),
    .I3(\reg_file.reg_storage[15][6] ),
    .S0(_0860_),
    .S1(_0837_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5345_ (.I0(\reg_file.reg_storage[8][6] ),
    .I1(\reg_file.reg_storage[9][6] ),
    .I2(\reg_file.reg_storage[10][6] ),
    .I3(\reg_file.reg_storage[11][6] ),
    .S0(_0860_),
    .S1(_0837_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5346_ (.I0(_1255_),
    .I1(_1259_),
    .I2(_1260_),
    .I3(_1261_),
    .S0(_0785_),
    .S1(_0825_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5347_ (.A1(_0890_),
    .A2(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5348_ (.A1(_1254_),
    .A2(_1263_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5349_ (.I(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5350_ (.A1(_1265_),
    .A2(_0910_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5351_ (.A1(_1252_),
    .A2(_1253_),
    .B(_1266_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5352_ (.I(_1182_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5353_ (.I(_1268_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5354_ (.I(net92),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5355_ (.I(_0640_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5356_ (.I0(\reg_file.reg_storage[4][5] ),
    .I1(\reg_file.reg_storage[5][5] ),
    .I2(\reg_file.reg_storage[6][5] ),
    .I3(\reg_file.reg_storage[7][5] ),
    .S0(_0770_),
    .S1(_1271_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5357_ (.I0(\reg_file.reg_storage[2][5] ),
    .I1(\reg_file.reg_storage[3][5] ),
    .S(_0637_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5358_ (.I0(\reg_file.reg_storage[1][5] ),
    .I1(_1273_),
    .S(_1271_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5359_ (.I0(\reg_file.reg_storage[12][5] ),
    .I1(\reg_file.reg_storage[13][5] ),
    .I2(\reg_file.reg_storage[14][5] ),
    .I3(\reg_file.reg_storage[15][5] ),
    .S0(_0637_),
    .S1(_0634_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5360_ (.I0(\reg_file.reg_storage[8][5] ),
    .I1(\reg_file.reg_storage[9][5] ),
    .I2(\reg_file.reg_storage[10][5] ),
    .I3(\reg_file.reg_storage[11][5] ),
    .S0(_0637_),
    .S1(_0634_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5361_ (.I0(_1272_),
    .I1(_1274_),
    .I2(_1275_),
    .I3(_1276_),
    .S0(_0625_),
    .S1(_0823_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5362_ (.I(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5363_ (.A1(_1270_),
    .A2(_0620_),
    .B1(_0834_),
    .B2(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5364_ (.I(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5365_ (.I(_1280_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5366_ (.I(_1058_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5367_ (.A1(_1281_),
    .A2(_1282_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5368_ (.I0(\reg_file.reg_storage[4][4] ),
    .I1(\reg_file.reg_storage[5][4] ),
    .I2(\reg_file.reg_storage[6][4] ),
    .I3(\reg_file.reg_storage[7][4] ),
    .S0(_1020_),
    .S1(_1141_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5369_ (.I0(\reg_file.reg_storage[2][4] ),
    .I1(\reg_file.reg_storage[3][4] ),
    .S(_0809_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5370_ (.I0(\reg_file.reg_storage[1][4] ),
    .I1(_1285_),
    .S(_1141_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5371_ (.I0(\reg_file.reg_storage[12][4] ),
    .I1(\reg_file.reg_storage[13][4] ),
    .I2(\reg_file.reg_storage[14][4] ),
    .I3(\reg_file.reg_storage[15][4] ),
    .S0(_1020_),
    .S1(_0902_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5372_ (.I0(\reg_file.reg_storage[8][4] ),
    .I1(\reg_file.reg_storage[9][4] ),
    .I2(\reg_file.reg_storage[10][4] ),
    .I3(\reg_file.reg_storage[11][4] ),
    .S0(_1020_),
    .S1(_0902_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5373_ (.I0(_1284_),
    .I1(_1286_),
    .I2(_1287_),
    .I3(_1288_),
    .S0(_0964_),
    .S1(_0946_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5374_ (.I(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5375_ (.A1(net91),
    .A2(_0888_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5376_ (.A1(_1218_),
    .A2(_1290_),
    .B(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5377_ (.I(_1292_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5378_ (.I(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5379_ (.I(_0850_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5380_ (.A1(_1294_),
    .A2(_1295_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5381_ (.A1(_1269_),
    .A2(_1283_),
    .A3(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5382_ (.A1(_1242_),
    .A2(_1267_),
    .B(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5383_ (.I(_1178_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5384_ (.I(net87),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5385_ (.I(_0759_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5386_ (.I0(\reg_file.reg_storage[8][2] ),
    .I1(\reg_file.reg_storage[9][2] ),
    .I2(\reg_file.reg_storage[10][2] ),
    .I3(\reg_file.reg_storage[11][2] ),
    .S0(_0809_),
    .S1(_1301_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5387_ (.I0(\reg_file.reg_storage[2][2] ),
    .I1(\reg_file.reg_storage[3][2] ),
    .S(_0628_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5388_ (.I0(\reg_file.reg_storage[1][2] ),
    .I1(_1303_),
    .S(_1301_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5389_ (.I0(\reg_file.reg_storage[12][2] ),
    .I1(\reg_file.reg_storage[13][2] ),
    .I2(\reg_file.reg_storage[14][2] ),
    .I3(\reg_file.reg_storage[15][2] ),
    .S0(_0919_),
    .S1(_1301_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5390_ (.I0(\reg_file.reg_storage[4][2] ),
    .I1(\reg_file.reg_storage[5][2] ),
    .I2(\reg_file.reg_storage[6][2] ),
    .I3(\reg_file.reg_storage[7][2] ),
    .S0(_0809_),
    .S1(_1301_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5391_ (.I0(_1302_),
    .I1(_1304_),
    .I2(_1305_),
    .I3(_1306_),
    .S0(_0914_),
    .S1(net9),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5392_ (.I(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5393_ (.A1(_1300_),
    .A2(_0621_),
    .B1(_1218_),
    .B2(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5394_ (.I(_1309_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5395_ (.A1(_1310_),
    .A2(_1030_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5396_ (.A1(net90),
    .A2(_0798_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5397_ (.I0(\reg_file.reg_storage[4][3] ),
    .I1(\reg_file.reg_storage[5][3] ),
    .I2(\reg_file.reg_storage[6][3] ),
    .I3(\reg_file.reg_storage[7][3] ),
    .S0(_0866_),
    .S1(_0867_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5398_ (.I(\reg_file.reg_storage[1][3] ),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5399_ (.A1(\reg_file.reg_storage[3][3] ),
    .A2(_0999_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5400_ (.A1(\reg_file.reg_storage[2][3] ),
    .A2(_0813_),
    .B(_0814_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5401_ (.A1(_1314_),
    .A2(_0775_),
    .B1(_1315_),
    .B2(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5402_ (.I0(\reg_file.reg_storage[12][3] ),
    .I1(\reg_file.reg_storage[13][3] ),
    .I2(\reg_file.reg_storage[14][3] ),
    .I3(\reg_file.reg_storage[15][3] ),
    .S0(_1122_),
    .S1(_1123_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5403_ (.I0(\reg_file.reg_storage[8][3] ),
    .I1(\reg_file.reg_storage[9][3] ),
    .I2(\reg_file.reg_storage[10][3] ),
    .I3(\reg_file.reg_storage[11][3] ),
    .S0(_1122_),
    .S1(_0867_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5404_ (.I0(_1313_),
    .I1(_1317_),
    .I2(_1318_),
    .I3(_1319_),
    .S0(_0870_),
    .S1(_0871_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5405_ (.A1(_0800_),
    .A2(_1320_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5406_ (.A1(_1312_),
    .A2(_1321_),
    .A3(_1282_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5407_ (.A1(_1311_),
    .A2(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5408_ (.I(net76),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5409_ (.I0(\reg_file.reg_storage[4][1] ),
    .I1(\reg_file.reg_storage[5][1] ),
    .I2(\reg_file.reg_storage[6][1] ),
    .I3(\reg_file.reg_storage[7][1] ),
    .S0(_0632_),
    .S1(_0641_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5410_ (.I(\reg_file.reg_storage[1][1] ),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5411_ (.A1(\reg_file.reg_storage[3][1] ),
    .A2(_0628_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5412_ (.A1(\reg_file.reg_storage[2][1] ),
    .A2(_0771_),
    .B(_0624_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5413_ (.A1(_1326_),
    .A2(_0624_),
    .B1(_1327_),
    .B2(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5414_ (.I0(\reg_file.reg_storage[12][1] ),
    .I1(\reg_file.reg_storage[13][1] ),
    .I2(\reg_file.reg_storage[14][1] ),
    .I3(\reg_file.reg_storage[15][1] ),
    .S0(_0770_),
    .S1(_1271_),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5415_ (.I0(\reg_file.reg_storage[8][1] ),
    .I1(\reg_file.reg_storage[9][1] ),
    .I2(\reg_file.reg_storage[10][1] ),
    .I3(\reg_file.reg_storage[11][1] ),
    .S0(_0770_),
    .S1(_1271_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5416_ (.I0(_1325_),
    .I1(_1329_),
    .I2(_1330_),
    .I3(_1331_),
    .S0(_0648_),
    .S1(_0823_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5417_ (.A1(_1014_),
    .A2(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5418_ (.A1(_1324_),
    .A2(_0913_),
    .B(_1333_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5419_ (.I(_1334_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5420_ (.A1(_1335_),
    .A2(_0831_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5421_ (.I(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5422_ (.A1(_0678_),
    .A2(_1030_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5423_ (.A1(_1337_),
    .A2(_1338_),
    .B(_0973_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5424_ (.A1(_1299_),
    .A2(_1323_),
    .B(_1339_),
    .C(_1241_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5425_ (.A1(_1241_),
    .A2(_1298_),
    .B(_1340_),
    .C(_1111_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5426_ (.A1(_1234_),
    .A2(_1341_),
    .B(_0744_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5427_ (.A1(_0745_),
    .A2(_1112_),
    .B(_1113_),
    .C(_1342_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5428_ (.I(_0721_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5429_ (.A1(net24),
    .A2(_0704_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5430_ (.A1(_0729_),
    .A2(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5431_ (.A1(_1344_),
    .A2(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5432_ (.A1(_0731_),
    .A2(_1345_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5433_ (.A1(_0697_),
    .A2(_1348_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5434_ (.A1(_1338_),
    .A2(_1347_),
    .B(_0733_),
    .C(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5435_ (.I(_0736_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5436_ (.I(net25),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5437_ (.I(_1352_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5438_ (.A1(_0593_),
    .A2(_0746_),
    .A3(_0706_),
    .A4(_0657_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5439_ (.I(_1354_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5440_ (.I0(_1353_),
    .I1(net19),
    .S(_1355_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5441_ (.I(_0534_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5442_ (.I(_1357_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5443_ (.I(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5444_ (.I(_1359_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5445_ (.I(_0539_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5446_ (.I(_1361_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5447_ (.I(_1362_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5448_ (.I(_1363_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5449_ (.I0(\reg_file.reg_storage[4][26] ),
    .I1(\reg_file.reg_storage[5][26] ),
    .I2(\reg_file.reg_storage[6][26] ),
    .I3(\reg_file.reg_storage[7][26] ),
    .S0(_1360_),
    .S1(_1364_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5450_ (.I0(\reg_file.reg_storage[2][26] ),
    .I1(\reg_file.reg_storage[3][26] ),
    .S(_1359_),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5451_ (.I0(\reg_file.reg_storage[1][26] ),
    .I1(_1366_),
    .S(_1364_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5452_ (.I(_0659_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5453_ (.I(_1368_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5454_ (.I0(\reg_file.reg_storage[12][26] ),
    .I1(\reg_file.reg_storage[13][26] ),
    .I2(\reg_file.reg_storage[14][26] ),
    .I3(\reg_file.reg_storage[15][26] ),
    .S0(_1369_),
    .S1(_1364_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5455_ (.I0(\reg_file.reg_storage[8][26] ),
    .I1(\reg_file.reg_storage[9][26] ),
    .I2(\reg_file.reg_storage[10][26] ),
    .I3(\reg_file.reg_storage[11][26] ),
    .S0(_1360_),
    .S1(_1364_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5456_ (.I(_0509_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5457_ (.I0(_1365_),
    .I1(_1367_),
    .I2(_1370_),
    .I3(_1371_),
    .S0(_1372_),
    .S1(_1105_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5458_ (.A1(_0492_),
    .A2(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5459_ (.A1(_0672_),
    .A2(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5460_ (.A1(_1351_),
    .A2(_1356_),
    .B(_1375_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5461_ (.A1(_1084_),
    .A2(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5462_ (.I(_1115_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5463_ (.I(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5464_ (.I(net25),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5465_ (.I(_1380_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5466_ (.I(net18),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5467_ (.I(_1355_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5468_ (.I0(_1381_),
    .I1(_1382_),
    .S(_1383_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5469_ (.I(_0671_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5470_ (.I(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5471_ (.I(_1359_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5472_ (.I(_1363_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5473_ (.I0(\reg_file.reg_storage[4][25] ),
    .I1(\reg_file.reg_storage[5][25] ),
    .I2(\reg_file.reg_storage[6][25] ),
    .I3(\reg_file.reg_storage[7][25] ),
    .S0(_1387_),
    .S1(_1388_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5474_ (.I(_0659_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5475_ (.I0(\reg_file.reg_storage[2][25] ),
    .I1(\reg_file.reg_storage[3][25] ),
    .S(_1390_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5476_ (.I0(\reg_file.reg_storage[1][25] ),
    .I1(_1391_),
    .S(_1388_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5477_ (.I0(\reg_file.reg_storage[12][25] ),
    .I1(\reg_file.reg_storage[13][25] ),
    .I2(\reg_file.reg_storage[14][25] ),
    .I3(\reg_file.reg_storage[15][25] ),
    .S0(_1387_),
    .S1(_1388_),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5478_ (.I0(\reg_file.reg_storage[8][25] ),
    .I1(\reg_file.reg_storage[9][25] ),
    .I2(\reg_file.reg_storage[10][25] ),
    .I3(\reg_file.reg_storage[11][25] ),
    .S0(_1387_),
    .S1(_1388_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5479_ (.I(_1105_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5480_ (.I0(_1389_),
    .I1(_1392_),
    .I2(_1393_),
    .I3(_1394_),
    .S0(_1372_),
    .S1(_1395_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5481_ (.A1(_0492_),
    .A2(_1396_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5482_ (.A1(_1386_),
    .A2(_1397_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5483_ (.A1(_1379_),
    .A2(_1384_),
    .B(_1398_),
    .C(_1071_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5484_ (.I(_1378_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5485_ (.I(_1400_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5486_ (.I(_1355_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5487_ (.I0(_1353_),
    .I1(net18),
    .S(_1402_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5488_ (.I(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5489_ (.A1(_1378_),
    .A2(_1397_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5490_ (.A1(_1060_),
    .A2(_1070_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5491_ (.A1(_1401_),
    .A2(_1404_),
    .B(_1405_),
    .C(_1406_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5492_ (.A1(_1399_),
    .A2(_1407_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5493_ (.I(_1098_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5494_ (.A1(_0608_),
    .A2(_0746_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5495_ (.A1(_0728_),
    .A2(_0682_),
    .A3(_0683_),
    .A4(_1410_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5496_ (.I(_1411_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5497_ (.A1(_1352_),
    .A2(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5498_ (.I(_1413_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5499_ (.A1(net20),
    .A2(_1402_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5500_ (.A1(_1414_),
    .A2(_1415_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5501_ (.I(_1385_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5502_ (.I(_1390_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5503_ (.I(_1418_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5504_ (.I(_0539_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5505_ (.I(_1420_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5506_ (.I(_1421_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5507_ (.I(_1422_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5508_ (.I0(\reg_file.reg_storage[4][27] ),
    .I1(\reg_file.reg_storage[5][27] ),
    .I2(\reg_file.reg_storage[6][27] ),
    .I3(\reg_file.reg_storage[7][27] ),
    .S0(_1419_),
    .S1(_1423_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5509_ (.I(_1421_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5510_ (.I(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5511_ (.I(_1426_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5512_ (.I(_1359_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5513_ (.I(_1428_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5514_ (.A1(_1429_),
    .A2(\reg_file.reg_storage[3][27] ),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5515_ (.I(_0688_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5516_ (.I(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5517_ (.A1(_1432_),
    .A2(\reg_file.reg_storage[2][27] ),
    .B(_1427_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5518_ (.A1(_1427_),
    .A2(_1090_),
    .B1(_1430_),
    .B2(_1433_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5519_ (.I0(\reg_file.reg_storage[12][27] ),
    .I1(\reg_file.reg_storage[13][27] ),
    .I2(\reg_file.reg_storage[14][27] ),
    .I3(\reg_file.reg_storage[15][27] ),
    .S0(_1419_),
    .S1(_1423_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5520_ (.I0(\reg_file.reg_storage[8][27] ),
    .I1(\reg_file.reg_storage[9][27] ),
    .I2(\reg_file.reg_storage[10][27] ),
    .I3(\reg_file.reg_storage[11][27] ),
    .S0(_1419_),
    .S1(_1423_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _5521_ (.I(_1372_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5522_ (.I(_1105_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5523_ (.I0(_1424_),
    .I1(_1434_),
    .I2(_1435_),
    .I3(_1436_),
    .S0(_1437_),
    .S1(_1438_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5524_ (.A1(_0493_),
    .A2(_1417_),
    .A3(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5525_ (.A1(_1114_),
    .A2(_1416_),
    .B(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5526_ (.A1(_1409_),
    .A2(_1441_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5527_ (.I(_1412_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5528_ (.A1(_0740_),
    .A2(_1443_),
    .B(_1414_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5529_ (.I(_0491_),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5530_ (.I(_1390_),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5531_ (.I(_1363_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5532_ (.I0(\reg_file.reg_storage[4][24] ),
    .I1(\reg_file.reg_storage[5][24] ),
    .I2(\reg_file.reg_storage[6][24] ),
    .I3(\reg_file.reg_storage[7][24] ),
    .S0(_1446_),
    .S1(_1447_),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5533_ (.I0(\reg_file.reg_storage[2][24] ),
    .I1(\reg_file.reg_storage[3][24] ),
    .S(_1360_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5534_ (.I(_1421_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5535_ (.I(_1450_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5536_ (.I0(\reg_file.reg_storage[1][24] ),
    .I1(_1449_),
    .S(_1451_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5537_ (.I0(\reg_file.reg_storage[12][24] ),
    .I1(\reg_file.reg_storage[13][24] ),
    .I2(\reg_file.reg_storage[14][24] ),
    .I3(\reg_file.reg_storage[15][24] ),
    .S0(_1428_),
    .S1(_1451_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5538_ (.I0(\reg_file.reg_storage[8][24] ),
    .I1(\reg_file.reg_storage[9][24] ),
    .I2(\reg_file.reg_storage[10][24] ),
    .I3(\reg_file.reg_storage[11][24] ),
    .S0(_1446_),
    .S1(_1451_),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5539_ (.I(_1372_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5540_ (.I0(_1448_),
    .I1(_1452_),
    .I2(_1453_),
    .I3(_1454_),
    .S0(_1455_),
    .S1(_1395_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5541_ (.A1(_1445_),
    .A2(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5542_ (.A1(_1386_),
    .A2(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5543_ (.A1(_1114_),
    .A2(_1444_),
    .B(_1458_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5544_ (.A1(_1459_),
    .A2(_1056_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5545_ (.A1(_1442_),
    .A2(_1460_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5546_ (.I(_0492_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5547_ (.I(_1390_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5548_ (.I(_1463_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5549_ (.I(_1450_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5550_ (.I0(\reg_file.reg_storage[4][31] ),
    .I1(\reg_file.reg_storage[5][31] ),
    .I2(\reg_file.reg_storage[6][31] ),
    .I3(\reg_file.reg_storage[7][31] ),
    .S0(_1464_),
    .S1(_1465_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5551_ (.A1(_1429_),
    .A2(\reg_file.reg_storage[3][31] ),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5552_ (.I(_1426_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5553_ (.A1(_1432_),
    .A2(\reg_file.reg_storage[2][31] ),
    .B(_1468_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5554_ (.A1(_1427_),
    .A2(_1016_),
    .B1(_1467_),
    .B2(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5555_ (.I(_1360_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5556_ (.I0(\reg_file.reg_storage[12][31] ),
    .I1(\reg_file.reg_storage[13][31] ),
    .I2(\reg_file.reg_storage[14][31] ),
    .I3(\reg_file.reg_storage[15][31] ),
    .S0(_1471_),
    .S1(_1465_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5557_ (.I0(\reg_file.reg_storage[8][31] ),
    .I1(\reg_file.reg_storage[9][31] ),
    .I2(\reg_file.reg_storage[10][31] ),
    .I3(\reg_file.reg_storage[11][31] ),
    .S0(_1464_),
    .S1(_1465_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5558_ (.I0(_1466_),
    .I1(_1470_),
    .I2(_1472_),
    .I3(_1473_),
    .S0(_1437_),
    .S1(_1438_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5559_ (.A1(_1462_),
    .A2(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5560_ (.A1(_1353_),
    .A2(_1400_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5561_ (.A1(_1379_),
    .A2(_1475_),
    .B(_1476_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5562_ (.A1(_1029_),
    .A2(_1477_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5563_ (.I(_1411_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5564_ (.I(_1479_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5565_ (.A1(_0722_),
    .A2(_1480_),
    .B(_1413_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5566_ (.I(_1369_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5567_ (.I(_1450_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5568_ (.I0(\reg_file.reg_storage[4][30] ),
    .I1(\reg_file.reg_storage[5][30] ),
    .I2(\reg_file.reg_storage[6][30] ),
    .I3(\reg_file.reg_storage[7][30] ),
    .S0(_1482_),
    .S1(_1483_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5569_ (.A1(_1419_),
    .A2(\reg_file.reg_storage[3][30] ),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5570_ (.I(_1426_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5571_ (.A1(_1432_),
    .A2(\reg_file.reg_storage[2][30] ),
    .B(_1486_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5572_ (.A1(_1468_),
    .A2(_1033_),
    .B1(_1485_),
    .B2(_1487_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5573_ (.I(_1363_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5574_ (.I0(\reg_file.reg_storage[12][30] ),
    .I1(\reg_file.reg_storage[13][30] ),
    .I2(\reg_file.reg_storage[14][30] ),
    .I3(\reg_file.reg_storage[15][30] ),
    .S0(_1482_),
    .S1(_1489_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5575_ (.I0(\reg_file.reg_storage[8][30] ),
    .I1(\reg_file.reg_storage[9][30] ),
    .I2(\reg_file.reg_storage[10][30] ),
    .I3(\reg_file.reg_storage[11][30] ),
    .S0(_1482_),
    .S1(_1483_),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5576_ (.I0(_1484_),
    .I1(_1488_),
    .I2(_1490_),
    .I3(_1491_),
    .S0(_1455_),
    .S1(_1438_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5577_ (.A1(_1462_),
    .A2(_1492_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5578_ (.A1(_1386_),
    .A2(_1493_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5579_ (.A1(_1114_),
    .A2(_1481_),
    .B(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5580_ (.A1(_1495_),
    .A2(_1041_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5581_ (.I(net22),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5582_ (.A1(_1497_),
    .A2(_1480_),
    .B(_1413_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5583_ (.I0(\reg_file.reg_storage[4][29] ),
    .I1(\reg_file.reg_storage[5][29] ),
    .I2(\reg_file.reg_storage[6][29] ),
    .I3(\reg_file.reg_storage[7][29] ),
    .S0(_1482_),
    .S1(_1489_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5584_ (.A1(_1464_),
    .A2(\reg_file.reg_storage[3][29] ),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5585_ (.A1(_1431_),
    .A2(\reg_file.reg_storage[2][29] ),
    .B(_1486_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5586_ (.A1(_1468_),
    .A2(_1001_),
    .B1(_1500_),
    .B2(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5587_ (.I0(\reg_file.reg_storage[12][29] ),
    .I1(\reg_file.reg_storage[13][29] ),
    .I2(\reg_file.reg_storage[14][29] ),
    .I3(\reg_file.reg_storage[15][29] ),
    .S0(_1418_),
    .S1(_1489_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5588_ (.I0(\reg_file.reg_storage[8][29] ),
    .I1(\reg_file.reg_storage[9][29] ),
    .I2(\reg_file.reg_storage[10][29] ),
    .I3(\reg_file.reg_storage[11][29] ),
    .S0(_1418_),
    .S1(_1489_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5589_ (.I0(_1499_),
    .I1(_1502_),
    .I2(_1503_),
    .I3(_1504_),
    .S0(_1455_),
    .S1(_1395_),
    .Z(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5590_ (.A1(_1505_),
    .A2(_1462_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5591_ (.A1(_1351_),
    .A2(_1506_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5592_ (.A1(_1417_),
    .A2(_1498_),
    .B(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5593_ (.A1(_1009_),
    .A2(_1508_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5594_ (.A1(net21),
    .A2(_1402_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5595_ (.A1(_1413_),
    .A2(_1510_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5596_ (.I0(\reg_file.reg_storage[4][28] ),
    .I1(\reg_file.reg_storage[5][28] ),
    .I2(\reg_file.reg_storage[6][28] ),
    .I3(\reg_file.reg_storage[7][28] ),
    .S0(_1418_),
    .S1(_1447_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5597_ (.A1(_1464_),
    .A2(\reg_file.reg_storage[3][28] ),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5598_ (.A1(_1431_),
    .A2(\reg_file.reg_storage[2][28] ),
    .B(_1486_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5599_ (.A1(_1468_),
    .A2(_0986_),
    .B1(_1513_),
    .B2(_1514_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5600_ (.I0(\reg_file.reg_storage[12][28] ),
    .I1(\reg_file.reg_storage[13][28] ),
    .I2(\reg_file.reg_storage[14][28] ),
    .I3(\reg_file.reg_storage[15][28] ),
    .S0(_1446_),
    .S1(_1447_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5601_ (.I0(\reg_file.reg_storage[8][28] ),
    .I1(\reg_file.reg_storage[9][28] ),
    .I2(\reg_file.reg_storage[10][28] ),
    .I3(\reg_file.reg_storage[11][28] ),
    .S0(_1446_),
    .S1(_1447_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5602_ (.I0(_1512_),
    .I1(_1515_),
    .I2(_1516_),
    .I3(_1517_),
    .S0(_1455_),
    .S1(_1395_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5603_ (.A1(_1445_),
    .A2(_1518_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5604_ (.A1(_1351_),
    .A2(_1519_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5605_ (.A1(_1417_),
    .A2(_1511_),
    .B(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5606_ (.A1(_0995_),
    .A2(_1521_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5607_ (.A1(_1478_),
    .A2(_1496_),
    .A3(_1509_),
    .A4(_1522_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _5608_ (.A1(_1377_),
    .A2(_1408_),
    .A3(_1461_),
    .A4(_1523_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5609_ (.I0(_1423_),
    .I1(_1352_),
    .S(_1479_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5610_ (.I0(\reg_file.reg_storage[8][21] ),
    .I1(\reg_file.reg_storage[9][21] ),
    .I2(\reg_file.reg_storage[10][21] ),
    .I3(\reg_file.reg_storage[11][21] ),
    .S0(_1368_),
    .S1(_1425_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5611_ (.I0(\reg_file.reg_storage[2][21] ),
    .I1(\reg_file.reg_storage[3][21] ),
    .S(_0659_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5612_ (.I0(\reg_file.reg_storage[1][21] ),
    .I1(_1527_),
    .S(_1425_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5613_ (.I0(\reg_file.reg_storage[12][21] ),
    .I1(\reg_file.reg_storage[13][21] ),
    .I2(\reg_file.reg_storage[14][21] ),
    .I3(\reg_file.reg_storage[15][21] ),
    .S0(_1368_),
    .S1(_1421_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5614_ (.I0(\reg_file.reg_storage[4][21] ),
    .I1(\reg_file.reg_storage[5][21] ),
    .I2(\reg_file.reg_storage[6][21] ),
    .I3(\reg_file.reg_storage[7][21] ),
    .S0(_1368_),
    .S1(_1425_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5615_ (.I(_0528_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5616_ (.I(_1531_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5617_ (.I(_1532_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5618_ (.I(_1533_),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5619_ (.I(_0563_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5620_ (.I(_1535_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5621_ (.I(_1536_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5622_ (.I0(_1526_),
    .I1(_1528_),
    .I2(_1529_),
    .I3(_1530_),
    .S0(_1534_),
    .S1(_1537_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5623_ (.A1(_0491_),
    .A2(_1538_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5624_ (.A1(_0736_),
    .A2(_1539_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5625_ (.A1(_1385_),
    .A2(_1525_),
    .B(_1540_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5626_ (.I(_1541_),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5627_ (.A1(_0828_),
    .A2(_1542_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5628_ (.I(_0874_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5629_ (.I0(\reg_file.reg_storage[8][23] ),
    .I1(\reg_file.reg_storage[9][23] ),
    .I2(\reg_file.reg_storage[10][23] ),
    .I3(\reg_file.reg_storage[11][23] ),
    .S0(_1471_),
    .S1(_1465_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5630_ (.A1(_1429_),
    .A2(\reg_file.reg_storage[3][23] ),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5631_ (.A1(_1432_),
    .A2(\reg_file.reg_storage[2][23] ),
    .B(_1486_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5632_ (.A1(_1427_),
    .A2(_0859_),
    .B1(_1546_),
    .B2(_1547_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5633_ (.I0(\reg_file.reg_storage[12][23] ),
    .I1(\reg_file.reg_storage[13][23] ),
    .I2(\reg_file.reg_storage[14][23] ),
    .I3(\reg_file.reg_storage[15][23] ),
    .S0(_1471_),
    .S1(_1483_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5634_ (.I0(\reg_file.reg_storage[4][23] ),
    .I1(\reg_file.reg_storage[5][23] ),
    .I2(\reg_file.reg_storage[6][23] ),
    .I3(\reg_file.reg_storage[7][23] ),
    .S0(_1471_),
    .S1(_1483_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5635_ (.I0(_1545_),
    .I1(_1548_),
    .I2(_1549_),
    .I3(_1550_),
    .S0(_1534_),
    .S1(_1537_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5636_ (.A1(_1462_),
    .A2(_1551_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5637_ (.I0(_1438_),
    .I1(_1353_),
    .S(_1412_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5638_ (.A1(_1116_),
    .A2(_1553_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5639_ (.A1(_1400_),
    .A2(_1552_),
    .B(_1554_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5640_ (.A1(_1544_),
    .A2(_1555_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5641_ (.I0(_1429_),
    .I1(_1352_),
    .S(_1479_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5642_ (.I0(\reg_file.reg_storage[8][20] ),
    .I1(\reg_file.reg_storage[9][20] ),
    .I2(\reg_file.reg_storage[10][20] ),
    .I3(\reg_file.reg_storage[11][20] ),
    .S0(_1428_),
    .S1(_1451_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5643_ (.I0(\reg_file.reg_storage[2][20] ),
    .I1(\reg_file.reg_storage[3][20] ),
    .S(_1369_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5644_ (.I0(\reg_file.reg_storage[1][20] ),
    .I1(_1559_),
    .S(_1422_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5645_ (.I0(\reg_file.reg_storage[12][20] ),
    .I1(\reg_file.reg_storage[13][20] ),
    .I2(\reg_file.reg_storage[14][20] ),
    .I3(\reg_file.reg_storage[15][20] ),
    .S0(_1463_),
    .S1(_1422_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5646_ (.I0(\reg_file.reg_storage[4][20] ),
    .I1(\reg_file.reg_storage[5][20] ),
    .I2(\reg_file.reg_storage[6][20] ),
    .I3(\reg_file.reg_storage[7][20] ),
    .S0(_1428_),
    .S1(_1422_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5647_ (.I0(_1558_),
    .I1(_1560_),
    .I2(_1561_),
    .I3(_1562_),
    .S0(_1534_),
    .S1(_1537_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5648_ (.A1(_1445_),
    .A2(_1563_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5649_ (.A1(_1386_),
    .A2(_1564_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5650_ (.A1(_1417_),
    .A2(_1557_),
    .B(_1565_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5651_ (.A1(_0791_),
    .A2(_1566_),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5652_ (.I0(_1437_),
    .I1(_1380_),
    .S(_1412_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5653_ (.I(_1450_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5654_ (.I0(\reg_file.reg_storage[8][22] ),
    .I1(\reg_file.reg_storage[9][22] ),
    .I2(\reg_file.reg_storage[10][22] ),
    .I3(\reg_file.reg_storage[11][22] ),
    .S0(_1463_),
    .S1(_1569_),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5655_ (.I0(\reg_file.reg_storage[2][22] ),
    .I1(\reg_file.reg_storage[3][22] ),
    .S(_1369_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5656_ (.I0(\reg_file.reg_storage[1][22] ),
    .I1(_1571_),
    .S(_1569_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5657_ (.I0(\reg_file.reg_storage[12][22] ),
    .I1(\reg_file.reg_storage[13][22] ),
    .I2(\reg_file.reg_storage[14][22] ),
    .I3(\reg_file.reg_storage[15][22] ),
    .S0(_1387_),
    .S1(_1569_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5658_ (.I0(\reg_file.reg_storage[4][22] ),
    .I1(\reg_file.reg_storage[5][22] ),
    .I2(\reg_file.reg_storage[6][22] ),
    .I3(\reg_file.reg_storage[7][22] ),
    .S0(_1463_),
    .S1(_1569_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5659_ (.I0(_1570_),
    .I1(_1572_),
    .I2(_1573_),
    .I3(_1574_),
    .S0(_1534_),
    .S1(_1537_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5660_ (.A1(_1445_),
    .A2(_1385_),
    .A3(_1575_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5661_ (.A1(_0672_),
    .A2(_1568_),
    .B(_1576_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5662_ (.A1(_0849_),
    .A2(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5663_ (.A1(_1543_),
    .A2(_1556_),
    .A3(_1567_),
    .A4(_1578_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5664_ (.I(_0933_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _5665_ (.A1(_0728_),
    .A2(_0681_),
    .A3(_0683_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5666_ (.I(_1581_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _5667_ (.A1(_0706_),
    .A2(_0652_),
    .A3(_0657_),
    .B(net25),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5668_ (.I(_1583_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5669_ (.A1(_0806_),
    .A2(_1582_),
    .B(_1584_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5670_ (.I(_0792_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5671_ (.I(_1357_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5672_ (.I(_1361_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5673_ (.I0(\reg_file.reg_storage[8][16] ),
    .I1(\reg_file.reg_storage[9][16] ),
    .I2(\reg_file.reg_storage[10][16] ),
    .I3(\reg_file.reg_storage[11][16] ),
    .S0(_1587_),
    .S1(_1588_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5674_ (.I(_0566_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5675_ (.I0(\reg_file.reg_storage[2][16] ),
    .I1(\reg_file.reg_storage[3][16] ),
    .S(_1590_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5676_ (.I0(\reg_file.reg_storage[1][16] ),
    .I1(_1591_),
    .S(_1420_),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5677_ (.I0(\reg_file.reg_storage[12][16] ),
    .I1(\reg_file.reg_storage[13][16] ),
    .I2(\reg_file.reg_storage[14][16] ),
    .I3(\reg_file.reg_storage[15][16] ),
    .S0(_1587_),
    .S1(_1420_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5678_ (.I0(\reg_file.reg_storage[4][16] ),
    .I1(\reg_file.reg_storage[5][16] ),
    .I2(\reg_file.reg_storage[6][16] ),
    .I3(\reg_file.reg_storage[7][16] ),
    .S0(_1587_),
    .S1(_1420_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5679_ (.I(_1531_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5680_ (.I(_1235_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5681_ (.I0(_1589_),
    .I1(_1592_),
    .I2(_1593_),
    .I3(_1594_),
    .S0(_1595_),
    .S1(_1596_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5682_ (.A1(_1597_),
    .A2(_0490_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5683_ (.A1(_1586_),
    .A2(_1598_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5684_ (.A1(_0670_),
    .A2(_1585_),
    .B(_1599_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5685_ (.I(_1600_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5686_ (.A1(_1580_),
    .A2(_1601_),
    .Z(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5687_ (.I0(_0914_),
    .I1(_1380_),
    .S(_1581_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5688_ (.I(_0690_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _5689_ (.I(_0534_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5690_ (.I(_1605_),
    .Z(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5691_ (.I(_1606_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5692_ (.I(_0518_),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5693_ (.I(_1608_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5694_ (.I0(\reg_file.reg_storage[8][18] ),
    .I1(\reg_file.reg_storage[9][18] ),
    .I2(\reg_file.reg_storage[10][18] ),
    .I3(\reg_file.reg_storage[11][18] ),
    .S0(_1607_),
    .S1(_1609_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5695_ (.I(_0685_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5696_ (.I0(\reg_file.reg_storage[2][18] ),
    .I1(\reg_file.reg_storage[3][18] ),
    .S(_1611_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5697_ (.I0(\reg_file.reg_storage[1][18] ),
    .I1(_1612_),
    .S(_1609_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5698_ (.I(_0577_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5699_ (.I(_1614_),
    .Z(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5700_ (.I0(\reg_file.reg_storage[12][18] ),
    .I1(\reg_file.reg_storage[13][18] ),
    .I2(\reg_file.reg_storage[14][18] ),
    .I3(\reg_file.reg_storage[15][18] ),
    .S0(_1615_),
    .S1(_0879_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5701_ (.I0(\reg_file.reg_storage[4][18] ),
    .I1(\reg_file.reg_storage[5][18] ),
    .I2(\reg_file.reg_storage[6][18] ),
    .I3(\reg_file.reg_storage[7][18] ),
    .S0(_1615_),
    .S1(_1609_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5702_ (.I0(_1610_),
    .I1(_1613_),
    .I2(_1616_),
    .I3(_1617_),
    .S0(_1533_),
    .S1(_1536_),
    .Z(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5703_ (.A1(_1604_),
    .A2(_1586_),
    .A3(_1618_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5704_ (.A1(_0735_),
    .A2(_1603_),
    .B(_1619_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5705_ (.A1(_0950_),
    .A2(_1620_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5706_ (.I(_0488_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5707_ (.I(_0570_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5708_ (.I0(\reg_file.reg_storage[8][17] ),
    .I1(\reg_file.reg_storage[9][17] ),
    .I2(\reg_file.reg_storage[10][17] ),
    .I3(\reg_file.reg_storage[11][17] ),
    .S0(_0658_),
    .S1(_1623_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5709_ (.I0(\reg_file.reg_storage[2][17] ),
    .I1(\reg_file.reg_storage[3][17] ),
    .S(_0577_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5710_ (.I0(\reg_file.reg_storage[1][17] ),
    .I1(_1625_),
    .S(_1623_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5711_ (.I(_0535_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5712_ (.I0(\reg_file.reg_storage[12][17] ),
    .I1(\reg_file.reg_storage[13][17] ),
    .I2(\reg_file.reg_storage[14][17] ),
    .I3(\reg_file.reg_storage[15][17] ),
    .S0(_0658_),
    .S1(_1627_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5713_ (.I0(\reg_file.reg_storage[4][17] ),
    .I1(\reg_file.reg_storage[5][17] ),
    .I2(\reg_file.reg_storage[6][17] ),
    .I3(\reg_file.reg_storage[7][17] ),
    .S0(_0658_),
    .S1(_1627_),
    .Z(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5714_ (.I0(_1624_),
    .I1(_1626_),
    .I2(_1628_),
    .I3(_1629_),
    .S0(_1531_),
    .S1(_1235_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5715_ (.A1(_1630_),
    .A2(_1622_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5716_ (.A1(_0734_),
    .A2(_1631_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5717_ (.A1(net9),
    .A2(_0701_),
    .A3(_0682_),
    .A4(_0684_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5718_ (.A1(_0680_),
    .A2(_1583_),
    .A3(_1633_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5719_ (.A1(_0908_),
    .A2(_1632_),
    .A3(_1634_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5720_ (.A1(_1632_),
    .A2(_1634_),
    .B(_0908_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5721_ (.A1(_0626_),
    .A2(_1582_),
    .B(_1583_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5722_ (.I0(\reg_file.reg_storage[8][19] ),
    .I1(\reg_file.reg_storage[9][19] ),
    .I2(\reg_file.reg_storage[10][19] ),
    .I3(\reg_file.reg_storage[11][19] ),
    .S0(_1614_),
    .S1(_0878_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5723_ (.I0(\reg_file.reg_storage[2][19] ),
    .I1(\reg_file.reg_storage[3][19] ),
    .S(_1357_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5724_ (.I0(\reg_file.reg_storage[1][19] ),
    .I1(_1639_),
    .S(_0878_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5725_ (.I0(\reg_file.reg_storage[12][19] ),
    .I1(\reg_file.reg_storage[13][19] ),
    .I2(\reg_file.reg_storage[14][19] ),
    .I3(\reg_file.reg_storage[15][19] ),
    .S0(_0685_),
    .S1(_1623_),
    .Z(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5726_ (.I(_0567_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5727_ (.I0(\reg_file.reg_storage[4][19] ),
    .I1(\reg_file.reg_storage[5][19] ),
    .I2(\reg_file.reg_storage[6][19] ),
    .I3(\reg_file.reg_storage[7][19] ),
    .S0(_1590_),
    .S1(_1642_),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5728_ (.I0(_1638_),
    .I1(_1640_),
    .I2(_1641_),
    .I3(_1643_),
    .S0(_1532_),
    .S1(_1535_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5729_ (.A1(_1644_),
    .A2(_1622_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5730_ (.A1(_0734_),
    .A2(_1645_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5731_ (.A1(_1586_),
    .A2(_1637_),
    .B(_1646_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5732_ (.I(_1647_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5733_ (.A1(_0968_),
    .A2(net238),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5734_ (.A1(_1635_),
    .A2(_1636_),
    .B(_1649_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5735_ (.A1(_1579_),
    .A2(_1602_),
    .A3(_1621_),
    .A4(_1650_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5736_ (.A1(_0682_),
    .A2(_0684_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5737_ (.A1(_0747_),
    .A2(_0684_),
    .A3(_1410_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5738_ (.A1(_1431_),
    .A2(_0716_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5739_ (.A1(net30),
    .A2(_0716_),
    .B1(_1653_),
    .B2(_1654_),
    .C(_1652_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5740_ (.A1(_1380_),
    .A2(_1652_),
    .B(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5741_ (.I(_1627_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5742_ (.I0(\reg_file.reg_storage[8][11] ),
    .I1(\reg_file.reg_storage[9][11] ),
    .I2(\reg_file.reg_storage[10][11] ),
    .I3(\reg_file.reg_storage[11][11] ),
    .S0(_1358_),
    .S1(_1657_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5743_ (.I0(\reg_file.reg_storage[2][11] ),
    .I1(\reg_file.reg_storage[3][11] ),
    .S(_1614_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5744_ (.I0(\reg_file.reg_storage[1][11] ),
    .I1(_1659_),
    .S(_1657_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5745_ (.I0(\reg_file.reg_storage[12][11] ),
    .I1(\reg_file.reg_storage[13][11] ),
    .I2(\reg_file.reg_storage[14][11] ),
    .I3(\reg_file.reg_storage[15][11] ),
    .S0(_0686_),
    .S1(_1588_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5746_ (.I0(\reg_file.reg_storage[4][11] ),
    .I1(\reg_file.reg_storage[5][11] ),
    .I2(\reg_file.reg_storage[6][11] ),
    .I3(\reg_file.reg_storage[7][11] ),
    .S0(_0686_),
    .S1(_1588_),
    .Z(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5747_ (.I0(_1658_),
    .I1(_1660_),
    .I2(_1661_),
    .I3(_1662_),
    .S0(_1595_),
    .S1(_1596_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5748_ (.A1(_0490_),
    .A2(_1663_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5749_ (.A1(_0670_),
    .A2(_1664_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5750_ (.A1(_0735_),
    .A2(_1656_),
    .B(_1665_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5751_ (.I(_1666_),
    .Z(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5752_ (.A1(_1193_),
    .A2(_1667_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5753_ (.A1(_1195_),
    .A2(_1204_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5754_ (.I(_0734_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5755_ (.A1(_0722_),
    .A2(_1355_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5756_ (.I(_1627_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5757_ (.I0(\reg_file.reg_storage[8][10] ),
    .I1(\reg_file.reg_storage[9][10] ),
    .I2(\reg_file.reg_storage[10][10] ),
    .I3(\reg_file.reg_storage[11][10] ),
    .S0(_1358_),
    .S1(_1672_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5758_ (.I0(\reg_file.reg_storage[2][10] ),
    .I1(\reg_file.reg_storage[3][10] ),
    .S(_1614_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5759_ (.I0(\reg_file.reg_storage[1][10] ),
    .I1(_1674_),
    .S(_1672_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5760_ (.I0(\reg_file.reg_storage[12][10] ),
    .I1(\reg_file.reg_storage[13][10] ),
    .I2(\reg_file.reg_storage[14][10] ),
    .I3(\reg_file.reg_storage[15][10] ),
    .S0(_0686_),
    .S1(_1657_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5761_ (.I0(\reg_file.reg_storage[4][10] ),
    .I1(\reg_file.reg_storage[5][10] ),
    .I2(\reg_file.reg_storage[6][10] ),
    .I3(\reg_file.reg_storage[7][10] ),
    .S0(_1358_),
    .S1(_1657_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5762_ (.I0(_1673_),
    .I1(_1675_),
    .I2(_1676_),
    .I3(_1677_),
    .S0(_1595_),
    .S1(_1596_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5763_ (.A1(_1604_),
    .A2(_1678_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5764_ (.A1(_0670_),
    .A2(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5765_ (.A1(_1670_),
    .A2(_1671_),
    .B(_1680_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5766_ (.I(_1681_),
    .Z(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5767_ (.A1(_1669_),
    .A2(_1682_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5768_ (.I0(\reg_file.reg_storage[8][12] ),
    .I1(\reg_file.reg_storage[9][12] ),
    .I2(\reg_file.reg_storage[10][12] ),
    .I3(\reg_file.reg_storage[11][12] ),
    .S0(_1606_),
    .S1(_1608_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5769_ (.I0(\reg_file.reg_storage[2][12] ),
    .I1(\reg_file.reg_storage[3][12] ),
    .S(_1357_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5770_ (.I0(\reg_file.reg_storage[1][12] ),
    .I1(_1685_),
    .S(_1608_),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5771_ (.I0(\reg_file.reg_storage[12][12] ),
    .I1(\reg_file.reg_storage[13][12] ),
    .I2(\reg_file.reg_storage[14][12] ),
    .I3(\reg_file.reg_storage[15][12] ),
    .S0(_1606_),
    .S1(_0878_),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5772_ (.I0(\reg_file.reg_storage[4][12] ),
    .I1(\reg_file.reg_storage[5][12] ),
    .I2(\reg_file.reg_storage[6][12] ),
    .I3(\reg_file.reg_storage[7][12] ),
    .S0(_1606_),
    .S1(_1608_),
    .Z(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5773_ (.I0(_1684_),
    .I1(_1686_),
    .I2(_1687_),
    .I3(_1688_),
    .S0(_1532_),
    .S1(_1535_),
    .Z(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5774_ (.A1(_1622_),
    .A2(_1689_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5775_ (.I(_1690_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5776_ (.A1(_0705_),
    .A2(_1581_),
    .B(_1583_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5777_ (.I0(_1691_),
    .I1(_1692_),
    .S(_0978_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5778_ (.A1(_1131_),
    .A2(_1693_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5779_ (.I(_1588_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5780_ (.I0(\reg_file.reg_storage[8][13] ),
    .I1(\reg_file.reg_storage[9][13] ),
    .I2(\reg_file.reg_storage[10][13] ),
    .I3(\reg_file.reg_storage[11][13] ),
    .S0(_0687_),
    .S1(_1695_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5781_ (.I0(\reg_file.reg_storage[2][13] ),
    .I1(\reg_file.reg_storage[3][13] ),
    .S(_1611_),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5782_ (.I0(\reg_file.reg_storage[1][13] ),
    .I1(_1697_),
    .S(_1695_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5783_ (.I0(\reg_file.reg_storage[12][13] ),
    .I1(\reg_file.reg_storage[13][13] ),
    .I2(\reg_file.reg_storage[14][13] ),
    .I3(\reg_file.reg_storage[15][13] ),
    .S0(_0687_),
    .S1(_1695_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5784_ (.I0(\reg_file.reg_storage[4][13] ),
    .I1(\reg_file.reg_storage[5][13] ),
    .I2(\reg_file.reg_storage[6][13] ),
    .I3(\reg_file.reg_storage[7][13] ),
    .S0(_0687_),
    .S1(_1695_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5785_ (.I0(_1696_),
    .I1(_1698_),
    .I2(_1699_),
    .I3(_1700_),
    .S0(_1533_),
    .S1(_1536_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5786_ (.A1(_0491_),
    .A2(_1701_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5787_ (.A1(_1670_),
    .A2(_1702_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5788_ (.I(_1582_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5789_ (.I(_1584_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5790_ (.A1(_0727_),
    .A2(_1704_),
    .B(_1705_),
    .C(_1115_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5791_ (.A1(_1703_),
    .A2(_1706_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5792_ (.A1(_1146_),
    .A2(_1707_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5793_ (.I(_0712_),
    .Z(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5794_ (.A1(_1709_),
    .A2(_1582_),
    .B(_1584_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5795_ (.I0(\reg_file.reg_storage[8][14] ),
    .I1(\reg_file.reg_storage[9][14] ),
    .I2(\reg_file.reg_storage[10][14] ),
    .I3(\reg_file.reg_storage[11][14] ),
    .S0(_1607_),
    .S1(_1362_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5796_ (.I0(\reg_file.reg_storage[2][14] ),
    .I1(\reg_file.reg_storage[3][14] ),
    .S(_1611_),
    .Z(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5797_ (.I0(\reg_file.reg_storage[1][14] ),
    .I1(_1712_),
    .S(_1362_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5798_ (.I0(\reg_file.reg_storage[12][14] ),
    .I1(\reg_file.reg_storage[13][14] ),
    .I2(\reg_file.reg_storage[14][14] ),
    .I3(\reg_file.reg_storage[15][14] ),
    .S0(_1607_),
    .S1(_1609_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5799_ (.I0(\reg_file.reg_storage[4][14] ),
    .I1(\reg_file.reg_storage[5][14] ),
    .I2(\reg_file.reg_storage[6][14] ),
    .I3(\reg_file.reg_storage[7][14] ),
    .S0(_1607_),
    .S1(_1362_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5800_ (.I0(_1711_),
    .I1(_1713_),
    .I2(_1714_),
    .I3(_1715_),
    .S0(_1533_),
    .S1(_1536_),
    .Z(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5801_ (.A1(_1604_),
    .A2(_1716_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5802_ (.A1(_1670_),
    .A2(_1717_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5803_ (.A1(_0671_),
    .A2(_1710_),
    .B(_1718_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5804_ (.I(_1719_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5805_ (.A1(_1161_),
    .A2(_1720_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5806_ (.A1(_0863_),
    .A2(_1704_),
    .B(_1584_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5807_ (.I0(\reg_file.reg_storage[8][15] ),
    .I1(\reg_file.reg_storage[9][15] ),
    .I2(\reg_file.reg_storage[10][15] ),
    .I3(\reg_file.reg_storage[11][15] ),
    .S0(_1615_),
    .S1(_0879_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5808_ (.I0(\reg_file.reg_storage[2][15] ),
    .I1(\reg_file.reg_storage[3][15] ),
    .S(_1587_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5809_ (.I0(\reg_file.reg_storage[1][15] ),
    .I1(_1724_),
    .S(_0879_),
    .Z(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5810_ (.I0(\reg_file.reg_storage[12][15] ),
    .I1(\reg_file.reg_storage[13][15] ),
    .I2(\reg_file.reg_storage[14][15] ),
    .I3(\reg_file.reg_storage[15][15] ),
    .S0(_1611_),
    .S1(_1672_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5811_ (.I0(\reg_file.reg_storage[4][15] ),
    .I1(\reg_file.reg_storage[5][15] ),
    .I2(\reg_file.reg_storage[6][15] ),
    .I3(\reg_file.reg_storage[7][15] ),
    .S0(_1615_),
    .S1(_1672_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5812_ (.I0(_1723_),
    .I1(_1725_),
    .I2(_1726_),
    .I3(_1727_),
    .S0(_1595_),
    .S1(_1596_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5813_ (.A1(_1604_),
    .A2(_1728_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5814_ (.A1(_0735_),
    .A2(_1729_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5815_ (.A1(_1670_),
    .A2(_1722_),
    .B(_1730_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5816_ (.A1(_1175_),
    .A2(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5817_ (.A1(_1694_),
    .A2(_1708_),
    .A3(_1721_),
    .A4(_1732_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5818_ (.I(_1227_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5819_ (.A1(net21),
    .A2(_1411_),
    .B(_0669_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5820_ (.I0(\reg_file.reg_storage[8][8] ),
    .I1(\reg_file.reg_storage[9][8] ),
    .I2(\reg_file.reg_storage[10][8] ),
    .I3(\reg_file.reg_storage[11][8] ),
    .S0(_1605_),
    .S1(_1361_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5821_ (.I0(\reg_file.reg_storage[2][8] ),
    .I1(\reg_file.reg_storage[3][8] ),
    .S(_0572_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5822_ (.I0(\reg_file.reg_storage[1][8] ),
    .I1(_1737_),
    .S(_1361_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5823_ (.I0(\reg_file.reg_storage[12][8] ),
    .I1(\reg_file.reg_storage[13][8] ),
    .I2(\reg_file.reg_storage[14][8] ),
    .I3(\reg_file.reg_storage[15][8] ),
    .S0(_0577_),
    .S1(_0578_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5824_ (.I0(\reg_file.reg_storage[4][8] ),
    .I1(\reg_file.reg_storage[5][8] ),
    .I2(\reg_file.reg_storage[6][8] ),
    .I3(\reg_file.reg_storage[7][8] ),
    .S0(_1605_),
    .S1(_0578_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5825_ (.I0(_1736_),
    .I1(_1738_),
    .I2(_1739_),
    .I3(_1740_),
    .S0(_1531_),
    .S1(_1235_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5826_ (.A1(_1741_),
    .A2(_0690_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5827_ (.A1(_0669_),
    .A2(_1742_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5828_ (.A1(_1735_),
    .A2(_1743_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5829_ (.A1(_1734_),
    .A2(_1744_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5830_ (.I0(\reg_file.reg_storage[8][9] ),
    .I1(\reg_file.reg_storage[9][9] ),
    .I2(\reg_file.reg_storage[10][9] ),
    .I3(\reg_file.reg_storage[11][9] ),
    .S0(_1590_),
    .S1(_1642_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5831_ (.I0(\reg_file.reg_storage[2][9] ),
    .I1(\reg_file.reg_storage[3][9] ),
    .S(_1605_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5832_ (.I0(\reg_file.reg_storage[1][9] ),
    .I1(_1747_),
    .S(_1642_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5833_ (.I0(\reg_file.reg_storage[12][9] ),
    .I1(\reg_file.reg_storage[13][9] ),
    .I2(\reg_file.reg_storage[14][9] ),
    .I3(\reg_file.reg_storage[15][9] ),
    .S0(_0685_),
    .S1(_1623_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5834_ (.I0(\reg_file.reg_storage[4][9] ),
    .I1(\reg_file.reg_storage[5][9] ),
    .I2(\reg_file.reg_storage[6][9] ),
    .I3(\reg_file.reg_storage[7][9] ),
    .S0(_1590_),
    .S1(_1642_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5835_ (.I0(_1746_),
    .I1(_1748_),
    .I2(_1749_),
    .I3(_1750_),
    .S0(_1532_),
    .S1(_1535_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5836_ (.A1(_1622_),
    .A2(_0715_),
    .A3(_0692_),
    .A4(_1751_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _5837_ (.A1(_1497_),
    .A2(_0736_),
    .A3(_1402_),
    .B(net213),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5838_ (.A1(_1216_),
    .A2(_1753_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5839_ (.A1(_1745_),
    .A2(_1754_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5840_ (.A1(_1668_),
    .A2(_1683_),
    .A3(_1733_),
    .A4(_1755_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5841_ (.A1(_1309_),
    .A2(_1240_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5842_ (.A1(net19),
    .A2(_1116_),
    .A3(_1480_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5843_ (.A1(_0489_),
    .A2(_0575_),
    .A3(_0691_),
    .A4(_0674_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5844_ (.A1(_1758_),
    .A2(_1759_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5845_ (.A1(_1264_),
    .A2(_1760_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5846_ (.A1(_0489_),
    .A2(_0564_),
    .A3(_0673_),
    .A4(_0674_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _5847_ (.A1(_1382_),
    .A2(_0792_),
    .A3(_1354_),
    .B(_1762_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5848_ (.A1(_1280_),
    .A2(_1763_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5849_ (.I0(net160),
    .I1(_0741_),
    .S(_0680_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5850_ (.I(_1765_),
    .Z(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5851_ (.A1(_1293_),
    .A2(_1766_),
    .Z(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5852_ (.A1(_1293_),
    .A2(_1766_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5853_ (.I(net20),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5854_ (.A1(_0690_),
    .A2(_0584_),
    .A3(_0691_),
    .A4(_0692_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _5855_ (.A1(_1769_),
    .A2(_0792_),
    .A3(_1354_),
    .B(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5856_ (.I(_1771_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5857_ (.A1(_1251_),
    .A2(_1772_),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5858_ (.A1(_1767_),
    .A2(_1768_),
    .B(_1773_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5859_ (.A1(_1761_),
    .A2(_1764_),
    .A3(_1774_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5860_ (.A1(_1335_),
    .A2(_1178_),
    .Z(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5861_ (.A1(_1312_),
    .A2(_1321_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5862_ (.A1(_1777_),
    .A2(_1118_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5863_ (.A1(_1778_),
    .A2(_0697_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5864_ (.A1(_1757_),
    .A2(_1775_),
    .A3(_1776_),
    .A4(_1779_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5865_ (.A1(_1756_),
    .A2(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5866_ (.A1(_1524_),
    .A2(_1651_),
    .A3(_1781_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5867_ (.A1(net24),
    .A2(_0717_),
    .A3(_0703_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5868_ (.A1(_1344_),
    .A2(_1783_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5869_ (.A1(_1242_),
    .A2(_1253_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5870_ (.I(_1103_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5871_ (.I(_1766_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5872_ (.A1(net24),
    .A2(_0701_),
    .A3(_0715_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5873_ (.A1(_0703_),
    .A2(_1788_),
    .A3(_0723_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5874_ (.A1(_1787_),
    .A2(_1789_),
    .A3(_0719_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5875_ (.A1(_1119_),
    .A2(_1786_),
    .A3(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5876_ (.A1(_1253_),
    .A2(_1784_),
    .B1(_1785_),
    .B2(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5877_ (.A1(_1782_),
    .A2(_0726_),
    .B1(_1792_),
    .B2(_0678_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5878_ (.A1(_1343_),
    .A2(_1350_),
    .A3(_1793_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5879_ (.A1(net76),
    .A2(_0747_),
    .B1(_0752_),
    .B2(_1332_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5880_ (.A1(_0885_),
    .A2(_0676_),
    .B(_1795_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5881_ (.A1(_0885_),
    .A2(_0677_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5882_ (.A1(_1310_),
    .A2(_0979_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5883_ (.A1(_1796_),
    .A2(_1757_),
    .A3(_1797_),
    .B(_1798_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5884_ (.I(_1777_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5885_ (.A1(_1800_),
    .A2(_1119_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5886_ (.A1(_1778_),
    .A2(_1799_),
    .B(_1801_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5887_ (.A1(_1279_),
    .A2(_1763_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5888_ (.A1(net18),
    .A2(_1115_),
    .A3(_1479_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5889_ (.A1(_1804_),
    .A2(_1762_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5890_ (.A1(_1803_),
    .A2(_1293_),
    .A3(_0743_),
    .B1(_1805_),
    .B2(_1279_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5891_ (.A1(_1265_),
    .A2(_1760_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5892_ (.A1(_1761_),
    .A2(_1806_),
    .B(_1807_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5893_ (.I(_1251_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5894_ (.I(_1809_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5895_ (.A1(_1810_),
    .A2(_1772_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5896_ (.A1(_1802_),
    .A2(_1775_),
    .B1(_1808_),
    .B2(_1773_),
    .C(_1811_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5897_ (.A1(_1756_),
    .A2(_1812_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5898_ (.I(_1732_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5899_ (.A1(_1703_),
    .A2(_1706_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5900_ (.A1(_1147_),
    .A2(_1815_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5901_ (.I(_1131_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5902_ (.I(_1693_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5903_ (.A1(_1817_),
    .A2(_1818_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5904_ (.I(_1147_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5905_ (.A1(_1820_),
    .A2(_1815_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5906_ (.A1(_1816_),
    .A2(_1819_),
    .B(_1821_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5907_ (.A1(_1162_),
    .A2(_1720_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5908_ (.A1(_1721_),
    .A2(_1822_),
    .B(_1823_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5909_ (.I(_1193_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5910_ (.A1(_1825_),
    .A2(_1667_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5911_ (.I(_1744_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5912_ (.A1(_0493_),
    .A2(_1751_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5913_ (.A1(net22),
    .A2(_1411_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5914_ (.I0(_1828_),
    .I1(_1829_),
    .S(_1379_),
    .Z(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5915_ (.A1(_1228_),
    .A2(_1827_),
    .A3(_1754_),
    .B1(_1830_),
    .B2(_1216_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5916_ (.I(_1682_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5917_ (.A1(_1669_),
    .A2(_1832_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5918_ (.A1(_1683_),
    .A2(_1831_),
    .B(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5919_ (.I(_1667_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5920_ (.A1(_1194_),
    .A2(_1835_),
    .Z(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5921_ (.A1(_1826_),
    .A2(_1834_),
    .B(_1836_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5922_ (.I(_1175_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5923_ (.I(_1731_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5924_ (.A1(_1838_),
    .A2(_1839_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5925_ (.A1(_1814_),
    .A2(_1824_),
    .B1(_1837_),
    .B2(net224),
    .C(_1840_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5926_ (.A1(_1813_),
    .A2(_1841_),
    .B(_1651_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5927_ (.I(_1544_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5928_ (.I(_1555_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5929_ (.A1(_1843_),
    .A2(_1844_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5930_ (.I(_1578_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5931_ (.I(_0829_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5932_ (.I(_1541_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5933_ (.I(_0791_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5934_ (.A1(_1849_),
    .A2(_1566_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5935_ (.A1(_1847_),
    .A2(_1848_),
    .B1(_1543_),
    .B2(_1850_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5936_ (.I(_0849_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5937_ (.I(_1577_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5938_ (.A1(_1852_),
    .A2(_1853_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5939_ (.A1(_1846_),
    .A2(_1851_),
    .B(_1854_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5940_ (.A1(_1556_),
    .A2(_1855_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5941_ (.A1(_0969_),
    .A2(_1647_),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5942_ (.I(_1620_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5943_ (.A1(_0950_),
    .A2(_1858_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5944_ (.A1(net73),
    .A2(_0889_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5945_ (.A1(_0891_),
    .A2(_0907_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5946_ (.A1(_1860_),
    .A2(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5947_ (.A1(_1632_),
    .A2(_1634_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5948_ (.A1(_1862_),
    .A2(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5949_ (.A1(_1635_),
    .A2(_1636_),
    .B(_1580_),
    .C(_1601_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5950_ (.A1(_1864_),
    .A2(_1865_),
    .B(_1621_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5951_ (.A1(_1859_),
    .A2(_1866_),
    .B(_1649_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5952_ (.A1(_1857_),
    .A2(_1867_),
    .B(_1579_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5953_ (.A1(_1845_),
    .A2(_1856_),
    .A3(_1868_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5954_ (.I(_1524_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5955_ (.A1(_1842_),
    .A2(_1869_),
    .B(_1870_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5956_ (.A1(_1029_),
    .A2(_1477_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5957_ (.I(_1478_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5958_ (.I(_1495_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5959_ (.A1(_1873_),
    .A2(_1031_),
    .A3(_1040_),
    .A4(_1874_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5960_ (.A1(_1409_),
    .A2(_1441_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5961_ (.A1(_1085_),
    .A2(_1376_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5962_ (.I(_1406_),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5963_ (.A1(_1400_),
    .A2(_1403_),
    .B(_1405_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5964_ (.A1(_1878_),
    .A2(_1879_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _5965_ (.I0(_0740_),
    .I1(_1381_),
    .S(_1480_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5966_ (.A1(_1351_),
    .A2(_1457_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5967_ (.A1(_1401_),
    .A2(_1881_),
    .B(_1882_),
    .C(_1056_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5968_ (.A1(_1399_),
    .A2(_1407_),
    .B(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5969_ (.A1(_1880_),
    .A2(_1884_),
    .B(_1377_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5970_ (.A1(_1877_),
    .A2(_1885_),
    .B(_1442_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5971_ (.A1(net205),
    .A2(_1522_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5972_ (.A1(_1876_),
    .A2(_1886_),
    .B(_1887_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5973_ (.A1(_1401_),
    .A2(_1511_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5974_ (.A1(_1401_),
    .A2(_1519_),
    .B(_1889_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5975_ (.A1(net204),
    .A2(_0997_),
    .A3(_1890_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5976_ (.A1(_1010_),
    .A2(_1508_),
    .B(_1891_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5977_ (.A1(_1888_),
    .A2(_1892_),
    .B(_1873_),
    .C(net237),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5978_ (.A1(_1872_),
    .A2(_1875_),
    .A3(_1893_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5979_ (.A1(_1873_),
    .A2(_0721_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5980_ (.A1(_1871_),
    .A2(_1894_),
    .B(_1895_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5981_ (.A1(_1782_),
    .A2(_0718_),
    .A3(_1789_),
    .Z(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5982_ (.A1(_1895_),
    .A2(_1871_),
    .A3(_1894_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5983_ (.A1(_1896_),
    .A2(_1897_),
    .A3(_1898_),
    .Z(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5984_ (.A1(_0697_),
    .A2(_0733_),
    .B1(_1794_),
    .B2(_1899_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5985_ (.I(_1900_),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5986_ (.I(_1901_),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5987_ (.I(_0696_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5988_ (.A1(_0702_),
    .A2(_0724_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5989_ (.A1(_1903_),
    .A2(_0730_),
    .B(_0695_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5990_ (.A1(_1795_),
    .A2(net227),
    .A3(_1904_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5991_ (.A1(_1902_),
    .A2(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5992_ (.A1(_0720_),
    .A2(_0726_),
    .A3(_0732_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5993_ (.A1(_1862_),
    .A2(_0910_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5994_ (.A1(_0949_),
    .A2(_0951_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5995_ (.A1(_0968_),
    .A2(_1163_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5996_ (.A1(_0791_),
    .A2(_1148_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5997_ (.A1(_1268_),
    .A2(_1910_),
    .A3(_1911_),
    .Z(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5998_ (.A1(_0973_),
    .A2(_1908_),
    .A3(_1909_),
    .B(_1912_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5999_ (.A1(_1057_),
    .A2(_0970_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6000_ (.A1(_1544_),
    .A2(_0851_),
    .B(_1914_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6001_ (.A1(_1847_),
    .A2(_1148_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6002_ (.A1(_0849_),
    .A2(_0796_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6003_ (.A1(_1916_),
    .A2(_1917_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6004_ (.I0(_1915_),
    .I1(_1918_),
    .S(_1268_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6005_ (.I0(_1913_),
    .I1(_1919_),
    .S(_1240_),
    .Z(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6006_ (.A1(_1041_),
    .A2(_0910_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6007_ (.A1(_1010_),
    .A2(_0831_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6008_ (.A1(_1921_),
    .A2(_1922_),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6009_ (.I(_1042_),
    .Z(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6010_ (.A1(_1029_),
    .A2(_1183_),
    .A3(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6011_ (.A1(_1269_),
    .A2(_1923_),
    .B(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6012_ (.A1(_1084_),
    .A2(_1058_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6013_ (.A1(_1071_),
    .A2(_1086_),
    .B(_1927_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6014_ (.A1(_0996_),
    .A2(_1163_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6015_ (.A1(_1098_),
    .A2(_0850_),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6016_ (.A1(_1929_),
    .A2(_1930_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6017_ (.I0(_1928_),
    .I1(_1931_),
    .S(_1178_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6018_ (.A1(_0980_),
    .A2(_1932_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6019_ (.A1(_0980_),
    .A2(_1926_),
    .B(_1933_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6020_ (.I0(_1920_),
    .I1(_1934_),
    .S(_1110_),
    .Z(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6021_ (.A1(_1281_),
    .A2(_1295_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6022_ (.I(_1936_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6023_ (.I(_1265_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6024_ (.A1(_1938_),
    .A2(_1295_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6025_ (.A1(_1252_),
    .A2(_1086_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6026_ (.A1(_1734_),
    .A2(_1282_),
    .B(_1940_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6027_ (.A1(_1299_),
    .A2(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6028_ (.A1(_1299_),
    .A2(_1937_),
    .A3(_1939_),
    .B(_1942_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6029_ (.A1(_1294_),
    .A2(_1282_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6030_ (.A1(_1800_),
    .A2(_1924_),
    .B(_1944_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6031_ (.A1(_1795_),
    .A2(_1295_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6032_ (.I(_1310_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6033_ (.A1(_1947_),
    .A2(_0851_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6034_ (.A1(_1269_),
    .A2(_1946_),
    .A3(_1948_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6035_ (.A1(_1269_),
    .A2(_1945_),
    .B(_1949_),
    .C(_0980_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6036_ (.A1(_1786_),
    .A2(_1943_),
    .B(_1950_),
    .C(_1119_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6037_ (.A1(_1175_),
    .A2(_1163_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6038_ (.A1(_0933_),
    .A2(_0970_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6039_ (.A1(_1952_),
    .A2(_1953_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6040_ (.I(_1162_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6041_ (.A1(_1147_),
    .A2(_1042_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6042_ (.A1(_1955_),
    .A2(_1030_),
    .B(_1956_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6043_ (.I0(_1954_),
    .I1(_1957_),
    .S(_1268_),
    .Z(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6044_ (.I(_1669_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6045_ (.A1(_1217_),
    .A2(_0875_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6046_ (.A1(_1959_),
    .A2(_0951_),
    .B(_1960_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6047_ (.A1(_1193_),
    .A2(_0909_),
    .Z(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6048_ (.A1(_1121_),
    .A2(_1130_),
    .A3(_0909_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6049_ (.A1(_1962_),
    .A2(_1963_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6050_ (.A1(_0886_),
    .A2(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6051_ (.A1(_0973_),
    .A2(_1961_),
    .B(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6052_ (.I0(_1958_),
    .I1(_1966_),
    .S(_1103_),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6053_ (.A1(_1111_),
    .A2(_1967_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6054_ (.A1(_0744_),
    .A2(_1951_),
    .A3(_1968_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6055_ (.A1(_0744_),
    .A2(_1935_),
    .B(_1969_),
    .C(_1113_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6056_ (.I(_1299_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6057_ (.A1(_1795_),
    .A2(_1242_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6058_ (.A1(_0721_),
    .A2(_1783_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6059_ (.A1(_1972_),
    .A2(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6060_ (.A1(_1972_),
    .A2(_1348_),
    .B(_1974_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6061_ (.A1(_1335_),
    .A2(_1971_),
    .B1(_1347_),
    .B2(_1975_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6062_ (.I(_1242_),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6063_ (.A1(_1977_),
    .A2(_1902_),
    .A3(_1946_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6064_ (.A1(_1791_),
    .A2(_1978_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6065_ (.A1(_1907_),
    .A2(_1970_),
    .A3(_1976_),
    .A4(_1979_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6066_ (.A1(_0733_),
    .A2(_1906_),
    .B(_1980_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6067_ (.I(_1981_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6068_ (.I(_1982_),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6069_ (.I(_1907_),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6070_ (.I(_1983_),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6071_ (.A1(_1182_),
    .A2(_1904_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6072_ (.A1(_1335_),
    .A2(_1985_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6073_ (.A1(_1902_),
    .A2(_1905_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6074_ (.A1(_1182_),
    .A2(_0694_),
    .B1(_1903_),
    .B2(_0730_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6075_ (.A1(_0979_),
    .A2(_1988_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6076_ (.A1(_1310_),
    .A2(_1989_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6077_ (.A1(_1986_),
    .A2(_1987_),
    .B(_1990_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6078_ (.A1(_1334_),
    .A2(_1985_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6079_ (.A1(_0696_),
    .A2(_1905_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6080_ (.A1(_1309_),
    .A2(_1989_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6081_ (.A1(_1992_),
    .A2(_1993_),
    .A3(_1994_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6082_ (.A1(_1991_),
    .A2(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6083_ (.I(_1907_),
    .Z(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6084_ (.I(_0745_),
    .Z(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6085_ (.I(_1998_),
    .Z(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6086_ (.I(_1999_),
    .Z(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6087_ (.I(_1120_),
    .Z(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6088_ (.I(_2001_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6089_ (.I(_1241_),
    .Z(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6090_ (.I(_2003_),
    .Z(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6091_ (.I(_2004_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6092_ (.I(_1977_),
    .Z(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6093_ (.I(_2006_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6094_ (.I(_2007_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6095_ (.I0(_1012_),
    .I1(_1101_),
    .S(_2008_),
    .Z(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6096_ (.I(_2003_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6097_ (.I(_2006_),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6098_ (.I(_2011_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6099_ (.A1(_2012_),
    .A2(_1044_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6100_ (.A1(_2010_),
    .A2(_2013_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6101_ (.A1(_2005_),
    .A2(_2009_),
    .B(_2014_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6102_ (.I(_1120_),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6103_ (.I(_2016_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6104_ (.I(_1971_),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6105_ (.I0(_0877_),
    .I1(_1073_),
    .S(_2018_),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6106_ (.I0(_0833_),
    .I1(_0972_),
    .S(_2011_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6107_ (.I(_1786_),
    .Z(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6108_ (.I(_2021_),
    .Z(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6109_ (.I0(_2019_),
    .I1(_2020_),
    .S(_2022_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6110_ (.A1(_2017_),
    .A2(_2023_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6111_ (.A1(_2002_),
    .A2(_2015_),
    .B(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6112_ (.I(_1998_),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6113_ (.I(_2016_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6114_ (.I(_1977_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6115_ (.I(_2028_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6116_ (.I(_2007_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6117_ (.A1(_2030_),
    .A2(_1267_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6118_ (.A1(_2029_),
    .A2(_1230_),
    .B(_2031_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6119_ (.A1(_2005_),
    .A2(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6120_ (.I(_1971_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6121_ (.I(_2034_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6122_ (.I(_2035_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6123_ (.I(_2034_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6124_ (.I(_2037_),
    .Z(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6125_ (.A1(_2038_),
    .A2(_1283_),
    .A3(_1296_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6126_ (.I(_2021_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6127_ (.I(_2040_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6128_ (.A1(_2036_),
    .A2(_1323_),
    .B(_2039_),
    .C(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6129_ (.A1(_2027_),
    .A2(_2033_),
    .A3(_2042_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6130_ (.I(_1111_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6131_ (.I(_2044_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6132_ (.I(_2045_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6133_ (.I(_2006_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6134_ (.I0(_0935_),
    .I1(_1177_),
    .S(_2047_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6135_ (.I(_2034_),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6136_ (.A1(_2037_),
    .A2(_1150_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6137_ (.A1(_2049_),
    .A2(_1206_),
    .B(_2050_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6138_ (.I(_2021_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6139_ (.I0(_2048_),
    .I1(_2051_),
    .S(_2052_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6140_ (.A1(_2046_),
    .A2(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6141_ (.A1(_2026_),
    .A2(_2043_),
    .A3(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6142_ (.I(_1113_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6143_ (.I(_2056_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6144_ (.A1(_2000_),
    .A2(_2025_),
    .B(_2055_),
    .C(_2057_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6145_ (.I(_2044_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6146_ (.I(_2059_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6147_ (.I(_2060_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6148_ (.I(_1241_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6149_ (.I(_2062_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6150_ (.I(_2063_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6151_ (.I(_0745_),
    .Z(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6152_ (.A1(_1789_),
    .A2(_0719_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6153_ (.I(_2066_),
    .Z(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6154_ (.A1(_2065_),
    .A2(_2067_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6155_ (.A1(_2061_),
    .A2(_2064_),
    .A3(_2068_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6156_ (.A1(_1311_),
    .A2(_1337_),
    .B(_2018_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6157_ (.A1(_2049_),
    .A2(_0677_),
    .B(_2070_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6158_ (.A1(_2069_),
    .A2(_2071_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6159_ (.I(_1347_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6160_ (.I(_2073_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6161_ (.I(_2074_),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6162_ (.I(_1348_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6163_ (.I(_2076_),
    .Z(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6164_ (.A1(_1947_),
    .A2(_2064_),
    .B(_2077_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6165_ (.I(_2004_),
    .Z(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6166_ (.I(_1973_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6167_ (.I(_2080_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6168_ (.A1(_1947_),
    .A2(_2079_),
    .A3(_2081_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6169_ (.A1(_2075_),
    .A2(_2078_),
    .A3(_2082_),
    .B1(_2064_),
    .B2(_1947_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6170_ (.A1(_1997_),
    .A2(_2058_),
    .A3(_2072_),
    .A4(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6171_ (.A1(_1984_),
    .A2(_1996_),
    .B(_2084_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _6172_ (.I(_2085_),
    .ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6173_ (.I(_0733_),
    .Z(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6174_ (.I(_2086_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _6175_ (.A1(_1239_),
    .A2(_0884_),
    .A3(_0793_),
    .B1(_0729_),
    .B2(_0725_),
    .B3(_0713_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6176_ (.A1(_1110_),
    .A2(net203),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6177_ (.A1(_1800_),
    .A2(_2089_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6178_ (.A1(_1777_),
    .A2(_2089_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6179_ (.A1(_2090_),
    .A2(_2091_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6180_ (.A1(_1309_),
    .A2(_1989_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6181_ (.A1(_1992_),
    .A2(_1993_),
    .B(_1994_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6182_ (.A1(_2093_),
    .A2(_2094_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6183_ (.A1(_2092_),
    .A2(_2095_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6184_ (.I(_1971_),
    .Z(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6185_ (.I0(_1915_),
    .I1(_1928_),
    .S(_2097_),
    .Z(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6186_ (.A1(_2097_),
    .A2(_1918_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6187_ (.A1(_2034_),
    .A2(_1910_),
    .A3(_1911_),
    .B(_2099_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6188_ (.I(_2040_),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6189_ (.I0(_2098_),
    .I1(_2100_),
    .S(_2101_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6190_ (.I(_1028_),
    .Z(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6191_ (.I(_1977_),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6192_ (.I(_2104_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6193_ (.I(_1253_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6194_ (.I(_2106_),
    .Z(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6195_ (.A1(_2103_),
    .A2(_2105_),
    .A3(_2107_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6196_ (.I(_1786_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6197_ (.I(_2109_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6198_ (.I0(_1931_),
    .I1(_1923_),
    .S(_2097_),
    .Z(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6199_ (.A1(_2110_),
    .A2(_2111_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6200_ (.A1(_2041_),
    .A2(_2108_),
    .B(_2112_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6201_ (.I(_2044_),
    .Z(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6202_ (.I0(_2102_),
    .I1(_2113_),
    .S(_2114_),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6203_ (.I(_2060_),
    .Z(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6204_ (.I(_2008_),
    .Z(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6205_ (.A1(_2012_),
    .A2(_1941_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6206_ (.A1(_2117_),
    .A2(_1961_),
    .B(_2118_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6207_ (.I(_2109_),
    .Z(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6208_ (.I(_2097_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6209_ (.I(_2121_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6210_ (.A1(_1937_),
    .A2(_1939_),
    .B(_2122_),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6211_ (.A1(_2120_),
    .A2(_2123_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6212_ (.A1(_2117_),
    .A2(_1945_),
    .B(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6213_ (.A1(_2079_),
    .A2(_2119_),
    .B(_2125_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6214_ (.A1(_2006_),
    .A2(_1954_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6215_ (.A1(_2104_),
    .A2(_1908_),
    .A3(_1909_),
    .B(_2127_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6216_ (.I0(_1957_),
    .I1(_1964_),
    .S(_2028_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6217_ (.I0(_2128_),
    .I1(_2129_),
    .S(_2022_),
    .Z(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6218_ (.A1(_2046_),
    .A2(_2130_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6219_ (.A1(_2116_),
    .A2(_2126_),
    .B(_2131_),
    .C(_2026_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6220_ (.A1(_2000_),
    .A2(_2115_),
    .B(_2132_),
    .C(_2057_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6221_ (.I(_1800_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6222_ (.I(_2060_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6223_ (.A1(_2134_),
    .A2(_2135_),
    .B(_2077_),
    .ZN(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6224_ (.I(_2059_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6225_ (.A1(_2134_),
    .A2(_2137_),
    .A3(_2081_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6226_ (.I(_2059_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6227_ (.I(_2139_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6228_ (.A1(_2075_),
    .A2(_2136_),
    .A3(_2138_),
    .B1(_2140_),
    .B2(_2134_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6229_ (.I(_1924_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6230_ (.A1(_2134_),
    .A2(_2142_),
    .B(_1948_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6231_ (.A1(_2121_),
    .A2(_1902_),
    .A3(_1946_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6232_ (.A1(_2035_),
    .A2(_2143_),
    .B(_2144_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6233_ (.A1(_2069_),
    .A2(_2145_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _6234_ (.A1(_2133_),
    .A2(_2141_),
    .A3(_2146_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6235_ (.A1(_2087_),
    .A2(_2096_),
    .B(_2147_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _6236_ (.I(_2148_),
    .ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6237_ (.A1(_2093_),
    .A2(_2091_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6238_ (.A1(_1777_),
    .A2(_2089_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6239_ (.A1(_2094_),
    .A2(_2149_),
    .B(_2150_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6240_ (.A1(_1903_),
    .A2(_0730_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6241_ (.I(_2152_),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _6242_ (.A1(_1109_),
    .A2(_1239_),
    .A3(_0883_),
    .A4(_0793_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6243_ (.I(_2154_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6244_ (.A1(_2153_),
    .A2(_2155_),
    .B(_1766_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6245_ (.A1(_1903_),
    .A2(_0731_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6246_ (.A1(_1110_),
    .A2(_1240_),
    .A3(_0884_),
    .A4(_0794_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6247_ (.A1(_0743_),
    .A2(_2157_),
    .A3(_2158_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6248_ (.A1(_2156_),
    .A2(_2159_),
    .B(_1292_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6249_ (.I(_2160_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6250_ (.A1(_1292_),
    .A2(_2156_),
    .A3(_2159_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6251_ (.A1(_2161_),
    .A2(_2162_),
    .Z(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6252_ (.A1(_2151_),
    .A2(_2163_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6253_ (.I(_2086_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6254_ (.A1(_2151_),
    .A2(_2163_),
    .B(_2165_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6255_ (.I(_1784_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6256_ (.I(_2167_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6257_ (.I(_2168_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6258_ (.A1(_0731_),
    .A2(_1345_),
    .Z(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6259_ (.I(_2170_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6260_ (.A1(_1768_),
    .A2(_2171_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6261_ (.A1(_1344_),
    .A2(_1346_),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6262_ (.I(_2173_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6263_ (.A1(_1768_),
    .A2(_2169_),
    .B(_2172_),
    .C(_2174_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6264_ (.I(_2065_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6265_ (.I(_2045_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6266_ (.I0(_0887_),
    .I1(_1102_),
    .S(_2063_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6267_ (.I(_2044_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6268_ (.A1(_2041_),
    .A2(_1045_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6269_ (.A1(_2179_),
    .A2(_2180_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6270_ (.A1(_2177_),
    .A2(_2178_),
    .B(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6271_ (.I(_2040_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6272_ (.I0(_1232_),
    .I1(_1298_),
    .S(_2183_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6273_ (.I(_2021_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6274_ (.A1(_2185_),
    .A2(_0974_),
    .Z(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6275_ (.A1(_2063_),
    .A2(_1179_),
    .B(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6276_ (.A1(_2114_),
    .A2(_2187_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6277_ (.I(_1998_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6278_ (.A1(_2177_),
    .A2(_2184_),
    .B(_2188_),
    .C(_2189_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6279_ (.A1(_2176_),
    .A2(_2182_),
    .B(_2190_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6280_ (.I(_1790_),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6281_ (.I(_2192_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6282_ (.I(_2121_),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6283_ (.A1(_1296_),
    .A2(_1322_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6284_ (.A1(_2049_),
    .A2(_1311_),
    .A3(_1337_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6285_ (.A1(_2194_),
    .A2(_2195_),
    .B(_2196_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6286_ (.I(_2109_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6287_ (.A1(_2198_),
    .A2(_2194_),
    .A3(_0677_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6288_ (.A1(_2041_),
    .A2(_2197_),
    .B(_2199_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6289_ (.A1(_2140_),
    .A2(_2200_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _6290_ (.A1(_1767_),
    .A2(_2175_),
    .B1(_2191_),
    .B2(_2057_),
    .C1(_2193_),
    .C2(_2201_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6291_ (.A1(_2164_),
    .A2(_2166_),
    .B(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6292_ (.I(_2203_),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6293_ (.A1(_1765_),
    .A2(_2155_),
    .B(_2153_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6294_ (.A1(_1280_),
    .A2(_1805_),
    .A3(_2204_),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6295_ (.I(_2164_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6296_ (.A1(_2161_),
    .A2(_2206_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6297_ (.A1(_2205_),
    .A2(_2207_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6298_ (.I(_0745_),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6299_ (.I(_2209_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6300_ (.I0(_1919_),
    .I1(_1932_),
    .S(_2062_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6301_ (.A1(_2004_),
    .A2(_1926_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6302_ (.I0(_2211_),
    .I1(_2212_),
    .S(_2045_),
    .Z(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6303_ (.I(_2016_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6304_ (.I0(_1958_),
    .I1(_1913_),
    .S(_2062_),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6305_ (.A1(_2214_),
    .A2(_2215_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6306_ (.I(_2062_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6307_ (.A1(_2052_),
    .A2(_1943_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6308_ (.A1(_2217_),
    .A2(_1966_),
    .B(_2218_),
    .C(_2045_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6309_ (.A1(_2216_),
    .A2(_2219_),
    .B(_1999_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6310_ (.A1(_2210_),
    .A2(_2213_),
    .B(_2220_),
    .C(_2056_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6311_ (.A1(_1944_),
    .A2(_1936_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6312_ (.I0(_2143_),
    .I1(_2222_),
    .S(_2105_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6313_ (.I0(_1978_),
    .I1(_2223_),
    .S(_2198_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6314_ (.A1(_2046_),
    .A2(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6315_ (.A1(_1281_),
    .A2(_1805_),
    .A3(_0718_),
    .B1(_1764_),
    .B2(_1344_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6316_ (.A1(_2192_),
    .A2(_2225_),
    .B1(_2226_),
    .B2(_1345_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6317_ (.A1(_1997_),
    .A2(_2208_),
    .B(_2221_),
    .C(_2227_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6318_ (.I(_2228_),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6319_ (.I(net19),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6320_ (.A1(_2229_),
    .A2(_0669_),
    .A3(_1354_),
    .B(_1759_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6321_ (.I(_2230_),
    .Z(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _6322_ (.A1(_1765_),
    .A2(_1763_),
    .Z(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6323_ (.A1(_2155_),
    .A2(_2232_),
    .B(_2152_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6324_ (.A1(_2231_),
    .A2(_2233_),
    .Z(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6325_ (.A1(_1264_),
    .A2(_2234_),
    .Z(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6326_ (.I(_2235_),
    .Z(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6327_ (.A1(_2161_),
    .A2(_2162_),
    .A3(_2205_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6328_ (.A1(_2094_),
    .A2(_2149_),
    .B(_2237_),
    .C(_2150_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6329_ (.A1(_1805_),
    .A2(_2204_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6330_ (.A1(_1281_),
    .A2(_2239_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6331_ (.A1(_1280_),
    .A2(_2239_),
    .B(_2160_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6332_ (.A1(_2240_),
    .A2(_2241_),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6333_ (.A1(_2238_),
    .A2(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6334_ (.A1(_2236_),
    .A2(_2243_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6335_ (.I(_2183_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6336_ (.I(_2120_),
    .Z(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6337_ (.A1(_2246_),
    .A2(_2032_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6338_ (.I(_2001_),
    .Z(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6339_ (.A1(_2245_),
    .A2(_2051_),
    .B(_2247_),
    .C(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6340_ (.I0(_2048_),
    .I1(_2020_),
    .S(_2063_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6341_ (.I(_1787_),
    .Z(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6342_ (.A1(_2116_),
    .A2(_2250_),
    .B(_2251_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6343_ (.I0(_2019_),
    .I1(_2009_),
    .S(_2010_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6344_ (.A1(_2110_),
    .A2(_2029_),
    .A3(_1044_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6345_ (.A1(_2179_),
    .A2(_2254_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6346_ (.A1(_2135_),
    .A2(_2253_),
    .B(_2255_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6347_ (.I(_1787_),
    .Z(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6348_ (.A1(_0704_),
    .A2(_0719_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6349_ (.I(_2258_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6350_ (.A1(_2249_),
    .A2(_2252_),
    .B1(_2256_),
    .B2(_2257_),
    .C(_2259_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6351_ (.I(_2214_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6352_ (.A1(_2104_),
    .A2(_1283_),
    .A3(_1266_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6353_ (.A1(_2028_),
    .A2(_2195_),
    .B(_2262_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6354_ (.I0(_2071_),
    .I1(_2263_),
    .S(_2022_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6355_ (.A1(_2261_),
    .A2(_2264_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6356_ (.I(_2073_),
    .Z(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6357_ (.A1(_1938_),
    .A2(_2231_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6358_ (.I(_2167_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6359_ (.I(_2170_),
    .Z(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6360_ (.A1(_2267_),
    .A2(_2269_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6361_ (.A1(_2267_),
    .A2(_2268_),
    .B(_2270_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6362_ (.A1(_1938_),
    .A2(_2231_),
    .B1(_2266_),
    .B2(_2271_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6363_ (.A1(_2068_),
    .A2(_2265_),
    .B(_2272_),
    .C(_1983_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6364_ (.A1(_2260_),
    .A2(_2273_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6365_ (.A1(_2087_),
    .A2(_2244_),
    .B(_2274_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6366_ (.I(_2275_),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6367_ (.A1(_2231_),
    .A2(_2154_),
    .A3(_2232_),
    .B(_2152_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6368_ (.A1(_1771_),
    .A2(_2276_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6369_ (.A1(_1809_),
    .A2(_2277_),
    .Z(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6370_ (.I(_2278_),
    .Z(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6371_ (.A1(_1938_),
    .A2(_2234_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6372_ (.A1(_2238_),
    .A2(_2242_),
    .B(_2236_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6373_ (.A1(_2280_),
    .A2(_2281_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6374_ (.A1(_2279_),
    .A2(_2282_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6375_ (.I(_2189_),
    .Z(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6376_ (.I0(_2098_),
    .I1(_2111_),
    .S(_2003_),
    .Z(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6377_ (.A1(_2079_),
    .A2(_2108_),
    .B(_2179_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6378_ (.A1(_2116_),
    .A2(_2285_),
    .B(_2286_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6379_ (.I(_2016_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6380_ (.I(_2288_),
    .Z(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6381_ (.I0(_2128_),
    .I1(_2100_),
    .S(_2003_),
    .Z(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6382_ (.A1(_2246_),
    .A2(_2119_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6383_ (.A1(_2079_),
    .A2(_2129_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6384_ (.A1(_2248_),
    .A2(_2291_),
    .A3(_2292_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6385_ (.A1(_2289_),
    .A2(_2290_),
    .B(_2293_),
    .C(_2176_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6386_ (.A1(_2284_),
    .A2(_2287_),
    .B(_2294_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6387_ (.I(_2056_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6388_ (.I(_2104_),
    .Z(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6389_ (.A1(_1939_),
    .A2(_1940_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6390_ (.A1(_2047_),
    .A2(_2298_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6391_ (.A1(_2297_),
    .A2(_2222_),
    .B(_2299_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6392_ (.I0(_2145_),
    .I1(_2300_),
    .S(_2185_),
    .Z(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6393_ (.A1(_2261_),
    .A2(_2301_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6394_ (.A1(_1252_),
    .A2(_1772_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6395_ (.I(_2170_),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6396_ (.A1(_2303_),
    .A2(_2304_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6397_ (.A1(_2303_),
    .A2(_2169_),
    .B(_2305_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6398_ (.A1(_1252_),
    .A2(_1772_),
    .B1(_2075_),
    .B2(_2306_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6399_ (.A1(_2068_),
    .A2(_2302_),
    .B(_2307_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6400_ (.A1(_2087_),
    .A2(_2283_),
    .B1(_2295_),
    .B2(_2296_),
    .C(_2308_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _6401_ (.I(_2309_),
    .ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6402_ (.A1(_2235_),
    .A2(_2279_),
    .Z(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6403_ (.A1(_1265_),
    .A2(_2234_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6404_ (.A1(_1810_),
    .A2(_2277_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6405_ (.A1(_2311_),
    .A2(_2312_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6406_ (.A1(_1810_),
    .A2(_2277_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6407_ (.A1(_2240_),
    .A2(_2235_),
    .A3(_2241_),
    .A4(_2278_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6408_ (.A1(_2238_),
    .A2(_2310_),
    .B1(_2313_),
    .B2(_2314_),
    .C(_2315_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6409_ (.A1(_2230_),
    .A2(_1771_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _6410_ (.A1(_2155_),
    .A2(_2232_),
    .A3(net217),
    .B(_2152_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6411_ (.A1(_1744_),
    .A2(_2318_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6412_ (.A1(_1228_),
    .A2(_2319_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6413_ (.A1(_2316_),
    .A2(_2320_),
    .Z(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6414_ (.A1(_2316_),
    .A2(_2320_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6415_ (.A1(_2165_),
    .A2(_2321_),
    .A3(_2322_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6416_ (.I(_2139_),
    .Z(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6417_ (.A1(_2324_),
    .A2(_1233_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6418_ (.I(_2209_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6419_ (.A1(_2261_),
    .A2(_0981_),
    .B(_2326_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6420_ (.A1(_2065_),
    .A2(_2114_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6421_ (.A1(_1104_),
    .A2(_2328_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6422_ (.A1(_2325_),
    .A2(_2327_),
    .B(_2329_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6423_ (.A1(_2245_),
    .A2(_1797_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6424_ (.I(_1120_),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6425_ (.I(_2332_),
    .Z(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6426_ (.A1(_2037_),
    .A2(_1283_),
    .A3(_1266_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6427_ (.I(_1924_),
    .Z(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6428_ (.A1(_1810_),
    .A2(_2335_),
    .B(_1229_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6429_ (.A1(_2028_),
    .A2(_2336_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6430_ (.A1(_2334_),
    .A2(_2337_),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6431_ (.I0(_2197_),
    .I1(_2338_),
    .S(_2183_),
    .Z(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6432_ (.A1(_2333_),
    .A2(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6433_ (.A1(_2289_),
    .A2(_2331_),
    .B(_2340_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6434_ (.I(_2192_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6435_ (.I(_1734_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6436_ (.A1(_2343_),
    .A2(_1827_),
    .B(_2171_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6437_ (.I(_2073_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6438_ (.A1(_2343_),
    .A2(_1827_),
    .A3(_2268_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6439_ (.A1(_2345_),
    .A2(_2346_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6440_ (.A1(_2343_),
    .A2(_1827_),
    .B1(_2344_),
    .B2(_2347_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6441_ (.A1(_2296_),
    .A2(_2330_),
    .B1(_2341_),
    .B2(_2342_),
    .C(_2348_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6442_ (.A1(_2323_),
    .A2(_2349_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _6443_ (.I(_2350_),
    .ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6444_ (.I(_1907_),
    .Z(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6445_ (.I(_2351_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6446_ (.A1(_1744_),
    .A2(_2157_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6447_ (.A1(_2318_),
    .A2(_2353_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6448_ (.A1(_1215_),
    .A2(_1753_),
    .A3(_2354_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6449_ (.A1(_2343_),
    .A2(_2319_),
    .B(_2321_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6450_ (.A1(_2355_),
    .A2(_2356_),
    .Z(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6451_ (.I0(_1967_),
    .I1(_1920_),
    .S(_2137_),
    .Z(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6452_ (.A1(_1934_),
    .A2(_2328_),
    .B1(_2358_),
    .B2(_2284_),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6453_ (.I(_2004_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6454_ (.A1(_2360_),
    .A2(_1978_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6455_ (.I(_2022_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6456_ (.I(_2106_),
    .Z(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6457_ (.A1(_1228_),
    .A2(_2363_),
    .B(_1960_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6458_ (.A1(_2018_),
    .A2(_2298_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6459_ (.A1(_2035_),
    .A2(_2364_),
    .B(_2365_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6460_ (.A1(_2110_),
    .A2(_2366_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6461_ (.A1(_2362_),
    .A2(_2223_),
    .B(_2367_),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6462_ (.A1(_2333_),
    .A2(_2368_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6463_ (.A1(_2289_),
    .A2(_2361_),
    .B(_2369_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6464_ (.I(_1217_),
    .Z(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6465_ (.I(_2173_),
    .Z(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6466_ (.I(_2080_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6467_ (.I(_2076_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6468_ (.A1(_2371_),
    .A2(_1830_),
    .B(_2374_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6469_ (.A1(_2371_),
    .A2(_1830_),
    .A3(_2373_),
    .B(_2375_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6470_ (.A1(_2371_),
    .A2(_1830_),
    .B1(_2372_),
    .B2(_2376_),
    .ZN(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6471_ (.A1(_2342_),
    .A2(_2370_),
    .B(_2377_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6472_ (.A1(_2352_),
    .A2(_2357_),
    .B1(_2359_),
    .B2(_2259_),
    .C(_2378_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6473_ (.I(_2379_),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6474_ (.A1(_2110_),
    .A2(_2071_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6475_ (.A1(_1216_),
    .A2(_2363_),
    .B(_1205_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6476_ (.A1(_2121_),
    .A2(_2336_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6477_ (.A1(_2037_),
    .A2(_2381_),
    .B(_2382_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6478_ (.I0(_2263_),
    .I1(_2383_),
    .S(_2109_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6479_ (.A1(_2332_),
    .A2(_2384_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6480_ (.A1(_2288_),
    .A2(_2380_),
    .B(_2385_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6481_ (.I(_1959_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6482_ (.A1(_2387_),
    .A2(_1832_),
    .B(_2077_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6483_ (.A1(_2387_),
    .A2(_1832_),
    .A3(_2373_),
    .B(_2388_),
    .ZN(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6484_ (.A1(_2387_),
    .A2(_1832_),
    .B1(_2372_),
    .B2(_2389_),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6485_ (.A1(_2320_),
    .A2(_2355_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6486_ (.A1(_1753_),
    .A2(_2318_),
    .A3(_2353_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6487_ (.A1(_2318_),
    .A2(_2353_),
    .B(_1753_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6488_ (.A1(_2392_),
    .A2(_2393_),
    .B(_2371_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6489_ (.A1(_1217_),
    .A2(_2392_),
    .A3(_2393_),
    .B1(_2319_),
    .B2(_1734_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6490_ (.A1(_2394_),
    .A2(_2395_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6491_ (.A1(_2316_),
    .A2(_2391_),
    .B(_2396_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6492_ (.I(_2157_),
    .Z(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _6493_ (.A1(_1735_),
    .A2(_1743_),
    .B1(_1829_),
    .B2(_1586_),
    .C(_1752_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6494_ (.A1(_2154_),
    .A2(_2232_),
    .A3(_2317_),
    .A4(_2399_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6495_ (.A1(_2398_),
    .A2(net207),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6496_ (.A1(_1669_),
    .A2(_1681_),
    .A3(_2401_),
    .Z(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6497_ (.A1(_2397_),
    .A2(_2402_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6498_ (.I(_2086_),
    .Z(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6499_ (.A1(_2397_),
    .A2(_2402_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6500_ (.A1(_2404_),
    .A2(_2405_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6501_ (.A1(_1787_),
    .A2(_2001_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6502_ (.A1(_2114_),
    .A2(_2053_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6503_ (.A1(_2027_),
    .A2(_2023_),
    .B(_2065_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6504_ (.A1(_2015_),
    .A2(_2407_),
    .B1(_2408_),
    .B2(_2409_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6505_ (.A1(_2057_),
    .A2(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6506_ (.A1(_2403_),
    .A2(_2406_),
    .B(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6507_ (.A1(_2342_),
    .A2(_2386_),
    .B(_2390_),
    .C(_2412_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6508_ (.I(net233),
    .ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6509_ (.A1(_1681_),
    .A2(net208),
    .B(_2157_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6510_ (.A1(_1192_),
    .A2(_1666_),
    .A3(_2414_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6511_ (.A1(_1682_),
    .A2(_2401_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6512_ (.A1(_1959_),
    .A2(_2416_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6513_ (.A1(_2417_),
    .A2(_2405_),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6514_ (.A1(_2415_),
    .A2(_2418_),
    .Z(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6515_ (.I0(_2130_),
    .I1(_2102_),
    .S(_2179_),
    .Z(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6516_ (.I(_1999_),
    .Z(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6517_ (.A1(_2113_),
    .A2(_2328_),
    .B1(_2420_),
    .B2(_2421_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6518_ (.A1(_2246_),
    .A2(_2145_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6519_ (.I(_2332_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6520_ (.A1(_2387_),
    .A2(_2335_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6521_ (.A1(_1962_),
    .A2(_2425_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6522_ (.A1(_2011_),
    .A2(_2426_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6523_ (.A1(_2297_),
    .A2(_2364_),
    .B(_2427_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6524_ (.I0(_2300_),
    .I1(_2428_),
    .S(_2198_),
    .Z(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6525_ (.A1(_2424_),
    .A2(_2429_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6526_ (.A1(_2002_),
    .A2(_2423_),
    .B(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6527_ (.I(_1825_),
    .Z(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6528_ (.A1(_2432_),
    .A2(_1835_),
    .B(_2076_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6529_ (.A1(_2432_),
    .A2(_1835_),
    .A3(_2080_),
    .B(_2433_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6530_ (.A1(_2432_),
    .A2(_1835_),
    .B1(_2173_),
    .B2(_2434_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6531_ (.A1(_2193_),
    .A2(_2431_),
    .B(_2435_),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6532_ (.A1(_2259_),
    .A2(_2422_),
    .B(_2436_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6533_ (.A1(_2087_),
    .A2(_2419_),
    .B(_2437_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _6534_ (.I(_2438_),
    .ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6535_ (.I(_2153_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6536_ (.A1(_1666_),
    .A2(_1682_),
    .A3(net206),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6537_ (.A1(_2439_),
    .A2(_2440_),
    .Z(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6538_ (.A1(_1818_),
    .A2(_2441_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6539_ (.A1(_1132_),
    .A2(_2442_),
    .Z(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6540_ (.I(_2443_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6541_ (.A1(_2402_),
    .A2(_2415_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6542_ (.A1(_1667_),
    .A2(_2414_),
    .Z(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _6543_ (.A1(_1959_),
    .A2(_2416_),
    .B1(_2446_),
    .B2(_1194_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6544_ (.A1(_1194_),
    .A2(_2446_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6545_ (.A1(_2391_),
    .A2(_2445_),
    .Z(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _6546_ (.A1(_2396_),
    .A2(_2445_),
    .B1(_2447_),
    .B2(_2448_),
    .C1(_2449_),
    .C2(_2316_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6547_ (.A1(_2444_),
    .A2(_2450_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6548_ (.A1(_2093_),
    .A2(_2091_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6549_ (.A1(_2161_),
    .A2(_2162_),
    .A3(_2205_),
    .Z(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6550_ (.A1(_1991_),
    .A2(_2452_),
    .B(_2453_),
    .C(_2090_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6551_ (.A1(_2236_),
    .A2(_2279_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6552_ (.A1(_2240_),
    .A2(_2236_),
    .A3(_2241_),
    .A4(_2279_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6553_ (.A1(_2311_),
    .A2(_2312_),
    .B(_2314_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6554_ (.A1(_2454_),
    .A2(_2455_),
    .B(_2456_),
    .C(_2457_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6555_ (.A1(_2391_),
    .A2(_2445_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6556_ (.A1(_2396_),
    .A2(_2445_),
    .B1(_2447_),
    .B2(_2448_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6557_ (.A1(_2458_),
    .A2(_2459_),
    .B(_2460_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6558_ (.A1(_2443_),
    .A2(_2461_),
    .B(_2351_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6559_ (.I(_2407_),
    .Z(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6560_ (.A1(_2027_),
    .A2(_2187_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6561_ (.A1(_2248_),
    .A2(_2178_),
    .B(_2464_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _6562_ (.A1(_2180_),
    .A2(_2463_),
    .B1(_2465_),
    .B2(_2257_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6563_ (.A1(_2432_),
    .A2(_2142_),
    .B(_1133_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6564_ (.A1(_2011_),
    .A2(_2467_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6565_ (.A1(_2297_),
    .A2(_2381_),
    .B(_2468_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6566_ (.I0(_2338_),
    .I1(_2469_),
    .S(_2052_),
    .Z(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6567_ (.A1(_2288_),
    .A2(_2470_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6568_ (.A1(_2017_),
    .A2(_2200_),
    .B(_2471_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6569_ (.A1(_2193_),
    .A2(_2472_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6570_ (.A1(_1132_),
    .A2(_1818_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6571_ (.A1(_2474_),
    .A2(_2269_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6572_ (.A1(_2474_),
    .A2(_2268_),
    .B(_2475_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6573_ (.A1(_1132_),
    .A2(_1818_),
    .B1(_2266_),
    .B2(_2476_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6574_ (.A1(_2473_),
    .A2(_2477_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6575_ (.A1(_2451_),
    .A2(_2462_),
    .B1(_2466_),
    .B2(_2296_),
    .C(_2478_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _6576_ (.I(_2479_),
    .ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6577_ (.A1(_1817_),
    .A2(_2442_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6578_ (.A1(_2444_),
    .A2(_2450_),
    .B(_2480_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6579_ (.I(_1820_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6580_ (.I(_1707_),
    .Z(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6581_ (.I(_2439_),
    .Z(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6582_ (.I(_1693_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6583_ (.A1(_1666_),
    .A2(_2485_),
    .A3(_1681_),
    .A4(net209),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6584_ (.A1(_2484_),
    .A2(_2486_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6585_ (.A1(_2483_),
    .A2(_2487_),
    .Z(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6586_ (.A1(_2482_),
    .A2(_2488_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6587_ (.A1(_2481_),
    .A2(_2489_),
    .Z(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6588_ (.I0(_2215_),
    .I1(_2211_),
    .S(_2060_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6589_ (.I(_2209_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6590_ (.A1(_2212_),
    .A2(_2328_),
    .B1(_2491_),
    .B2(_2492_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6591_ (.I(_1820_),
    .Z(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6592_ (.A1(_2494_),
    .A2(_2483_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6593_ (.I(_2170_),
    .Z(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6594_ (.A1(_2495_),
    .A2(_2496_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6595_ (.A1(_2495_),
    .A2(_2268_),
    .B(_2497_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _6596_ (.A1(_2494_),
    .A2(_2483_),
    .B1(_2266_),
    .B2(_2498_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6597_ (.A1(_2494_),
    .A2(_2142_),
    .B(_1963_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6598_ (.A1(_2018_),
    .A2(_2426_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6599_ (.A1(_2035_),
    .A2(_2500_),
    .B(_2501_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6600_ (.I0(_2366_),
    .I1(_2502_),
    .S(_2185_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6601_ (.A1(_2288_),
    .A2(_2503_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6602_ (.A1(_2017_),
    .A2(_2224_),
    .B(_2504_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6603_ (.A1(_2193_),
    .A2(_2505_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6604_ (.A1(_2259_),
    .A2(_2493_),
    .B(_2499_),
    .C(_2506_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6605_ (.A1(_2165_),
    .A2(_2490_),
    .B(_2507_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _6606_ (.I(_2508_),
    .ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6607_ (.I(_1955_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6608_ (.I(_1720_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6609_ (.A1(_2483_),
    .A2(_2486_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6610_ (.A1(_2398_),
    .A2(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6611_ (.A1(_2510_),
    .A2(_2512_),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6612_ (.I(_2513_),
    .Z(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6613_ (.A1(_1815_),
    .A2(_2487_),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6614_ (.A1(_1817_),
    .A2(_2442_),
    .B1(_2515_),
    .B2(_2482_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6615_ (.A1(_2494_),
    .A2(_2488_),
    .B(_2516_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6616_ (.A1(_2443_),
    .A2(_2461_),
    .A3(_2489_),
    .B(_2517_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6617_ (.A1(_2509_),
    .A2(_2514_),
    .A3(_2518_),
    .Z(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6618_ (.A1(_2135_),
    .A2(_2250_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6619_ (.A1(_2248_),
    .A2(_2253_),
    .B(_2026_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6620_ (.A1(_2254_),
    .A2(_2407_),
    .B1(_2520_),
    .B2(_2521_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6621_ (.A1(_1149_),
    .A2(_1164_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6622_ (.I0(_2467_),
    .I1(_2523_),
    .S(_2047_),
    .Z(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6623_ (.I0(_2383_),
    .I1(_2524_),
    .S(_2052_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6624_ (.I0(_2264_),
    .I1(_2525_),
    .S(_2001_),
    .Z(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6625_ (.A1(_2509_),
    .A2(_2510_),
    .B(_2374_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6626_ (.A1(_2509_),
    .A2(_2510_),
    .A3(_2081_),
    .B(_2527_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6627_ (.A1(_2509_),
    .A2(_2510_),
    .B1(_2372_),
    .B2(_2528_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6628_ (.A1(_2296_),
    .A2(_2522_),
    .B1(_2526_),
    .B2(_2342_),
    .C(_2529_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6629_ (.A1(_1984_),
    .A2(_2519_),
    .B(_2530_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6630_ (.I(_2531_),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6631_ (.I(_1838_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6632_ (.I(_1162_),
    .Z(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6633_ (.A1(_2533_),
    .A2(_2514_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6634_ (.A1(_2533_),
    .A2(_2514_),
    .Z(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6635_ (.A1(_2518_),
    .A2(_2534_),
    .B(_2535_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6636_ (.I(_2398_),
    .Z(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6637_ (.A1(_1720_),
    .A2(_2511_),
    .B(_2537_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6638_ (.A1(_1731_),
    .A2(_2538_),
    .Z(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6639_ (.I(_2539_),
    .Z(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6640_ (.A1(_2532_),
    .A2(_2536_),
    .A3(_2540_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6641_ (.A1(_2103_),
    .A2(_2158_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6642_ (.I0(_2290_),
    .I1(_2285_),
    .S(_2059_),
    .Z(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6643_ (.A1(_2251_),
    .A2(_2543_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6644_ (.A1(_2251_),
    .A2(_2542_),
    .B(_2544_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6645_ (.A1(_1955_),
    .A2(_2335_),
    .B(_1952_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6646_ (.A1(_2047_),
    .A2(_2546_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6647_ (.A1(_2297_),
    .A2(_2500_),
    .B(_2547_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6648_ (.I0(_2428_),
    .I1(_2548_),
    .S(_2185_),
    .Z(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6649_ (.I0(_2301_),
    .I1(_2549_),
    .S(_2332_),
    .Z(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6650_ (.I(_2532_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6651_ (.A1(_2551_),
    .A2(_1839_),
    .B(_2496_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6652_ (.A1(_2551_),
    .A2(_1839_),
    .A3(_2167_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6653_ (.A1(_2073_),
    .A2(_2553_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6654_ (.A1(_2551_),
    .A2(_1839_),
    .B1(_2552_),
    .B2(_2554_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6655_ (.A1(_2056_),
    .A2(_2545_),
    .B1(_2550_),
    .B2(_2192_),
    .C(_2555_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6656_ (.A1(_1997_),
    .A2(_2541_),
    .B(_2556_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6657_ (.I(_2557_),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6658_ (.A1(_2532_),
    .A2(_2540_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6659_ (.A1(_2532_),
    .A2(_2540_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6660_ (.A1(_2536_),
    .A2(_2558_),
    .B(_2559_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6661_ (.I(_2560_),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6662_ (.I(_1601_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6663_ (.A1(_1719_),
    .A2(_1731_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6664_ (.I(_2153_),
    .Z(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6665_ (.A1(_1707_),
    .A2(_2486_),
    .A3(_2563_),
    .B(_2564_),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6666_ (.A1(_2562_),
    .A2(_2565_),
    .Z(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6667_ (.A1(_1580_),
    .A2(_2566_),
    .Z(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6668_ (.A1(_2561_),
    .A2(_2567_),
    .B(_1983_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6669_ (.A1(_2561_),
    .A2(_2567_),
    .B(_2568_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6670_ (.A1(_2251_),
    .A2(_2258_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6671_ (.I(_2570_),
    .Z(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6672_ (.A1(_1112_),
    .A2(_2571_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6673_ (.I(_1580_),
    .Z(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6674_ (.I(_2345_),
    .Z(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6675_ (.A1(_2573_),
    .A2(_2562_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6676_ (.I(_2167_),
    .Z(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6677_ (.I(_2576_),
    .Z(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6678_ (.I(_2304_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6679_ (.A1(_2575_),
    .A2(_2578_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6680_ (.A1(_2575_),
    .A2(_2577_),
    .B(_2579_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6681_ (.A1(_2573_),
    .A2(_2562_),
    .B1(_2574_),
    .B2(_2580_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6682_ (.I(_2066_),
    .Z(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6683_ (.I(_2582_),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6684_ (.A1(_2261_),
    .A2(_2339_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6685_ (.I(_2139_),
    .Z(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6686_ (.A1(_0934_),
    .A2(_1176_),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6687_ (.I0(_2523_),
    .I1(_2586_),
    .S(_2105_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6688_ (.I0(_2469_),
    .I1(_2587_),
    .S(_2120_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6689_ (.A1(_2585_),
    .A2(_2588_),
    .B(_2326_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6690_ (.A1(_2463_),
    .A2(_2331_),
    .B1(_2584_),
    .B2(_2589_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6691_ (.A1(_2583_),
    .A2(_2590_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6692_ (.A1(_2569_),
    .A2(_2572_),
    .A3(_2581_),
    .A4(_2591_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6693_ (.I(_2592_),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6694_ (.I(_1862_),
    .Z(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6695_ (.A1(_1601_),
    .A2(_2398_),
    .B(_2565_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6696_ (.A1(_1863_),
    .A2(_2594_),
    .Z(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6697_ (.A1(_2593_),
    .A2(_2595_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6698_ (.A1(_2593_),
    .A2(_2595_),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6699_ (.A1(_2596_),
    .A2(_2597_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6700_ (.A1(_2573_),
    .A2(_2566_),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6701_ (.A1(_2561_),
    .A2(_2567_),
    .B(_2599_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6702_ (.A1(_2598_),
    .A2(_2600_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6703_ (.A1(_2424_),
    .A2(_2368_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6704_ (.A1(_0908_),
    .A2(_2363_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6705_ (.A1(_2573_),
    .A2(_2107_),
    .B(_2603_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6706_ (.A1(_2049_),
    .A2(_2546_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6707_ (.A1(_2194_),
    .A2(_2604_),
    .B(_2605_),
    .ZN(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6708_ (.I0(_2502_),
    .I1(_2606_),
    .S(_2198_),
    .Z(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6709_ (.A1(_2177_),
    .A2(_2607_),
    .B(_2189_),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6710_ (.A1(_2407_),
    .A2(_2361_),
    .B1(_2602_),
    .B2(_2608_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6711_ (.I(_2067_),
    .Z(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6712_ (.A1(_1635_),
    .A2(_2171_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6713_ (.A1(_1635_),
    .A2(_2169_),
    .B(_2611_),
    .C(_2174_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6714_ (.A1(_1935_),
    .A2(_2570_),
    .B1(_2609_),
    .B2(_2610_),
    .C1(_1636_),
    .C2(_2612_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6715_ (.A1(_1984_),
    .A2(_2601_),
    .B(_2613_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6716_ (.I(_2614_),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6717_ (.A1(_2025_),
    .A2(_2571_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6718_ (.I(_0949_),
    .Z(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6719_ (.A1(_2616_),
    .A2(_1858_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6720_ (.A1(_2617_),
    .A2(_2578_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6721_ (.A1(_2617_),
    .A2(_2577_),
    .B(_2618_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6722_ (.A1(_2616_),
    .A2(_1858_),
    .B1(_2574_),
    .B2(_2619_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6723_ (.A1(_2593_),
    .A2(_2595_),
    .Z(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6724_ (.A1(_2599_),
    .A2(_2621_),
    .Z(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6725_ (.I(_2567_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6726_ (.A1(_2623_),
    .A2(_2598_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6727_ (.A1(_2597_),
    .A2(_2622_),
    .B1(_2624_),
    .B2(_2560_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6728_ (.A1(_1600_),
    .A2(_1863_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6729_ (.A1(_2564_),
    .A2(_2626_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6730_ (.A1(_2565_),
    .A2(_2627_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6731_ (.A1(_1858_),
    .A2(_2628_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6732_ (.A1(_0950_),
    .A2(_2629_),
    .Z(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6733_ (.A1(_2625_),
    .A2(_2630_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6734_ (.A1(_2625_),
    .A2(_2630_),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6735_ (.A1(_1997_),
    .A2(_2632_),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6736_ (.I(_2214_),
    .Z(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6737_ (.A1(_2634_),
    .A2(_2384_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6738_ (.I0(_2616_),
    .I1(_2593_),
    .S(_2335_),
    .Z(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6739_ (.I0(_2586_),
    .I1(_2636_),
    .S(_2007_),
    .Z(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6740_ (.I0(_2524_),
    .I1(_2637_),
    .S(_2101_),
    .Z(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6741_ (.A1(_2324_),
    .A2(_2638_),
    .B(_2326_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6742_ (.A1(_2463_),
    .A2(_2380_),
    .B1(_2635_),
    .B2(_2639_),
    .ZN(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6743_ (.I(_2067_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6744_ (.A1(_2631_),
    .A2(_2633_),
    .B1(_2640_),
    .B2(_2641_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _6745_ (.A1(_2615_),
    .A2(_2620_),
    .A3(_2642_),
    .ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6746_ (.A1(_2115_),
    .A2(_2571_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6747_ (.I(_0969_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6748_ (.A1(_2644_),
    .A2(net239),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6749_ (.A1(_2645_),
    .A2(_2578_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6750_ (.A1(_2645_),
    .A2(_2577_),
    .B(_2646_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6751_ (.A1(_2644_),
    .A2(net240),
    .B1(_2574_),
    .B2(_2647_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6752_ (.A1(_1620_),
    .A2(_2439_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6753_ (.A1(_2565_),
    .A2(_2627_),
    .A3(_2649_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6754_ (.A1(_1647_),
    .A2(_2650_),
    .Z(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6755_ (.A1(_0969_),
    .A2(_2651_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6756_ (.A1(_2616_),
    .A2(_2629_),
    .B(_2632_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6757_ (.A1(_2652_),
    .A2(_2653_),
    .Z(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6758_ (.A1(_2634_),
    .A2(_2429_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6759_ (.A1(_1910_),
    .A2(_1909_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6760_ (.A1(_2030_),
    .A2(_2656_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6761_ (.A1(_2012_),
    .A2(_2604_),
    .B(_2657_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6762_ (.I0(_2548_),
    .I1(_2658_),
    .S(_2101_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6763_ (.A1(_2324_),
    .A2(_2659_),
    .B(_2210_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6764_ (.A1(_2463_),
    .A2(_2423_),
    .B1(_2655_),
    .B2(_2660_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6765_ (.A1(_2404_),
    .A2(_2654_),
    .B1(_2661_),
    .B2(_2641_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _6766_ (.A1(_2643_),
    .A2(_2648_),
    .A3(_2662_),
    .ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6767_ (.A1(_2623_),
    .A2(_2598_),
    .A3(_2630_),
    .A4(_2652_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6768_ (.A1(_2599_),
    .A2(_2621_),
    .B(_2597_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6769_ (.A1(_0949_),
    .A2(_2629_),
    .B1(_2651_),
    .B2(_2644_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6770_ (.A1(_2644_),
    .A2(_2651_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _6771_ (.A1(_2664_),
    .A2(_2630_),
    .A3(_2652_),
    .B1(_2665_),
    .B2(_2666_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6772_ (.A1(_2561_),
    .A2(_2663_),
    .B(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6773_ (.A1(_1378_),
    .A2(_1557_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6774_ (.A1(_1116_),
    .A2(_1564_),
    .B(_2669_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6775_ (.I(_2670_),
    .Z(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6776_ (.I(_2564_),
    .Z(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6777_ (.A1(_1620_),
    .A2(_1648_),
    .A3(_2626_),
    .Z(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _6778_ (.A1(_1707_),
    .A2(_2486_),
    .A3(_2563_),
    .A4(_2673_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6779_ (.A1(_2672_),
    .A2(_2674_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6780_ (.A1(_2671_),
    .A2(_2675_),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6781_ (.A1(_1849_),
    .A2(_2676_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6782_ (.A1(_2668_),
    .A2(_2677_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6783_ (.A1(_2668_),
    .A2(_2677_),
    .Z(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6784_ (.A1(_2165_),
    .A2(_2678_),
    .A3(_2679_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6785_ (.A1(_1998_),
    .A2(_1113_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6786_ (.I(_2681_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6787_ (.A1(_2182_),
    .A2(_2682_),
    .Z(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6788_ (.I(_1849_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6789_ (.A1(_2684_),
    .A2(_2671_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6790_ (.A1(_2685_),
    .A2(_2578_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6791_ (.A1(_2685_),
    .A2(_2577_),
    .B(_2686_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6792_ (.A1(_2684_),
    .A2(_2671_),
    .B1(_2574_),
    .B2(_2687_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6793_ (.A1(_2289_),
    .A2(_2470_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6794_ (.A1(_0797_),
    .A2(_0971_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6795_ (.I0(_2636_),
    .I1(_2690_),
    .S(_2008_),
    .Z(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6796_ (.I0(_2587_),
    .I1(_2691_),
    .S(_2183_),
    .Z(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6797_ (.A1(_2585_),
    .A2(_2692_),
    .B(_2492_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6798_ (.A1(_2176_),
    .A2(_2140_),
    .A3(_2200_),
    .B1(_2689_),
    .B2(_2693_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6799_ (.A1(_2583_),
    .A2(_2694_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6800_ (.A1(_2680_),
    .A2(_2683_),
    .A3(_2688_),
    .A4(_2695_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6801_ (.I(_2696_),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6802_ (.I(_1847_),
    .Z(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6803_ (.A1(_2671_),
    .A2(_2674_),
    .B(_2672_),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6804_ (.A1(_1848_),
    .A2(_2698_),
    .Z(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6805_ (.A1(_2697_),
    .A2(_2699_),
    .Z(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6806_ (.A1(_2684_),
    .A2(_2676_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6807_ (.A1(_2701_),
    .A2(_2679_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6808_ (.A1(_2700_),
    .A2(_2702_),
    .Z(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6809_ (.I(_2209_),
    .Z(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6810_ (.A1(_2002_),
    .A2(_2503_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6811_ (.I(_2106_),
    .Z(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6812_ (.A1(_2684_),
    .A2(_2706_),
    .B(_1916_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6813_ (.A1(_2122_),
    .A2(_2656_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6814_ (.A1(_2038_),
    .A2(_2707_),
    .B(_2708_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6815_ (.I0(_2606_),
    .I1(_2709_),
    .S(_2101_),
    .Z(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6816_ (.A1(_2061_),
    .A2(_2710_),
    .B(_2026_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6817_ (.A1(_2704_),
    .A2(_2140_),
    .A3(_2224_),
    .B1(_2705_),
    .B2(_2711_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6818_ (.A1(_2697_),
    .A2(_1542_),
    .B(_2374_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6819_ (.A1(_2697_),
    .A2(_1542_),
    .A3(_2373_),
    .B(_2713_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6820_ (.A1(_2697_),
    .A2(_1542_),
    .B1(_2372_),
    .B2(_2714_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6821_ (.A1(_2213_),
    .A2(_2571_),
    .B1(_2712_),
    .B2(_2641_),
    .C(_2715_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6822_ (.A1(_1984_),
    .A2(_2703_),
    .B(_2716_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6823_ (.I(_2717_),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6824_ (.A1(_1849_),
    .A2(_2676_),
    .B1(_2699_),
    .B2(_0829_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6825_ (.A1(_0829_),
    .A2(_2699_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6826_ (.A1(_2668_),
    .A2(_2677_),
    .A3(_2700_),
    .B1(_2718_),
    .B2(_2719_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _6827_ (.A1(_1848_),
    .A2(_2670_),
    .A3(_2674_),
    .B(_2564_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6828_ (.A1(_1853_),
    .A2(_2721_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6829_ (.A1(_1852_),
    .A2(_2722_),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6830_ (.A1(_2720_),
    .A2(_2723_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6831_ (.I(_2404_),
    .Z(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6832_ (.A1(_2720_),
    .A2(_2723_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6833_ (.A1(_2725_),
    .A2(_2726_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6834_ (.A1(_1852_),
    .A2(_2106_),
    .B(_0832_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6835_ (.I0(_2690_),
    .I1(_2728_),
    .S(_2007_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6836_ (.I0(_2637_),
    .I1(_2729_),
    .S(_2040_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6837_ (.A1(_2116_),
    .A2(_2730_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6838_ (.A1(_2634_),
    .A2(_2525_),
    .B(_2210_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6839_ (.A1(_2000_),
    .A2(_2265_),
    .B1(_2731_),
    .B2(_2732_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6840_ (.A1(_0848_),
    .A2(_1853_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6841_ (.A1(_2734_),
    .A2(_2304_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6842_ (.A1(_2734_),
    .A2(_2576_),
    .B(_2735_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6843_ (.A1(_0848_),
    .A2(_1853_),
    .B1(_2345_),
    .B2(_2736_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6844_ (.A1(_2256_),
    .A2(_2682_),
    .B(_2737_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6845_ (.A1(_2583_),
    .A2(_2733_),
    .B(_2738_),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6846_ (.A1(_2724_),
    .A2(_2727_),
    .B(_2739_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6847_ (.I(_2740_),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6848_ (.A1(_1852_),
    .A2(_2722_),
    .Z(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6849_ (.I(_0874_),
    .Z(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6850_ (.A1(_1577_),
    .A2(_2439_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6851_ (.A1(_2743_),
    .A2(_2721_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6852_ (.A1(_1844_),
    .A2(_2744_),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6853_ (.A1(_2742_),
    .A2(_2745_),
    .Z(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6854_ (.A1(_2741_),
    .A2(_2726_),
    .B(_2746_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6855_ (.A1(_2741_),
    .A2(_2726_),
    .A3(_2746_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6856_ (.A1(_2725_),
    .A2(_2748_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6857_ (.A1(_2634_),
    .A2(_2549_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6858_ (.A1(_1843_),
    .A2(_2706_),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6859_ (.A1(_2751_),
    .A2(_1917_),
    .Z(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6860_ (.A1(_2122_),
    .A2(_2707_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6861_ (.A1(_2038_),
    .A2(_2752_),
    .B(_2753_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6862_ (.A1(_2217_),
    .A2(_2658_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6863_ (.A1(_2360_),
    .A2(_2754_),
    .B(_2755_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6864_ (.A1(_2324_),
    .A2(_2756_),
    .B(_2210_),
    .ZN(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6865_ (.A1(_2000_),
    .A2(_2302_),
    .B1(_2750_),
    .B2(_2757_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6866_ (.A1(_2742_),
    .A2(_1844_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6867_ (.A1(_2759_),
    .A2(_2269_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6868_ (.A1(_2759_),
    .A2(_2576_),
    .B(_2760_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6869_ (.A1(_2742_),
    .A2(_1844_),
    .B1(_2345_),
    .B2(_2761_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6870_ (.A1(_2287_),
    .A2(_2682_),
    .B(_2762_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6871_ (.A1(_2583_),
    .A2(_2758_),
    .B(_2763_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6872_ (.A1(_2747_),
    .A2(_2749_),
    .B(_2764_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6873_ (.I(_2765_),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6874_ (.A1(_1555_),
    .A2(_2672_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6875_ (.A1(_2721_),
    .A2(_2743_),
    .A3(_2766_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6876_ (.A1(_1459_),
    .A2(_2767_),
    .Z(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6877_ (.A1(_1057_),
    .A2(_2768_),
    .Z(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6878_ (.A1(_1820_),
    .A2(_2488_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6879_ (.A1(_2444_),
    .A2(_2450_),
    .B(_2516_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6880_ (.A1(_2533_),
    .A2(_2513_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6881_ (.A1(_2533_),
    .A2(_2514_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6882_ (.A1(_2770_),
    .A2(_2771_),
    .A3(_2772_),
    .B(_2773_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6883_ (.A1(_1838_),
    .A2(_2539_),
    .Z(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6884_ (.A1(_1838_),
    .A2(_2540_),
    .Z(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6885_ (.A1(_2774_),
    .A2(_2775_),
    .B(_2776_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6886_ (.I(_2723_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6887_ (.A1(_2677_),
    .A2(_2700_),
    .A3(_2778_),
    .A4(_2746_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6888_ (.A1(_2663_),
    .A2(_2779_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6889_ (.A1(_2719_),
    .A2(_2718_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6890_ (.A1(_2778_),
    .A2(_2746_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6891_ (.A1(_1843_),
    .A2(_2745_),
    .B(_2741_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6892_ (.A1(_1843_),
    .A2(_2745_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _6893_ (.A1(_2781_),
    .A2(_2782_),
    .B1(_2783_),
    .B2(_2784_),
    .C1(_2779_),
    .C2(_2667_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6894_ (.A1(_2777_),
    .A2(_2780_),
    .B(_2785_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6895_ (.A1(_2769_),
    .A2(_2786_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6896_ (.A1(_2742_),
    .A2(_2706_),
    .B(_1059_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6897_ (.A1(_2012_),
    .A2(_2788_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6898_ (.A1(_2029_),
    .A2(_2728_),
    .B(_2789_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6899_ (.A1(_2362_),
    .A2(_2790_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6900_ (.A1(_2245_),
    .A2(_2691_),
    .B(_2791_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6901_ (.A1(_2137_),
    .A2(_2588_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6902_ (.A1(_2585_),
    .A2(_2792_),
    .B(_2793_),
    .C(_2492_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6903_ (.A1(_2284_),
    .A2(_2341_),
    .B(_2794_),
    .C(_2610_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6904_ (.A1(_2061_),
    .A2(_2681_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6905_ (.A1(_1379_),
    .A2(_1881_),
    .B(_1882_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6906_ (.I(_1057_),
    .Z(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6907_ (.A1(_2797_),
    .A2(_2798_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6908_ (.A1(_2799_),
    .A2(_2496_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6909_ (.A1(_2799_),
    .A2(_2168_),
    .B(_2800_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6910_ (.A1(_2797_),
    .A2(_2798_),
    .B1(_2266_),
    .B2(_2801_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6911_ (.A1(_1983_),
    .A2(_2802_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6912_ (.A1(_1104_),
    .A2(_2796_),
    .B(_2803_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _6913_ (.A1(_2725_),
    .A2(_2787_),
    .B1(_2795_),
    .B2(_2804_),
    .ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6914_ (.A1(_2798_),
    .A2(_2768_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6915_ (.A1(_2769_),
    .A2(_2786_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6916_ (.I(_1879_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6917_ (.A1(_2797_),
    .A2(_2767_),
    .B(_2484_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6918_ (.A1(_2807_),
    .A2(_2808_),
    .Z(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6919_ (.A1(_1878_),
    .A2(_2809_),
    .Z(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6920_ (.A1(_1878_),
    .A2(_2809_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6921_ (.A1(_2810_),
    .A2(_2811_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6922_ (.A1(_2805_),
    .A2(_2806_),
    .B(_2812_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6923_ (.A1(_2805_),
    .A2(_2806_),
    .A3(_2812_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6924_ (.A1(_2404_),
    .A2(_2814_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6925_ (.A1(_1071_),
    .A2(_2363_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6926_ (.A1(_2798_),
    .A2(_2107_),
    .B(_2816_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6927_ (.A1(_2038_),
    .A2(_2752_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6928_ (.A1(_2036_),
    .A2(_2817_),
    .B(_2818_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6929_ (.A1(_2217_),
    .A2(_2709_),
    .Z(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6930_ (.A1(_2246_),
    .A2(_2819_),
    .B(_2820_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6931_ (.A1(_2137_),
    .A2(_2607_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6932_ (.A1(_2585_),
    .A2(_2821_),
    .B(_2822_),
    .C(_2326_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6933_ (.A1(_2421_),
    .A2(_2370_),
    .B(_2823_),
    .C(_2582_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6934_ (.I0(_2269_),
    .I1(_2080_),
    .S(_1399_),
    .Z(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6935_ (.A1(_1878_),
    .A2(_2807_),
    .B1(_2074_),
    .B2(_2825_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6936_ (.I(_2826_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6937_ (.A1(_1934_),
    .A2(_2796_),
    .B(_2827_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6938_ (.A1(_2813_),
    .A2(_2815_),
    .B(_2824_),
    .C(_2828_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _6939_ (.I(_2829_),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6940_ (.A1(_2769_),
    .A2(_2810_),
    .A3(_2811_),
    .Z(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6941_ (.A1(_2805_),
    .A2(_2811_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6942_ (.A1(_2810_),
    .A2(_2831_),
    .Z(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6943_ (.A1(_2786_),
    .A2(_2830_),
    .B(_2832_),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6944_ (.I(_1376_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6945_ (.A1(_2807_),
    .A2(_2797_),
    .B(_2672_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _6946_ (.A1(_2721_),
    .A2(_2743_),
    .A3(_2766_),
    .A4(_2835_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6947_ (.A1(_2834_),
    .A2(_2836_),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6948_ (.A1(_1085_),
    .A2(_2837_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6949_ (.A1(_2833_),
    .A2(_2838_),
    .Z(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6950_ (.A1(_2833_),
    .A2(_2838_),
    .B(_2351_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6951_ (.I(_1085_),
    .Z(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6952_ (.A1(_2841_),
    .A2(_2142_),
    .B(_1072_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6953_ (.I0(_2788_),
    .I1(_2842_),
    .S(_2105_),
    .Z(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6954_ (.A1(_2010_),
    .A2(_2729_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6955_ (.A1(_2005_),
    .A2(_2843_),
    .B(_2844_),
    .C(_2214_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6956_ (.A1(_2424_),
    .A2(_2638_),
    .B(_2845_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6957_ (.A1(_2189_),
    .A2(_2386_),
    .B(_2067_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6958_ (.A1(_2176_),
    .A2(_2846_),
    .B(_2847_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6959_ (.A1(_2333_),
    .A2(_2570_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6960_ (.A1(_2841_),
    .A2(_2834_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6961_ (.A1(_2850_),
    .A2(_2496_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6962_ (.A1(_2850_),
    .A2(_2168_),
    .B(_2851_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6963_ (.A1(_2841_),
    .A2(_2834_),
    .B1(_2074_),
    .B2(_2852_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6964_ (.A1(_2015_),
    .A2(_2849_),
    .B(_2853_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6965_ (.A1(_2839_),
    .A2(_2840_),
    .B(_2848_),
    .C(_2854_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _6966_ (.I(_2855_),
    .ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6967_ (.I(_1441_),
    .Z(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6968_ (.A1(_2834_),
    .A2(_2484_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6969_ (.A1(_2836_),
    .A2(_2857_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6970_ (.A1(_2856_),
    .A2(_2858_),
    .Z(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6971_ (.A1(_1099_),
    .A2(_2859_),
    .Z(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6972_ (.A1(_2841_),
    .A2(_2837_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6973_ (.A1(_2861_),
    .A2(_2839_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6974_ (.A1(_2860_),
    .A2(_2862_),
    .Z(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6975_ (.A1(_1927_),
    .A2(_1930_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6976_ (.A1(_2008_),
    .A2(_2864_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6977_ (.A1(_2030_),
    .A2(_2817_),
    .B(_2865_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6978_ (.A1(_2005_),
    .A2(_2754_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6979_ (.A1(_2064_),
    .A2(_2866_),
    .B(_2867_),
    .C(_2017_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6980_ (.A1(_2177_),
    .A2(_2659_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6981_ (.A1(_2704_),
    .A2(_2868_),
    .A3(_2869_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6982_ (.A1(_2421_),
    .A2(_2431_),
    .B(_2870_),
    .C(_2582_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6983_ (.A1(_1099_),
    .A2(_2856_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6984_ (.A1(_2872_),
    .A2(_2077_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6985_ (.A1(_2872_),
    .A2(_2373_),
    .B(_2873_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6986_ (.A1(_1099_),
    .A2(_2856_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6987_ (.A1(_2174_),
    .A2(_2874_),
    .B(_2875_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6988_ (.A1(_2113_),
    .A2(_2796_),
    .B(_2876_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6989_ (.A1(_2352_),
    .A2(_2863_),
    .B(_2871_),
    .C(_2877_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6990_ (.I(_2878_),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6991_ (.I(_0997_),
    .Z(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6992_ (.A1(_2856_),
    .A2(_2484_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6993_ (.A1(_2836_),
    .A2(_2857_),
    .A3(_2880_),
    .Z(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6994_ (.A1(_1521_),
    .A2(_2881_),
    .Z(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6995_ (.A1(_2879_),
    .A2(_2882_),
    .Z(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6996_ (.A1(_2879_),
    .A2(_2882_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6997_ (.A1(_2883_),
    .A2(_2884_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6998_ (.A1(_2860_),
    .A2(_2838_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6999_ (.A1(_1409_),
    .A2(_2859_),
    .B(_2861_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7000_ (.A1(_1409_),
    .A2(_2859_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7001_ (.A1(_2830_),
    .A2(_2886_),
    .Z(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _7002_ (.A1(_2832_),
    .A2(net235),
    .B1(_2887_),
    .B2(_2888_),
    .C1(_2889_),
    .C2(_2786_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7003_ (.A1(_2885_),
    .A2(_2890_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7004_ (.A1(_2061_),
    .A2(_2692_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7005_ (.A1(_2879_),
    .A2(_2706_),
    .B(_1100_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7006_ (.A1(_2117_),
    .A2(_2893_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7007_ (.A1(_2117_),
    .A2(_2842_),
    .B(_2894_),
    .C(_2362_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7008_ (.A1(_2360_),
    .A2(_2790_),
    .ZN(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7009_ (.A1(_2333_),
    .A2(_2895_),
    .A3(_2896_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7010_ (.A1(_2704_),
    .A2(_2892_),
    .A3(_2897_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7011_ (.A1(_2284_),
    .A2(_2472_),
    .B(_2898_),
    .C(_2610_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7012_ (.A1(_0996_),
    .A2(_1890_),
    .B(_2374_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7013_ (.A1(_2879_),
    .A2(_1521_),
    .A3(_2168_),
    .B(_2173_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7014_ (.A1(_0996_),
    .A2(_1890_),
    .B1(_2900_),
    .B2(_2901_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7015_ (.A1(_2180_),
    .A2(_2849_),
    .B(_2902_),
    .C(_2351_),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7016_ (.I(_2903_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7017_ (.A1(_2725_),
    .A2(_2891_),
    .B1(_2899_),
    .B2(_2904_),
    .ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7018_ (.I(_1010_),
    .Z(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7019_ (.I(_2905_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7020_ (.A1(_1521_),
    .A2(_2537_),
    .B(_2881_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7021_ (.A1(_1508_),
    .A2(_2907_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7022_ (.A1(_2906_),
    .A2(_2908_),
    .Z(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7023_ (.A1(_2885_),
    .A2(_2890_),
    .B(_2883_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7024_ (.A1(_2909_),
    .A2(_2910_),
    .Z(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7025_ (.I(_1508_),
    .Z(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7026_ (.A1(_2906_),
    .A2(_2912_),
    .B(_2076_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7027_ (.A1(_2906_),
    .A2(_2912_),
    .A3(_2081_),
    .B(_2913_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7028_ (.A1(_2906_),
    .A2(_2912_),
    .B1(_2174_),
    .B2(_2914_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7029_ (.A1(_2212_),
    .A2(_2796_),
    .B(_2915_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7030_ (.A1(_2036_),
    .A2(_2864_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7031_ (.A1(_1929_),
    .A2(_1922_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7032_ (.A1(_2029_),
    .A2(_2918_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7033_ (.A1(_2362_),
    .A2(_2917_),
    .A3(_2919_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7034_ (.A1(_2245_),
    .A2(_2819_),
    .B(_2920_),
    .C(_2424_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7035_ (.A1(_2135_),
    .A2(_2710_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7036_ (.A1(_2704_),
    .A2(_2921_),
    .A3(_2922_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7037_ (.A1(_2421_),
    .A2(_2505_),
    .B(_2923_),
    .C(_2610_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7038_ (.A1(_2352_),
    .A2(_2911_),
    .B(_2916_),
    .C(_2924_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7039_ (.I(_2925_),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7040_ (.I(_1041_),
    .Z(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7041_ (.A1(_2912_),
    .A2(_2537_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7042_ (.A1(_2907_),
    .A2(_2927_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7043_ (.A1(_1874_),
    .A2(_2928_),
    .Z(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7044_ (.A1(_2926_),
    .A2(_2929_),
    .Z(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7045_ (.A1(_2905_),
    .A2(_2908_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7046_ (.A1(_2883_),
    .A2(_2931_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7047_ (.A1(_2905_),
    .A2(_2908_),
    .B(_2932_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7048_ (.A1(_2885_),
    .A2(_2890_),
    .A3(_2909_),
    .B(_2933_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7049_ (.A1(_2930_),
    .A2(net214),
    .B(_2086_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7050_ (.A1(_2930_),
    .A2(_2934_),
    .B(_2935_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7051_ (.A1(_2926_),
    .A2(_1874_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7052_ (.A1(_2937_),
    .A2(_2304_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7053_ (.A1(_2937_),
    .A2(_2576_),
    .B(_2938_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7054_ (.A1(_2926_),
    .A2(_1874_),
    .B1(_2075_),
    .B2(_2939_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7055_ (.A1(_2010_),
    .A2(_2843_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7056_ (.A1(_2905_),
    .A2(_2107_),
    .B(_2030_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7057_ (.A1(_2122_),
    .A2(_2893_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7058_ (.A1(_1043_),
    .A2(_2942_),
    .B(_2943_),
    .C(_2120_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7059_ (.A1(_2941_),
    .A2(_2944_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7060_ (.A1(_2139_),
    .A2(_2730_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7061_ (.A1(_2046_),
    .A2(_2945_),
    .B(_2946_),
    .C(_1999_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7062_ (.A1(_2492_),
    .A2(_2526_),
    .B(_2947_),
    .C(_2582_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7063_ (.A1(_2254_),
    .A2(_2849_),
    .B(_2940_),
    .C(_2948_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7064_ (.A1(_2936_),
    .A2(_2949_),
    .Z(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _7065_ (.I(_2950_),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7066_ (.A1(_2926_),
    .A2(_2929_),
    .B1(_2930_),
    .B2(_2934_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7067_ (.A1(_1495_),
    .A2(_2928_),
    .B(_2537_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7068_ (.A1(_1873_),
    .A2(_2951_),
    .A3(_2952_),
    .Z(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7069_ (.A1(_2194_),
    .A2(_1921_),
    .B(_2108_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7070_ (.A1(_2036_),
    .A2(_2918_),
    .B(_2954_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7071_ (.A1(_2217_),
    .A2(_2866_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7072_ (.A1(_2360_),
    .A2(_2955_),
    .B(_2956_),
    .C(_2027_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7073_ (.A1(_2002_),
    .A2(_2756_),
    .B(_2957_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7074_ (.A1(_2257_),
    .A2(_2550_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7075_ (.A1(_2257_),
    .A2(_2958_),
    .B(_2959_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7076_ (.A1(_2103_),
    .A2(_1477_),
    .ZN(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7077_ (.A1(_2961_),
    .A2(_2171_),
    .B(_2074_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7078_ (.A1(_2103_),
    .A2(_1477_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _7079_ (.A1(_2961_),
    .A2(_2169_),
    .B1(_2542_),
    .B2(_2682_),
    .C1(_2962_),
    .C2(_2963_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7080_ (.A1(_2641_),
    .A2(_2960_),
    .B(_2964_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7081_ (.A1(_2352_),
    .A2(_2953_),
    .B(_2965_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7082_ (.I(_2966_),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7083_ (.I(_1709_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7084_ (.I(_2967_),
    .Z(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7085_ (.I(_0727_),
    .Z(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7086_ (.I(_2969_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7087_ (.I(_2970_),
    .Z(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7088_ (.I(net4),
    .Z(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7089_ (.A1(_2968_),
    .A2(_2971_),
    .A3(_2972_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7090_ (.A1(net97),
    .A2(_2973_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7091_ (.I(_0705_),
    .Z(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7092_ (.A1(_1709_),
    .A2(_0714_),
    .A3(_2975_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7093_ (.I(_2976_),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7094_ (.I(_2977_),
    .Z(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7095_ (.I(_2978_),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7096_ (.I(_2979_),
    .Z(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7097_ (.A1(net108),
    .A2(_2974_),
    .B(_2980_),
    .ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7098_ (.A1(_2969_),
    .A2(_2972_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7099_ (.A1(net6),
    .A2(_2981_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7100_ (.A1(net97),
    .A2(_2982_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7101_ (.A1(net108),
    .A2(_2983_),
    .B(_2980_),
    .ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7102_ (.I(_1982_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7103_ (.A1(_2984_),
    .A2(_2974_),
    .B(_2980_),
    .ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7104_ (.A1(_2984_),
    .A2(_2983_),
    .B(_2980_),
    .ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7105_ (.A1(net6),
    .A2(_2970_),
    .A3(_2972_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7106_ (.A1(_2985_),
    .A2(_2982_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7107_ (.I(_2986_),
    .Z(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7108_ (.I(_2987_),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7109_ (.I(_2988_),
    .Z(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7110_ (.A1(net134),
    .A2(_2988_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7111_ (.A1(net212),
    .A2(_2989_),
    .B(_2990_),
    .ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7112_ (.A1(net145),
    .A2(_2988_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7113_ (.A1(_1828_),
    .A2(_2989_),
    .B(_2991_),
    .ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7114_ (.I(_2987_),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7115_ (.A1(net156),
    .A2(_2992_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7116_ (.A1(_1679_),
    .A2(_2989_),
    .B(_2993_),
    .ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7117_ (.A1(net159),
    .A2(_2992_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7118_ (.A1(_1664_),
    .A2(_2989_),
    .B(_2994_),
    .ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7119_ (.I(_2988_),
    .Z(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7120_ (.A1(net160),
    .A2(_2992_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7121_ (.A1(_1690_),
    .A2(_2995_),
    .B(_2996_),
    .ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7122_ (.A1(net161),
    .A2(_2992_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7123_ (.A1(_1702_),
    .A2(_2995_),
    .B(_2997_),
    .ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7124_ (.A1(net162),
    .A2(_2987_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7125_ (.A1(_1717_),
    .A2(_2995_),
    .B(_2998_),
    .ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7126_ (.A1(net163),
    .A2(_2987_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7127_ (.A1(_1729_),
    .A2(_2995_),
    .B(_2999_),
    .ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7128_ (.I(_2979_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7129_ (.I(_2978_),
    .Z(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7130_ (.I(_3001_),
    .Z(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7131_ (.A1(net134),
    .A2(_3002_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7132_ (.A1(net228),
    .A2(_3000_),
    .B(_3003_),
    .ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7133_ (.I(_3001_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7134_ (.A1(net145),
    .A2(_3004_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7135_ (.A1(net225),
    .A2(_3000_),
    .B(_3005_),
    .ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7136_ (.I(_0494_),
    .Z(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7137_ (.A1(_3006_),
    .A2(net222),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7138_ (.A1(net156),
    .A2(_3004_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7139_ (.A1(_3007_),
    .A2(_3000_),
    .B(_3008_),
    .ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7140_ (.A1(net159),
    .A2(_3004_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7141_ (.A1(_1645_),
    .A2(_3000_),
    .B(_3009_),
    .ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7142_ (.I(_2985_),
    .Z(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7143_ (.A1(_3006_),
    .A2(_1563_),
    .A3(_3010_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7144_ (.A1(_0555_),
    .A2(_3010_),
    .B(_3011_),
    .ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7145_ (.I(_3001_),
    .Z(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7146_ (.A1(net161),
    .A2(_3004_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7147_ (.A1(_1539_),
    .A2(_3012_),
    .B(_3013_),
    .ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7148_ (.A1(_3006_),
    .A2(_1575_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7149_ (.A1(net162),
    .A2(_2979_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7150_ (.A1(_3014_),
    .A2(_3012_),
    .B(_3015_),
    .ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7151_ (.A1(net163),
    .A2(_2979_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7152_ (.A1(_1552_),
    .A2(_3012_),
    .B(_3016_),
    .ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7153_ (.I(_2973_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7154_ (.A1(_1457_),
    .A2(_3012_),
    .B1(_3017_),
    .B2(net212),
    .C(_2990_),
    .ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7155_ (.I(_3001_),
    .Z(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7156_ (.A1(_1397_),
    .A2(_3018_),
    .B1(_3017_),
    .B2(_1828_),
    .C(_2991_),
    .ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7157_ (.A1(_1374_),
    .A2(_3018_),
    .B1(_3017_),
    .B2(_1679_),
    .C(_2993_),
    .ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7158_ (.A1(_3006_),
    .A2(net219),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7159_ (.A1(_3019_),
    .A2(_3018_),
    .B1(_3017_),
    .B2(_1664_),
    .C(_2994_),
    .ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7160_ (.I(_2973_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7161_ (.A1(net234),
    .A2(_3018_),
    .B1(_3020_),
    .B2(_1690_),
    .C(_2996_),
    .ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7162_ (.A1(net223),
    .A2(_3002_),
    .B1(_3020_),
    .B2(_1702_),
    .C(_2997_),
    .ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7163_ (.A1(net220),
    .A2(_3002_),
    .B1(_3020_),
    .B2(_1717_),
    .C(_2998_),
    .ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7164_ (.A1(_1475_),
    .A2(_3002_),
    .B1(_3020_),
    .B2(_1729_),
    .C(_2999_),
    .ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7165_ (.A1(_2970_),
    .A2(_1981_),
    .Z(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7166_ (.I(_3021_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7167_ (.I(_3022_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7168_ (.I(_3023_),
    .Z(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7169_ (.A1(_2969_),
    .A2(_2975_),
    .A3(_1900_),
    .Z(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7170_ (.I(_3025_),
    .Z(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7171_ (.I(_3026_),
    .Z(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7172_ (.I(_3027_),
    .Z(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7173_ (.I(_3028_),
    .Z(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7174_ (.A1(_3024_),
    .A2(_3029_),
    .ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7175_ (.A1(_2972_),
    .A2(net97),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7176_ (.A1(net108),
    .A2(_3030_),
    .B(_2971_),
    .ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7177_ (.A1(_2975_),
    .A2(_1901_),
    .ZN(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7178_ (.I(_3031_),
    .Z(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7179_ (.A1(_1982_),
    .A2(_3032_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7180_ (.A1(_2971_),
    .A2(_3033_),
    .ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7181_ (.A1(_2984_),
    .A2(_3030_),
    .B(_2971_),
    .ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7182_ (.I(_0746_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _7183_ (.A1(_0663_),
    .A2(_3034_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7184_ (.I(_2975_),
    .Z(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7185_ (.A1(_3036_),
    .A2(_1901_),
    .Z(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7186_ (.A1(_0701_),
    .A2(_3037_),
    .B(_1410_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7187_ (.I(_3038_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7188_ (.A1(_3035_),
    .A2(_3039_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7189_ (.I(_3040_),
    .Z(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7190_ (.I(_3041_),
    .Z(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7191_ (.A1(net65),
    .A2(_0689_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7192_ (.I(_3039_),
    .Z(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7193_ (.I(_3044_),
    .Z(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7194_ (.I(_3045_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7195_ (.A1(_0606_),
    .A2(_3042_),
    .B1(_3043_),
    .B2(_3046_),
    .ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7196_ (.I(_0613_),
    .Z(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7197_ (.I(_3047_),
    .Z(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7198_ (.A1(_0608_),
    .A2(_3048_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7199_ (.I(_3049_),
    .Z(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7200_ (.I(_3050_),
    .Z(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7201_ (.I(_3038_),
    .Z(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7202_ (.I(_3052_),
    .Z(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7203_ (.A1(net65),
    .A2(_0689_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7204_ (.A1(_1324_),
    .A2(_1180_),
    .Z(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7205_ (.A1(_3054_),
    .A2(_3055_),
    .Z(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7206_ (.A1(_3051_),
    .A2(_1982_),
    .B1(_3053_),
    .B2(_3056_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7207_ (.A1(_1324_),
    .A2(_3042_),
    .B(_3057_),
    .ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7208_ (.I(net87),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7209_ (.I(_3050_),
    .Z(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7210_ (.I(_3052_),
    .Z(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7211_ (.I(_3060_),
    .Z(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7212_ (.A1(net76),
    .A2(_1180_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7213_ (.A1(_3054_),
    .A2(_3055_),
    .B(_3062_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7214_ (.A1(_3058_),
    .A2(_1238_),
    .A3(_3063_),
    .Z(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7215_ (.A1(_3059_),
    .A2(net119),
    .B1(_3061_),
    .B2(_3064_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7216_ (.A1(_3058_),
    .A2(_3042_),
    .B(_3065_),
    .ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7217_ (.I(_1300_),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7218_ (.I(net90),
    .Z(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7219_ (.A1(_3066_),
    .A2(_3067_),
    .Z(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7220_ (.I(_1108_),
    .Z(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7221_ (.A1(_3066_),
    .A2(_0977_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7222_ (.A1(_3066_),
    .A2(_0977_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7223_ (.A1(_3070_),
    .A2(_3063_),
    .B(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7224_ (.A1(_3067_),
    .A2(_3069_),
    .A3(_3072_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7225_ (.A1(_3059_),
    .A2(net122),
    .B1(_3061_),
    .B2(_3073_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7226_ (.A1(_3042_),
    .A2(_3068_),
    .B(_3074_),
    .ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7227_ (.I(_3040_),
    .Z(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7228_ (.I(_3075_),
    .Z(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7229_ (.I(_3076_),
    .Z(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7230_ (.I(net91),
    .Z(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7231_ (.A1(_3058_),
    .A2(_3067_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7232_ (.A1(_3078_),
    .A2(_3079_),
    .Z(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7233_ (.I(_0741_),
    .Z(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7234_ (.A1(net90),
    .A2(_3069_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7235_ (.A1(_3067_),
    .A2(_3069_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7236_ (.A1(_3082_),
    .A2(_3072_),
    .B(_3083_),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7237_ (.A1(_3078_),
    .A2(_3081_),
    .A3(_3084_),
    .Z(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7238_ (.A1(_3059_),
    .A2(net123),
    .B1(_3061_),
    .B2(_3085_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7239_ (.A1(_3077_),
    .A2(_3080_),
    .B(_3086_),
    .ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7240_ (.I(net92),
    .Z(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7241_ (.A1(_3058_),
    .A2(net90),
    .A3(net91),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7242_ (.A1(_3087_),
    .A2(_3088_),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7243_ (.A1(_1382_),
    .A2(_1383_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7244_ (.A1(_3078_),
    .A2(_3081_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7245_ (.A1(_3078_),
    .A2(_3081_),
    .Z(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7246_ (.A1(_3092_),
    .A2(_3084_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7247_ (.A1(_3091_),
    .A2(_3093_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7248_ (.A1(_3087_),
    .A2(_3090_),
    .A3(_3094_),
    .Z(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7249_ (.A1(_3059_),
    .A2(net124),
    .B1(_3061_),
    .B2(_3095_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7250_ (.A1(_3077_),
    .A2(_3089_),
    .B(_3096_),
    .ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7251_ (.I(net93),
    .Z(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7252_ (.A1(_1270_),
    .A2(_3088_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7253_ (.A1(_3097_),
    .A2(_3098_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7254_ (.I(_3050_),
    .Z(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7255_ (.I(_3052_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7256_ (.A1(_2229_),
    .A2(_1383_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7257_ (.A1(net93),
    .A2(_3102_),
    .Z(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7258_ (.I(_3103_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7259_ (.A1(_3087_),
    .A2(_3090_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7260_ (.A1(_3087_),
    .A2(_3090_),
    .ZN(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7261_ (.A1(_3091_),
    .A2(_3106_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7262_ (.A1(_3092_),
    .A2(_3084_),
    .B(_3107_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7263_ (.A1(_3105_),
    .A2(_3108_),
    .Z(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7264_ (.A1(_3104_),
    .A2(_3109_),
    .Z(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7265_ (.A1(_3100_),
    .A2(net125),
    .B1(_3101_),
    .B2(_3110_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7266_ (.A1(_3077_),
    .A2(_3099_),
    .B(_3111_),
    .ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7267_ (.A1(net93),
    .A2(net94),
    .A3(_3098_),
    .Z(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7268_ (.I(net94),
    .Z(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7269_ (.A1(_3097_),
    .A2(_3098_),
    .B(_3113_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7270_ (.A1(_3112_),
    .A2(_3114_),
    .Z(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _7271_ (.A1(_1769_),
    .A2(_1383_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7272_ (.A1(_3097_),
    .A2(_3102_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7273_ (.A1(_3104_),
    .A2(_3109_),
    .B(_3117_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7274_ (.A1(_3113_),
    .A2(_3116_),
    .A3(_3118_),
    .Z(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7275_ (.A1(_3100_),
    .A2(net126),
    .B1(_3101_),
    .B2(_3119_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7276_ (.A1(_3077_),
    .A2(_3115_),
    .B(_3120_),
    .ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7277_ (.I(_3076_),
    .Z(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7278_ (.I(net95),
    .Z(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7279_ (.A1(_3122_),
    .A2(_3112_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7280_ (.A1(_3113_),
    .A2(_3116_),
    .Z(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7281_ (.A1(_3113_),
    .A2(_3116_),
    .B1(_3102_),
    .B2(_3097_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7282_ (.A1(_3105_),
    .A2(_3104_),
    .A3(_3108_),
    .B(_3125_),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7283_ (.A1(_3124_),
    .A2(_3126_),
    .Z(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7284_ (.A1(net21),
    .A2(_1443_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7285_ (.A1(_3122_),
    .A2(_3128_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7286_ (.A1(_3127_),
    .A2(_3129_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7287_ (.A1(_3100_),
    .A2(net127),
    .B1(_3101_),
    .B2(_3130_),
    .ZN(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7288_ (.A1(_3121_),
    .A2(_3123_),
    .B(_3131_),
    .ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7289_ (.A1(net95),
    .A2(net96),
    .A3(_3112_),
    .Z(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7290_ (.I(_3132_),
    .Z(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7291_ (.I(net96),
    .Z(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7292_ (.A1(_3122_),
    .A2(_3112_),
    .B(_3134_),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7293_ (.A1(_3133_),
    .A2(_3135_),
    .Z(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7294_ (.A1(_3134_),
    .A2(_1829_),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7295_ (.I(_1443_),
    .Z(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7296_ (.A1(_3122_),
    .A2(net21),
    .A3(_3138_),
    .ZN(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7297_ (.A1(_3127_),
    .A2(_3129_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7298_ (.A1(_3139_),
    .A2(_3140_),
    .Z(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7299_ (.A1(_3137_),
    .A2(_3141_),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7300_ (.A1(_3100_),
    .A2(net128),
    .B1(_3101_),
    .B2(_3142_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7301_ (.A1(_3121_),
    .A2(_3136_),
    .B(_3143_),
    .ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7302_ (.I(_3075_),
    .Z(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7303_ (.I(net66),
    .Z(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7304_ (.A1(_3145_),
    .A2(_3133_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7305_ (.A1(_3134_),
    .A2(net22),
    .A3(_3138_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7306_ (.A1(net22),
    .A2(_1443_),
    .B(_3134_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7307_ (.A1(_3147_),
    .A2(_3141_),
    .B(_3148_),
    .ZN(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7308_ (.A1(net66),
    .A2(_1671_),
    .Z(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7309_ (.A1(_3149_),
    .A2(_3150_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7310_ (.A1(_3149_),
    .A2(_3150_),
    .Z(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7311_ (.A1(_3060_),
    .A2(_3151_),
    .A3(_3152_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7312_ (.A1(_3035_),
    .A2(_2413_),
    .B1(_3144_),
    .B2(_3146_),
    .C(_3153_),
    .ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7313_ (.I(net67),
    .Z(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7314_ (.A1(_3145_),
    .A2(_3133_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7315_ (.A1(_3154_),
    .A2(_3155_),
    .Z(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7316_ (.I(_3050_),
    .Z(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7317_ (.I(_3052_),
    .Z(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7318_ (.A1(_3145_),
    .A2(_1671_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7319_ (.A1(_3159_),
    .A2(_3151_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7320_ (.I(_1656_),
    .Z(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7321_ (.A1(net67),
    .A2(_3161_),
    .Z(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7322_ (.A1(_3160_),
    .A2(_3162_),
    .Z(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7323_ (.A1(_3157_),
    .A2(net99),
    .B1(_3158_),
    .B2(_3163_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7324_ (.A1(_3121_),
    .A2(_3156_),
    .B(_3164_),
    .ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7325_ (.I(net68),
    .Z(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7326_ (.A1(_3145_),
    .A2(_3154_),
    .A3(_3133_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7327_ (.A1(_3165_),
    .A2(_3166_),
    .Z(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7328_ (.A1(_3165_),
    .A2(_1692_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7329_ (.A1(_3150_),
    .A2(_3162_),
    .ZN(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7330_ (.A1(_3139_),
    .A2(_3147_),
    .B(_3169_),
    .C(_3148_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7331_ (.A1(_3154_),
    .A2(_3161_),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7332_ (.A1(_3159_),
    .A2(_3171_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7333_ (.A1(_3154_),
    .A2(_3161_),
    .B(_3170_),
    .C(_3172_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7334_ (.A1(_3137_),
    .A2(_3169_),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _7335_ (.A1(_3124_),
    .A2(_3126_),
    .A3(_3129_),
    .A4(_3174_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7336_ (.A1(_3173_),
    .A2(_3175_),
    .Z(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7337_ (.A1(_3168_),
    .A2(_3176_),
    .Z(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7338_ (.A1(_3157_),
    .A2(net100),
    .B1(_3158_),
    .B2(_3177_),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7339_ (.A1(_3121_),
    .A2(_3167_),
    .B(_3178_),
    .ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7340_ (.I(_3041_),
    .Z(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7341_ (.I(net69),
    .Z(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7342_ (.A1(net66),
    .A2(net67),
    .A3(_3165_),
    .A4(_3132_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7343_ (.A1(_3180_),
    .A2(_3181_),
    .Z(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7344_ (.A1(_2969_),
    .A2(_1704_),
    .B(_1705_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7345_ (.I(_3183_),
    .Z(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7346_ (.A1(_3180_),
    .A2(_3184_),
    .Z(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7347_ (.A1(net69),
    .A2(_3183_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7348_ (.A1(_3185_),
    .A2(_3186_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7349_ (.A1(_3165_),
    .A2(_1692_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7350_ (.A1(_3168_),
    .A2(_3176_),
    .B(_3188_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7351_ (.A1(_3187_),
    .A2(_3189_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7352_ (.A1(_3157_),
    .A2(net101),
    .B1(_3158_),
    .B2(_3190_),
    .ZN(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7353_ (.A1(_3179_),
    .A2(_3182_),
    .B(_3191_),
    .ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7354_ (.I(net70),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7355_ (.A1(_1134_),
    .A2(_3181_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7356_ (.A1(_3192_),
    .A2(_3193_),
    .ZN(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7357_ (.A1(_3180_),
    .A2(_3184_),
    .Z(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7358_ (.A1(_3195_),
    .A2(_3189_),
    .B(_3185_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7359_ (.A1(_3192_),
    .A2(_1710_),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7360_ (.A1(_3196_),
    .A2(_3197_),
    .Z(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7361_ (.A1(_3157_),
    .A2(net102),
    .B1(_3158_),
    .B2(_3198_),
    .ZN(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7362_ (.A1(_3179_),
    .A2(_3194_),
    .B(_3199_),
    .ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7363_ (.I(_3075_),
    .Z(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7364_ (.A1(_3192_),
    .A2(_3193_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7365_ (.A1(net71),
    .A2(_3201_),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7366_ (.A1(_3192_),
    .A2(_1710_),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7367_ (.A1(_3196_),
    .A2(_3197_),
    .B(_3203_),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7368_ (.I(_1722_),
    .Z(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7369_ (.A1(_1165_),
    .A2(_3205_),
    .Z(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7370_ (.A1(_3204_),
    .A2(_3206_),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7371_ (.I(_3049_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7372_ (.I(_3208_),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7373_ (.A1(_3209_),
    .A2(net103),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7374_ (.A1(_3200_),
    .A2(_3202_),
    .B1(_3207_),
    .B2(_3046_),
    .C(_3210_),
    .ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7375_ (.A1(_1165_),
    .A2(_3201_),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7376_ (.A1(_0911_),
    .A2(_3211_),
    .Z(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7377_ (.A1(_0911_),
    .A2(_1585_),
    .Z(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7378_ (.A1(net71),
    .A2(_3205_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7379_ (.A1(_3197_),
    .A2(_3206_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7380_ (.A1(_3180_),
    .A2(_3184_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7381_ (.A1(_3188_),
    .A2(_3216_),
    .B(_3186_),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7382_ (.A1(_3215_),
    .A2(_3217_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7383_ (.A1(net71),
    .A2(_3205_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7384_ (.A1(_3203_),
    .A2(_3214_),
    .B(_3218_),
    .C(_3219_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7385_ (.A1(_3185_),
    .A2(_3186_),
    .A3(_3215_),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7386_ (.A1(_3173_),
    .A2(_3175_),
    .B(_3221_),
    .C(_3168_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7387_ (.A1(_3220_),
    .A2(_3222_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7388_ (.A1(_3213_),
    .A2(_3223_),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7389_ (.A1(_3208_),
    .A2(net104),
    .B1(_3060_),
    .B2(_3224_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7390_ (.A1(_3179_),
    .A2(_3212_),
    .B(_3225_),
    .ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7391_ (.I(_3044_),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7392_ (.I(net73),
    .Z(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7393_ (.A1(_1705_),
    .A2(_1633_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7394_ (.A1(_3227_),
    .A2(_3228_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7395_ (.A1(net72),
    .A2(_1585_),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7396_ (.A1(_3213_),
    .A2(_3223_),
    .B(_3230_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7397_ (.A1(_3229_),
    .A2(_3231_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7398_ (.A1(net72),
    .A2(net73),
    .A3(_3211_),
    .Z(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7399_ (.A1(net72),
    .A2(_3211_),
    .B(_3227_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7400_ (.A1(_3233_),
    .A2(_3234_),
    .Z(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7401_ (.A1(_3209_),
    .A2(net105),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7402_ (.A1(_3226_),
    .A2(_3232_),
    .B1(_3235_),
    .B2(_3179_),
    .C(_3236_),
    .ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7403_ (.A1(_0936_),
    .A2(_3233_),
    .Z(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7404_ (.A1(net74),
    .A2(_1603_),
    .Z(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7405_ (.A1(_3213_),
    .A2(_3229_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7406_ (.A1(_3220_),
    .A2(_3222_),
    .B(_3239_),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7407_ (.A1(_3227_),
    .A2(_3228_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7408_ (.A1(_3227_),
    .A2(_3228_),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7409_ (.A1(_3230_),
    .A2(_3241_),
    .B(_3242_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7410_ (.I(_3243_),
    .ZN(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7411_ (.A1(_3240_),
    .A2(_3244_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7412_ (.A1(_3238_),
    .A2(_3245_),
    .ZN(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7413_ (.A1(_3209_),
    .A2(net106),
    .ZN(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7414_ (.A1(_3200_),
    .A2(_3237_),
    .B1(_3246_),
    .B2(_3046_),
    .C(_3247_),
    .ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7415_ (.I(_3208_),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7416_ (.A1(_3248_),
    .A2(net107),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7417_ (.I(_3041_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7418_ (.A1(net74),
    .A2(_3233_),
    .ZN(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7419_ (.A1(_0952_),
    .A2(_3251_),
    .Z(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7420_ (.I(_1637_),
    .Z(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7421_ (.A1(_0952_),
    .A2(_3253_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7422_ (.A1(_0914_),
    .A2(_1704_),
    .B(_1705_),
    .ZN(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7423_ (.A1(net74),
    .A2(_3255_),
    .ZN(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7424_ (.A1(_3238_),
    .A2(_3245_),
    .B(_3256_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7425_ (.A1(_3254_),
    .A2(_3257_),
    .ZN(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7426_ (.A1(_3250_),
    .A2(_3252_),
    .B1(_3258_),
    .B2(_3053_),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7427_ (.A1(_3249_),
    .A2(_3259_),
    .ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7428_ (.I(net77),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7429_ (.A1(_0952_),
    .A2(_3251_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7430_ (.A1(_3260_),
    .A2(_3261_),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7431_ (.I(_1557_),
    .Z(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7432_ (.A1(net77),
    .A2(_3263_),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7433_ (.A1(_3240_),
    .A2(_3244_),
    .B(_3254_),
    .C(_3238_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7434_ (.A1(net75),
    .A2(_3253_),
    .ZN(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7435_ (.A1(net75),
    .A2(_3253_),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7436_ (.A1(_3256_),
    .A2(_3266_),
    .B(_3267_),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _7437_ (.A1(_3264_),
    .A2(_3265_),
    .A3(_3268_),
    .ZN(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7438_ (.A1(_3265_),
    .A2(_3268_),
    .B(_3264_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7439_ (.A1(_3060_),
    .A2(_3270_),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7440_ (.I(_3208_),
    .Z(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7441_ (.A1(_3272_),
    .A2(net109),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7442_ (.A1(_3200_),
    .A2(_3262_),
    .B1(_3269_),
    .B2(_3271_),
    .C(_3273_),
    .ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7443_ (.A1(net77),
    .A2(net78),
    .A3(_3261_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7444_ (.I(net78),
    .Z(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7445_ (.A1(_3260_),
    .A2(_3261_),
    .B(_3275_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7446_ (.A1(_3274_),
    .A2(_3276_),
    .Z(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7447_ (.I(_1525_),
    .Z(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7448_ (.A1(_3260_),
    .A2(_3263_),
    .ZN(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7449_ (.A1(_3279_),
    .A2(_3270_),
    .ZN(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7450_ (.A1(_3275_),
    .A2(_3278_),
    .A3(_3280_),
    .Z(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7451_ (.A1(_3053_),
    .A2(_3281_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7452_ (.A1(_3248_),
    .A2(net110),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7453_ (.A1(_3144_),
    .A2(_3277_),
    .B(_3282_),
    .C(_3283_),
    .ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7454_ (.I(net79),
    .Z(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7455_ (.A1(_3284_),
    .A2(_3274_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7456_ (.A1(net79),
    .A2(_1568_),
    .Z(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7457_ (.A1(net78),
    .A2(_1525_),
    .B1(_3263_),
    .B2(_3260_),
    .ZN(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7458_ (.A1(_3275_),
    .A2(_3278_),
    .ZN(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7459_ (.A1(_3270_),
    .A2(_3287_),
    .B(_3288_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7460_ (.A1(_3286_),
    .A2(_3289_),
    .Z(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7461_ (.A1(_3272_),
    .A2(net111),
    .ZN(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7462_ (.A1(_3076_),
    .A2(_3285_),
    .B1(_3290_),
    .B2(_3046_),
    .C(_3291_),
    .ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7463_ (.I(net80),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7464_ (.A1(_3284_),
    .A2(_3274_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7465_ (.A1(_3292_),
    .A2(_3293_),
    .Z(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7466_ (.I(_1553_),
    .Z(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7467_ (.A1(_3292_),
    .A2(_3295_),
    .ZN(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7468_ (.A1(_3270_),
    .A2(_3287_),
    .ZN(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7469_ (.A1(_3275_),
    .A2(_3278_),
    .B(_3297_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7470_ (.A1(_1437_),
    .A2(_3138_),
    .B(_1414_),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7471_ (.A1(_3284_),
    .A2(_3299_),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7472_ (.A1(_3286_),
    .A2(_3298_),
    .B(_3300_),
    .ZN(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7473_ (.A1(_3296_),
    .A2(_3301_),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7474_ (.A1(_3272_),
    .A2(net112),
    .ZN(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7475_ (.A1(_3076_),
    .A2(_3294_),
    .B1(_3302_),
    .B2(_3226_),
    .C(_3303_),
    .ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7476_ (.A1(net79),
    .A2(net80),
    .A3(_3274_),
    .ZN(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7477_ (.A1(net81),
    .A2(_3304_),
    .Z(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7478_ (.A1(_3248_),
    .A2(net113),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7479_ (.A1(net81),
    .A2(_1444_),
    .ZN(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7480_ (.A1(_1046_),
    .A2(_1881_),
    .ZN(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7481_ (.A1(_3307_),
    .A2(_3308_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7482_ (.A1(_3286_),
    .A2(_3296_),
    .ZN(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7483_ (.A1(_3292_),
    .A2(_3295_),
    .B(_3299_),
    .C(_3284_),
    .ZN(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7484_ (.I(_3311_),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7485_ (.A1(_3292_),
    .A2(_3295_),
    .B1(_3289_),
    .B2(_3310_),
    .C(_3312_),
    .ZN(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7486_ (.A1(_3309_),
    .A2(_3313_),
    .Z(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7487_ (.A1(_3053_),
    .A2(_3314_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7488_ (.A1(_3144_),
    .A2(_3305_),
    .B(_3306_),
    .C(_3315_),
    .ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7489_ (.A1(net82),
    .A2(_1404_),
    .Z(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7490_ (.I(net82),
    .Z(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7491_ (.A1(_3317_),
    .A2(_1404_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7492_ (.A1(_3316_),
    .A2(_3318_),
    .ZN(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7493_ (.A1(_3309_),
    .A2(_3313_),
    .B(_3307_),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7494_ (.A1(_3319_),
    .A2(_3320_),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7495_ (.A1(_1046_),
    .A2(_3304_),
    .ZN(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7496_ (.A1(_3317_),
    .A2(_3322_),
    .ZN(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7497_ (.I(_3041_),
    .Z(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7498_ (.A1(_3272_),
    .A2(net114),
    .ZN(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7499_ (.A1(_3226_),
    .A2(_3321_),
    .B1(_3323_),
    .B2(_3324_),
    .C(_3325_),
    .ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7500_ (.I(net83),
    .Z(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7501_ (.A1(_3317_),
    .A2(_3322_),
    .ZN(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7502_ (.A1(_3326_),
    .A2(_3327_),
    .Z(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7503_ (.I(_3318_),
    .ZN(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7504_ (.A1(_3329_),
    .A2(_3320_),
    .B(_3316_),
    .ZN(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7505_ (.A1(_3326_),
    .A2(_1356_),
    .ZN(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7506_ (.A1(_3330_),
    .A2(_3331_),
    .B(_3044_),
    .ZN(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7507_ (.A1(_3330_),
    .A2(_3331_),
    .B(_3332_),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7508_ (.A1(_3035_),
    .A2(_2855_),
    .B1(_3200_),
    .B2(_3328_),
    .C(_3333_),
    .ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7509_ (.A1(_1088_),
    .A2(_1416_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7510_ (.A1(_1414_),
    .A2(_1415_),
    .ZN(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7511_ (.A1(net84),
    .A2(_3335_),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7512_ (.A1(_3334_),
    .A2(_3336_),
    .ZN(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7513_ (.A1(_3326_),
    .A2(_1356_),
    .ZN(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7514_ (.A1(_3330_),
    .A2(_3331_),
    .B(_3338_),
    .ZN(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7515_ (.A1(_3337_),
    .A2(_3339_),
    .Z(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7516_ (.A1(net82),
    .A2(_3326_),
    .A3(_3322_),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7517_ (.A1(net84),
    .A2(_3341_),
    .Z(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7518_ (.A1(_3051_),
    .A2(net116),
    .ZN(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7519_ (.A1(_3226_),
    .A2(_3340_),
    .B1(_3342_),
    .B2(_3324_),
    .C(_3343_),
    .ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7520_ (.I(net85),
    .Z(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7521_ (.I(_3344_),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7522_ (.I(_1511_),
    .Z(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7523_ (.A1(_3331_),
    .A2(_3337_),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7524_ (.A1(_3309_),
    .A2(_3319_),
    .A3(_3347_),
    .Z(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7525_ (.A1(_3317_),
    .A2(_1404_),
    .ZN(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7526_ (.A1(_3307_),
    .A2(_3318_),
    .B(_3347_),
    .C(_3349_),
    .ZN(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7527_ (.A1(net84),
    .A2(_3335_),
    .ZN(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7528_ (.A1(_3338_),
    .A2(_3351_),
    .B(_3336_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7529_ (.A1(_3350_),
    .A2(_3352_),
    .ZN(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7530_ (.A1(_3313_),
    .A2(_3348_),
    .B(_3353_),
    .ZN(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7531_ (.A1(_3345_),
    .A2(_3346_),
    .A3(_3354_),
    .ZN(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7532_ (.A1(_1088_),
    .A2(_3341_),
    .ZN(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7533_ (.A1(_3345_),
    .A2(_3356_),
    .ZN(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7534_ (.A1(_3051_),
    .A2(net117),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7535_ (.A1(_3045_),
    .A2(_3355_),
    .B1(_3357_),
    .B2(_3324_),
    .C(_3358_),
    .ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7536_ (.I(net86),
    .Z(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7537_ (.I(_1498_),
    .Z(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7538_ (.A1(_3345_),
    .A2(_3346_),
    .Z(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7539_ (.A1(_3345_),
    .A2(_3346_),
    .Z(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7540_ (.A1(_3361_),
    .A2(_3354_),
    .B(_3362_),
    .ZN(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7541_ (.A1(_3359_),
    .A2(_3360_),
    .A3(_3363_),
    .Z(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7542_ (.A1(_3344_),
    .A2(_3356_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7543_ (.A1(_3359_),
    .A2(_3365_),
    .Z(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7544_ (.A1(_3051_),
    .A2(net118),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7545_ (.A1(_3045_),
    .A2(_3364_),
    .B1(_3366_),
    .B2(_3324_),
    .C(_3367_),
    .ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7546_ (.I(net88),
    .Z(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7547_ (.A1(_3344_),
    .A2(net86),
    .A3(_3356_),
    .ZN(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7548_ (.A1(_3368_),
    .A2(_3369_),
    .Z(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7549_ (.A1(_3248_),
    .A2(net120),
    .ZN(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7550_ (.A1(_3368_),
    .A2(_1481_),
    .Z(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7551_ (.A1(_3359_),
    .A2(_3360_),
    .ZN(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7552_ (.A1(_3359_),
    .A2(_3360_),
    .ZN(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7553_ (.A1(_3373_),
    .A2(_3363_),
    .B(_3374_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7554_ (.A1(_3372_),
    .A2(_3375_),
    .B(_3044_),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7555_ (.A1(_3372_),
    .A2(_3375_),
    .B(_3376_),
    .ZN(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7556_ (.A1(_3144_),
    .A2(_3370_),
    .B(_3371_),
    .C(_3377_),
    .ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7557_ (.A1(_3368_),
    .A2(_1481_),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7558_ (.A1(_3372_),
    .A2(_3375_),
    .ZN(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7559_ (.A1(net89),
    .A2(_1381_),
    .Z(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7560_ (.A1(_3378_),
    .A2(_3379_),
    .A3(_3380_),
    .Z(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7561_ (.A1(_3378_),
    .A2(_3379_),
    .B(_3380_),
    .ZN(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7562_ (.A1(_3344_),
    .A2(net86),
    .A3(_3368_),
    .A4(_3356_),
    .ZN(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7563_ (.A1(net89),
    .A2(_3383_),
    .Z(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7564_ (.A1(_3075_),
    .A2(_3384_),
    .ZN(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7565_ (.A1(_3209_),
    .A2(net121),
    .B(_3385_),
    .ZN(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7566_ (.A1(_3045_),
    .A2(_3381_),
    .A3(_3382_),
    .B(_3386_),
    .ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7567_ (.I(net2),
    .Z(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _7568_ (.A1(_1236_),
    .A2(_3387_),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7569_ (.I(net31),
    .Z(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7570_ (.I(net30),
    .Z(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7571_ (.A1(_0587_),
    .A2(_0605_),
    .B(_0707_),
    .ZN(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _7572_ (.A1(_0594_),
    .A2(_3034_),
    .A3(_3391_),
    .ZN(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _7573_ (.A1(_0609_),
    .A2(_0600_),
    .A3(_0611_),
    .A4(_0664_),
    .ZN(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7574_ (.A1(_3392_),
    .A2(_3393_),
    .B(net3),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7575_ (.I(_3394_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7576_ (.A1(_3390_),
    .A2(_3395_),
    .ZN(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _7577_ (.A1(_3389_),
    .A2(_3396_),
    .ZN(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7578_ (.A1(_3388_),
    .A2(_3397_),
    .ZN(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7579_ (.I(_3398_),
    .Z(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7580_ (.I(_3399_),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7581_ (.I(_3034_),
    .Z(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7582_ (.I(_3392_),
    .Z(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7583_ (.I(_3402_),
    .Z(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7584_ (.A1(_2970_),
    .A2(_1981_),
    .ZN(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7585_ (.I(_3404_),
    .Z(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7586_ (.I(_3026_),
    .Z(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7587_ (.I(_3406_),
    .Z(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7588_ (.I0(net40),
    .I1(net49),
    .S(_3407_),
    .Z(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7589_ (.A1(_3405_),
    .A2(_3408_),
    .ZN(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7590_ (.I(_3023_),
    .Z(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7591_ (.I(_3026_),
    .Z(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7592_ (.I(_3411_),
    .Z(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7593_ (.I0(net33),
    .I1(net63),
    .S(_3412_),
    .Z(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7594_ (.I(_0595_),
    .Z(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7595_ (.A1(_3410_),
    .A2(_3413_),
    .B(_3414_),
    .ZN(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7596_ (.I(_3391_),
    .Z(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7597_ (.I(_3416_),
    .Z(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7598_ (.A1(_1901_),
    .A2(_3417_),
    .ZN(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7599_ (.A1(_3409_),
    .A2(_3415_),
    .B(_3418_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7600_ (.A1(net65),
    .A2(_3401_),
    .B1(_0689_),
    .B2(_3403_),
    .C(_3419_),
    .ZN(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7601_ (.I(_3420_),
    .Z(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7602_ (.I(_3398_),
    .Z(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7603_ (.A1(\reg_file.reg_storage[5][0] ),
    .A2(_3422_),
    .ZN(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7604_ (.A1(_3400_),
    .A2(_3421_),
    .B(_3423_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7605_ (.A1(_0975_),
    .A2(_1106_),
    .ZN(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _7606_ (.A1(_0880_),
    .A2(_3390_),
    .A3(_3394_),
    .ZN(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7607_ (.A1(_3424_),
    .A2(_3425_),
    .ZN(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7608_ (.I(_3426_),
    .Z(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7609_ (.I(_3427_),
    .Z(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7610_ (.A1(_0600_),
    .A2(_0661_),
    .B(_0665_),
    .ZN(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7611_ (.I(_3429_),
    .Z(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7612_ (.I(_3430_),
    .Z(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7613_ (.I(_3431_),
    .Z(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7614_ (.I(_3411_),
    .Z(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7615_ (.I(_3023_),
    .Z(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _7616_ (.I0(net44),
    .I1(net64),
    .I2(net41),
    .I3(net50),
    .S0(_3433_),
    .S1(_3434_),
    .Z(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7617_ (.A1(net129),
    .A2(_3435_),
    .ZN(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7618_ (.A1(_0594_),
    .A2(_3034_),
    .ZN(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7619_ (.I(_3437_),
    .Z(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7620_ (.I(_3438_),
    .Z(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7621_ (.A1(net76),
    .A2(_3401_),
    .B1(_1180_),
    .B2(_3439_),
    .C(_3417_),
    .ZN(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7622_ (.A1(_3436_),
    .A2(_3440_),
    .ZN(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7623_ (.A1(_1981_),
    .A2(_3432_),
    .B(_3441_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7624_ (.I(_3442_),
    .Z(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7625_ (.I(_3426_),
    .Z(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7626_ (.A1(\reg_file.reg_storage[5][1] ),
    .A2(_3444_),
    .ZN(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7627_ (.A1(_3428_),
    .A2(_3443_),
    .B(_3445_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7628_ (.I(_3431_),
    .Z(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _7629_ (.I(net51),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7630_ (.A1(net42),
    .A2(_3433_),
    .ZN(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7631_ (.A1(_3447_),
    .A2(_3028_),
    .B(_3448_),
    .ZN(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _7632_ (.A1(_3405_),
    .A2(_3449_),
    .ZN(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7633_ (.I0(net55),
    .I1(net34),
    .S(_3412_),
    .Z(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7634_ (.A1(_3024_),
    .A2(_3451_),
    .B(_3414_),
    .ZN(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7635_ (.A1(_3066_),
    .A2(_3401_),
    .B1(_1238_),
    .B2(_3402_),
    .ZN(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7636_ (.A1(_2085_),
    .A2(_3446_),
    .B1(_3450_),
    .B2(_3452_),
    .C(_3453_),
    .ZN(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7637_ (.I(_3454_),
    .Z(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7638_ (.I(_3455_),
    .Z(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7639_ (.I(_3426_),
    .Z(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7640_ (.I(_3457_),
    .Z(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7641_ (.I0(\reg_file.reg_storage[5][2] ),
    .I1(_3456_),
    .S(_3458_),
    .Z(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7642_ (.I(_3459_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7643_ (.I(_3416_),
    .Z(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7644_ (.I(_3022_),
    .Z(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _7645_ (.I0(net58),
    .I1(net35),
    .I2(net43),
    .I3(net52),
    .S0(_3407_),
    .S1(_3461_),
    .Z(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7646_ (.A1(_3414_),
    .A2(_3462_),
    .ZN(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7647_ (.I(_3437_),
    .Z(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7648_ (.A1(_3047_),
    .A2(_3068_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7649_ (.I(_3416_),
    .Z(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7650_ (.A1(_3069_),
    .A2(_3464_),
    .B(_3465_),
    .C(_3466_),
    .ZN(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _7651_ (.A1(_2148_),
    .A2(_3460_),
    .B1(_3463_),
    .B2(_3467_),
    .ZN(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7652_ (.I(_3468_),
    .Z(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7653_ (.I(_3469_),
    .Z(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7654_ (.I0(\reg_file.reg_storage[5][3] ),
    .I1(_3470_),
    .S(_3458_),
    .Z(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7655_ (.I(_3471_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7656_ (.I(_3430_),
    .Z(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7657_ (.A1(_3081_),
    .A2(_3403_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7658_ (.A1(_3048_),
    .A2(_3080_),
    .B(_3472_),
    .C(_3473_),
    .ZN(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _7659_ (.I0(net59),
    .I1(net36),
    .I2(net45),
    .I3(net53),
    .S0(_3028_),
    .S1(_3410_),
    .Z(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7660_ (.A1(net129),
    .A2(_3475_),
    .Z(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7661_ (.A1(net123),
    .A2(_3432_),
    .B1(_3474_),
    .B2(_3476_),
    .ZN(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7662_ (.I(_3477_),
    .Z(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7663_ (.A1(\reg_file.reg_storage[5][4] ),
    .A2(_3444_),
    .ZN(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7664_ (.A1(_3428_),
    .A2(_3478_),
    .B(_3479_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7665_ (.I(net124),
    .ZN(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7666_ (.I(_3026_),
    .Z(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _7667_ (.I0(net60),
    .I1(net37),
    .I2(net46),
    .I3(net54),
    .S0(_3481_),
    .S1(_3461_),
    .Z(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _7668_ (.A1(_3414_),
    .A2(_3482_),
    .ZN(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7669_ (.I(_0613_),
    .Z(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7670_ (.I(_3484_),
    .Z(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7671_ (.I(_3429_),
    .Z(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7672_ (.A1(_3485_),
    .A2(_3089_),
    .B(_3486_),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7673_ (.A1(_3090_),
    .A2(_3403_),
    .B(_3487_),
    .ZN(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7674_ (.A1(_3480_),
    .A2(_3460_),
    .B1(_3483_),
    .B2(_3488_),
    .ZN(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7675_ (.I(_3489_),
    .Z(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7676_ (.I(_3490_),
    .Z(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7677_ (.I(_3427_),
    .Z(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7678_ (.I0(\reg_file.reg_storage[5][5] ),
    .I1(_3491_),
    .S(_3492_),
    .Z(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7679_ (.I(_3493_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _7680_ (.I0(net61),
    .I1(net38),
    .I2(net47),
    .I3(net56),
    .S0(_3433_),
    .S1(_3434_),
    .Z(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7681_ (.A1(net129),
    .A2(_3494_),
    .Z(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _7682_ (.A1(_3429_),
    .A2(_3437_),
    .ZN(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7683_ (.I(_3496_),
    .Z(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7684_ (.A1(net19),
    .A2(_3138_),
    .ZN(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7685_ (.I(_3486_),
    .Z(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7686_ (.A1(_3048_),
    .A2(_3099_),
    .B1(_3497_),
    .B2(_3498_),
    .C(_3499_),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7687_ (.A1(net125),
    .A2(_3432_),
    .B1(_3495_),
    .B2(_3500_),
    .ZN(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7688_ (.I(_3501_),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7689_ (.A1(\reg_file.reg_storage[5][6] ),
    .A2(_3444_),
    .ZN(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7690_ (.A1(_3428_),
    .A2(_3502_),
    .B(_3503_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _7691_ (.I(_3466_),
    .Z(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7692_ (.I(_3392_),
    .Z(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _7693_ (.I0(net62),
    .I1(net48),
    .I2(net39),
    .I3(net57),
    .S0(_3021_),
    .S1(_3025_),
    .Z(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7694_ (.A1(_3047_),
    .A2(_3115_),
    .B(_3430_),
    .ZN(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7695_ (.A1(_3116_),
    .A2(_3505_),
    .B1(_3506_),
    .B2(_0595_),
    .C(_3507_),
    .ZN(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7696_ (.A1(_2309_),
    .A2(_3504_),
    .B(_3508_),
    .ZN(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7697_ (.I(_3509_),
    .Z(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7698_ (.I(_3510_),
    .Z(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7699_ (.I0(\reg_file.reg_storage[5][7] ),
    .I1(_3511_),
    .S(_3492_),
    .Z(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7700_ (.I(_3512_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7701_ (.A1(_1709_),
    .A2(_0714_),
    .B(_2986_),
    .ZN(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7702_ (.I(_3513_),
    .Z(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7703_ (.I(_3514_),
    .Z(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7704_ (.I0(net63),
    .I1(net40),
    .S(_3027_),
    .Z(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7705_ (.I(_3022_),
    .Z(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7706_ (.I(_0714_),
    .Z(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7707_ (.A1(_3518_),
    .A2(_3032_),
    .B(net49),
    .ZN(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7708_ (.A1(_3517_),
    .A2(_3519_),
    .ZN(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7709_ (.A1(_2976_),
    .A2(_2981_),
    .ZN(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7710_ (.I(_3521_),
    .Z(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7711_ (.A1(_3434_),
    .A2(_3516_),
    .B(_3520_),
    .C(_3522_),
    .ZN(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7712_ (.A1(_3506_),
    .A2(_3513_),
    .Z(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7713_ (.A1(_0594_),
    .A2(_3524_),
    .ZN(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7714_ (.A1(_3515_),
    .A2(_3523_),
    .B(_3525_),
    .ZN(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7715_ (.A1(_3485_),
    .A2(_3123_),
    .B1(_3496_),
    .B2(_3128_),
    .C(_3486_),
    .ZN(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7716_ (.A1(_3526_),
    .A2(_3527_),
    .ZN(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7717_ (.A1(_2350_),
    .A2(_3504_),
    .B(_3528_),
    .ZN(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7718_ (.I(_3529_),
    .Z(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7719_ (.I(_3530_),
    .Z(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7720_ (.I0(\reg_file.reg_storage[5][8] ),
    .I1(_3531_),
    .S(_3492_),
    .Z(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7721_ (.I(_3532_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7722_ (.I0(net64),
    .I1(net41),
    .S(_3412_),
    .Z(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7723_ (.I(_3518_),
    .Z(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7724_ (.A1(_3534_),
    .A2(_3032_),
    .B(net50),
    .ZN(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7725_ (.A1(_3410_),
    .A2(_3535_),
    .ZN(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7726_ (.I(_3521_),
    .Z(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7727_ (.A1(_3024_),
    .A2(_3533_),
    .B(_3536_),
    .C(_3537_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7728_ (.I(_3525_),
    .Z(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7729_ (.A1(_3515_),
    .A2(_3538_),
    .B(_3539_),
    .ZN(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7730_ (.A1(_3048_),
    .A2(_3136_),
    .B1(_3497_),
    .B2(_1829_),
    .C(_3472_),
    .ZN(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _7731_ (.A1(net128),
    .A2(_3432_),
    .B1(_3540_),
    .B2(_3541_),
    .ZN(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7732_ (.I(_3542_),
    .Z(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7733_ (.I(_3457_),
    .Z(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7734_ (.A1(\reg_file.reg_storage[5][9] ),
    .A2(_3544_),
    .ZN(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7735_ (.A1(_3428_),
    .A2(_3543_),
    .B(_3545_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7736_ (.A1(_0595_),
    .A2(_3524_),
    .Z(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7737_ (.I(_3546_),
    .Z(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7738_ (.I0(net34),
    .I1(net42),
    .S(_3027_),
    .Z(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7739_ (.A1(_3447_),
    .A2(_3481_),
    .B(_3517_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7740_ (.A1(_3434_),
    .A2(_3548_),
    .B(_3549_),
    .C(_3522_),
    .ZN(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7741_ (.A1(_3514_),
    .A2(_3550_),
    .ZN(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7742_ (.A1(_1671_),
    .A2(_3402_),
    .B(_3416_),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7743_ (.A1(_3485_),
    .A2(_3146_),
    .B(_3552_),
    .ZN(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7744_ (.A1(_3547_),
    .A2(_3551_),
    .B(_3553_),
    .ZN(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7745_ (.A1(net233),
    .A2(_3504_),
    .B(_3554_),
    .ZN(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7746_ (.I(_3555_),
    .Z(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7747_ (.I(_3556_),
    .Z(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7748_ (.I0(\reg_file.reg_storage[5][10] ),
    .I1(_3557_),
    .S(_3492_),
    .Z(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7749_ (.I(_3558_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7750_ (.I0(net35),
    .I1(net43),
    .S(_3027_),
    .Z(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7751_ (.A1(_3518_),
    .A2(_3031_),
    .B(net52),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7752_ (.A1(_3517_),
    .A2(_3560_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7753_ (.A1(_3461_),
    .A2(_3559_),
    .B(_3561_),
    .C(_3522_),
    .ZN(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7754_ (.A1(_3514_),
    .A2(_3562_),
    .ZN(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7755_ (.A1(_3484_),
    .A2(_3156_),
    .B(_3430_),
    .ZN(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7756_ (.A1(_3161_),
    .A2(_3402_),
    .B1(_3546_),
    .B2(_3563_),
    .C(_3564_),
    .ZN(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7757_ (.A1(_2438_),
    .A2(_3504_),
    .B(_3565_),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7758_ (.I(_3566_),
    .Z(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7759_ (.I(_3567_),
    .Z(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7760_ (.I(_3457_),
    .Z(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7761_ (.I0(\reg_file.reg_storage[5][11] ),
    .I1(_3568_),
    .S(_3569_),
    .Z(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7762_ (.I(_3570_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7763_ (.A1(_2479_),
    .A2(_3460_),
    .ZN(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7764_ (.I(_3484_),
    .Z(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7765_ (.I(_3525_),
    .Z(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7766_ (.I(net53),
    .ZN(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7767_ (.I(net45),
    .ZN(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7768_ (.A1(_3575_),
    .A2(_3406_),
    .ZN(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7769_ (.A1(net36),
    .A2(_3411_),
    .B(_3576_),
    .C(_3404_),
    .ZN(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7770_ (.A1(_3574_),
    .A2(_3405_),
    .A3(_3407_),
    .B(_3577_),
    .ZN(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _7771_ (.I(_3514_),
    .ZN(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7772_ (.A1(_3537_),
    .A2(_3578_),
    .B(_3579_),
    .ZN(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7773_ (.A1(_1692_),
    .A2(_3464_),
    .B(_3466_),
    .ZN(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7774_ (.A1(_3572_),
    .A2(_3167_),
    .B1(_3573_),
    .B2(_3580_),
    .C(_3581_),
    .ZN(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7775_ (.A1(_3571_),
    .A2(_3582_),
    .Z(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7776_ (.I(_3583_),
    .Z(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7777_ (.I(_3584_),
    .Z(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7778_ (.I0(\reg_file.reg_storage[5][12] ),
    .I1(_3585_),
    .S(_3569_),
    .Z(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7779_ (.I(_3586_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7780_ (.A1(_2508_),
    .A2(_3460_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7781_ (.I(net54),
    .ZN(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7782_ (.I(net46),
    .ZN(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7783_ (.A1(_3589_),
    .A2(_3406_),
    .ZN(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7784_ (.A1(net37),
    .A2(_3411_),
    .B(_3590_),
    .C(_3404_),
    .ZN(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7785_ (.A1(_3588_),
    .A2(_3405_),
    .A3(_3407_),
    .B(_3591_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7786_ (.A1(_3537_),
    .A2(_3592_),
    .B(_3579_),
    .ZN(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7787_ (.A1(_3184_),
    .A2(_3438_),
    .B(_3466_),
    .ZN(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7788_ (.A1(_3572_),
    .A2(_3182_),
    .B1(_3573_),
    .B2(_3593_),
    .C(_3594_),
    .ZN(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7789_ (.A1(_3587_),
    .A2(_3595_),
    .Z(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7790_ (.I(_3596_),
    .Z(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7791_ (.I(_3597_),
    .Z(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7792_ (.I0(\reg_file.reg_storage[5][13] ),
    .I1(_3598_),
    .S(_3569_),
    .Z(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7793_ (.I(_3599_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7794_ (.I(_3427_),
    .Z(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7795_ (.I(_3472_),
    .Z(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7796_ (.I0(net38),
    .I1(net47),
    .S(_3412_),
    .Z(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7797_ (.A1(_3518_),
    .A2(_3032_),
    .B(net56),
    .ZN(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7798_ (.A1(_3410_),
    .A2(_3603_),
    .ZN(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7799_ (.A1(_3024_),
    .A2(_3602_),
    .B(_3604_),
    .C(_3537_),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7800_ (.A1(_3515_),
    .A2(_3605_),
    .B(_3539_),
    .ZN(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7801_ (.I(_3572_),
    .Z(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7802_ (.A1(_1710_),
    .A2(_3439_),
    .ZN(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7803_ (.A1(_3607_),
    .A2(_3194_),
    .B(_3446_),
    .C(_3608_),
    .ZN(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _7804_ (.A1(net102),
    .A2(_3601_),
    .B1(_3606_),
    .B2(_3609_),
    .ZN(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7805_ (.I(_3610_),
    .Z(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7806_ (.A1(\reg_file.reg_storage[5][14] ),
    .A2(_3544_),
    .ZN(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7807_ (.A1(_3600_),
    .A2(_3611_),
    .B(_3612_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7808_ (.A1(net103),
    .A2(_3472_),
    .ZN(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7809_ (.I(net57),
    .ZN(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7810_ (.A1(_3614_),
    .A2(_3433_),
    .B(_3461_),
    .ZN(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7811_ (.A1(net39),
    .A2(_3517_),
    .A3(_3481_),
    .Z(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7812_ (.A1(_3522_),
    .A2(_3615_),
    .A3(_3616_),
    .ZN(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7813_ (.A1(_3515_),
    .A2(_3617_),
    .ZN(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7814_ (.A1(_3205_),
    .A2(_3438_),
    .ZN(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7815_ (.A1(_3572_),
    .A2(_3202_),
    .B(_3486_),
    .C(_3619_),
    .ZN(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7816_ (.A1(_3547_),
    .A2(_3618_),
    .B(_3620_),
    .ZN(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7817_ (.A1(_3613_),
    .A2(_3621_),
    .ZN(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7818_ (.I(_3622_),
    .Z(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7819_ (.I(_3623_),
    .Z(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7820_ (.I0(\reg_file.reg_storage[5][15] ),
    .I1(_3624_),
    .S(_3569_),
    .Z(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7821_ (.I(_3625_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7822_ (.A1(_3010_),
    .A2(_3408_),
    .ZN(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7823_ (.A1(_3614_),
    .A2(_3022_),
    .ZN(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7824_ (.A1(net39),
    .A2(_3023_),
    .B(_3627_),
    .ZN(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7825_ (.A1(net48),
    .A2(_3404_),
    .A3(_3406_),
    .ZN(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7826_ (.A1(_3481_),
    .A2(_3628_),
    .B(_3629_),
    .ZN(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7827_ (.A1(_2982_),
    .A2(_3630_),
    .B(_3579_),
    .ZN(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7828_ (.I(_3631_),
    .Z(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7829_ (.A1(_3626_),
    .A2(_3632_),
    .B(_3539_),
    .ZN(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7830_ (.I(_3431_),
    .Z(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7831_ (.A1(_1585_),
    .A2(_3439_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7832_ (.A1(_3607_),
    .A2(_3212_),
    .B(_3634_),
    .C(_3635_),
    .ZN(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7833_ (.A1(net104),
    .A2(_3601_),
    .B1(_3633_),
    .B2(_3636_),
    .ZN(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7834_ (.I(_3637_),
    .Z(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7835_ (.A1(\reg_file.reg_storage[5][16] ),
    .A2(_3544_),
    .ZN(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7836_ (.A1(_3600_),
    .A2(_3638_),
    .B(_3639_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7837_ (.I(_3631_),
    .Z(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7838_ (.I(_3534_),
    .Z(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7839_ (.I(_3036_),
    .Z(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7840_ (.A1(_2968_),
    .A2(_3641_),
    .A3(_3642_),
    .A4(net41),
    .ZN(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7841_ (.A1(_3640_),
    .A2(_3643_),
    .B(_3539_),
    .ZN(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7842_ (.I(_3438_),
    .Z(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7843_ (.A1(_3228_),
    .A2(_3645_),
    .ZN(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7844_ (.A1(_3607_),
    .A2(_3235_),
    .B(_3634_),
    .C(_3646_),
    .ZN(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _7845_ (.A1(net105),
    .A2(_3601_),
    .B1(_3644_),
    .B2(_3647_),
    .ZN(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7846_ (.I(_3648_),
    .Z(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7847_ (.A1(\reg_file.reg_storage[5][17] ),
    .A2(_3544_),
    .ZN(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7848_ (.A1(_3600_),
    .A2(_3649_),
    .B(_3650_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7849_ (.A1(_3010_),
    .A2(_3449_),
    .ZN(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7850_ (.I(_3525_),
    .Z(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7851_ (.A1(_3640_),
    .A2(_3651_),
    .B(_3652_),
    .ZN(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7852_ (.A1(_3255_),
    .A2(_3645_),
    .ZN(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7853_ (.A1(_3607_),
    .A2(_3237_),
    .B(_3634_),
    .C(_3654_),
    .ZN(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7854_ (.A1(net106),
    .A2(_3601_),
    .B1(_3653_),
    .B2(_3655_),
    .ZN(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7855_ (.I(_3656_),
    .Z(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7856_ (.I(_3457_),
    .Z(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7857_ (.A1(\reg_file.reg_storage[5][18] ),
    .A2(_3658_),
    .ZN(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7858_ (.A1(_3600_),
    .A2(_3657_),
    .B(_3659_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7859_ (.I(_3427_),
    .Z(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7860_ (.I(_3431_),
    .Z(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7861_ (.A1(_2968_),
    .A2(_3641_),
    .A3(_3642_),
    .A4(net43),
    .ZN(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7862_ (.A1(_3640_),
    .A2(_3662_),
    .B(_3652_),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7863_ (.A1(_3401_),
    .A2(_3252_),
    .B1(_3439_),
    .B2(_3253_),
    .ZN(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7864_ (.A1(_3446_),
    .A2(_3664_),
    .ZN(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7865_ (.A1(net107),
    .A2(_3661_),
    .B1(_3663_),
    .B2(_3665_),
    .ZN(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7866_ (.I(_3666_),
    .Z(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7867_ (.A1(\reg_file.reg_storage[5][19] ),
    .A2(_3658_),
    .ZN(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7868_ (.A1(_3660_),
    .A2(_3667_),
    .B(_3668_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7869_ (.A1(_2968_),
    .A2(_3641_),
    .A3(_3642_),
    .A4(net45),
    .ZN(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7870_ (.A1(_3640_),
    .A2(_3669_),
    .B(_3652_),
    .ZN(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7871_ (.I(_3485_),
    .Z(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7872_ (.A1(_3263_),
    .A2(_3645_),
    .ZN(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7873_ (.A1(_3671_),
    .A2(_3262_),
    .B(_3634_),
    .C(_3672_),
    .ZN(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7874_ (.A1(net109),
    .A2(_3661_),
    .B1(_3670_),
    .B2(_3673_),
    .ZN(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7875_ (.I(_3674_),
    .Z(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7876_ (.A1(\reg_file.reg_storage[5][20] ),
    .A2(_3658_),
    .ZN(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7877_ (.A1(_3660_),
    .A2(_3675_),
    .B(_3676_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7878_ (.A1(_2967_),
    .A2(_3641_),
    .A3(_3642_),
    .A4(net46),
    .ZN(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7879_ (.A1(_3632_),
    .A2(_3677_),
    .B(_3652_),
    .ZN(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7880_ (.A1(_3278_),
    .A2(_3645_),
    .ZN(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7881_ (.A1(_3671_),
    .A2(_3277_),
    .B(_3499_),
    .C(_3679_),
    .ZN(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7882_ (.A1(net110),
    .A2(_3661_),
    .B1(_3678_),
    .B2(_3680_),
    .ZN(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7883_ (.I(_3681_),
    .Z(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7884_ (.A1(\reg_file.reg_storage[5][21] ),
    .A2(_3658_),
    .ZN(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7885_ (.A1(_3660_),
    .A2(_3682_),
    .B(_3683_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7886_ (.A1(_2967_),
    .A2(_3534_),
    .A3(_3036_),
    .A4(net47),
    .ZN(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7887_ (.A1(_3632_),
    .A2(_3684_),
    .B(_3573_),
    .ZN(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7888_ (.A1(_3299_),
    .A2(_3464_),
    .ZN(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7889_ (.A1(_3671_),
    .A2(_3285_),
    .B(_3499_),
    .C(_3686_),
    .ZN(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7890_ (.A1(net111),
    .A2(_3661_),
    .B1(_3685_),
    .B2(_3687_),
    .ZN(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7891_ (.I(_3688_),
    .Z(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7892_ (.A1(\reg_file.reg_storage[5][22] ),
    .A2(_3458_),
    .ZN(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7893_ (.A1(_3660_),
    .A2(_3689_),
    .B(_3690_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _7894_ (.A1(_2967_),
    .A2(_3534_),
    .A3(_3036_),
    .A4(net48),
    .ZN(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _7895_ (.A1(_3632_),
    .A2(_3691_),
    .B(_3573_),
    .ZN(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7896_ (.A1(_3295_),
    .A2(_3464_),
    .ZN(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7897_ (.A1(_3671_),
    .A2(_3294_),
    .B(_3499_),
    .C(_3693_),
    .ZN(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7898_ (.A1(net112),
    .A2(_3446_),
    .B1(_3692_),
    .B2(_3694_),
    .ZN(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7899_ (.I(_3695_),
    .Z(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7900_ (.A1(\reg_file.reg_storage[5][23] ),
    .A2(_3458_),
    .ZN(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7901_ (.A1(_3444_),
    .A2(_3696_),
    .B(_3697_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7902_ (.I(_3417_),
    .Z(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7903_ (.I(_3547_),
    .Z(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7904_ (.I(_3631_),
    .Z(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7905_ (.A1(_2978_),
    .A2(_3519_),
    .B(_3700_),
    .ZN(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7906_ (.I(_3484_),
    .Z(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _7907_ (.A1(_3702_),
    .A2(_3305_),
    .B1(_3497_),
    .B2(_1881_),
    .ZN(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7908_ (.A1(net113),
    .A2(_3698_),
    .B1(_3699_),
    .B2(_3701_),
    .C(_3703_),
    .ZN(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7909_ (.I(_3704_),
    .Z(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7910_ (.A1(\reg_file.reg_storage[5][24] ),
    .A2(_3422_),
    .ZN(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7911_ (.A1(_3400_),
    .A2(_3705_),
    .B(_3706_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7912_ (.A1(_2978_),
    .A2(_3535_),
    .B(_3700_),
    .ZN(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _7913_ (.A1(_3702_),
    .A2(_3323_),
    .B1(_3497_),
    .B2(_1384_),
    .ZN(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7914_ (.A1(net114),
    .A2(_3698_),
    .B1(_3699_),
    .B2(_3707_),
    .C(_3708_),
    .ZN(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7915_ (.I(_3709_),
    .Z(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7916_ (.A1(\reg_file.reg_storage[5][25] ),
    .A2(_3422_),
    .ZN(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7917_ (.A1(_3400_),
    .A2(_3710_),
    .B(_3711_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7918_ (.I(_2977_),
    .Z(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7919_ (.I(_3631_),
    .Z(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _7920_ (.A1(_3447_),
    .A2(_3712_),
    .A3(_3029_),
    .B(_3713_),
    .ZN(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7921_ (.I(_3047_),
    .Z(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7922_ (.A1(_1356_),
    .A2(_3403_),
    .ZN(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7923_ (.A1(_3715_),
    .A2(_3328_),
    .B(_3716_),
    .ZN(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7924_ (.A1(net115),
    .A2(_3698_),
    .B1(_3699_),
    .B2(_3714_),
    .C(_3717_),
    .ZN(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7925_ (.I(_3718_),
    .Z(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7926_ (.I(_3398_),
    .Z(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7927_ (.A1(\reg_file.reg_storage[5][26] ),
    .A2(_3720_),
    .ZN(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7928_ (.A1(_3400_),
    .A2(_3719_),
    .B(_3721_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7929_ (.I(_3399_),
    .Z(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7930_ (.A1(_3712_),
    .A2(_3560_),
    .B(_3700_),
    .ZN(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _7931_ (.A1(_3702_),
    .A2(_3342_),
    .B1(_3496_),
    .B2(_1416_),
    .ZN(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7932_ (.A1(net116),
    .A2(_3698_),
    .B1(_3699_),
    .B2(_3723_),
    .C(_3724_),
    .ZN(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7933_ (.I(_3725_),
    .Z(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7934_ (.A1(\reg_file.reg_storage[5][27] ),
    .A2(_3720_),
    .ZN(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7935_ (.A1(_3722_),
    .A2(_3726_),
    .B(_3727_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7936_ (.I(_3417_),
    .Z(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7937_ (.I(_3547_),
    .Z(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7938_ (.A1(_3574_),
    .A2(_3712_),
    .A3(_3029_),
    .B(_3713_),
    .ZN(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7939_ (.A1(_3346_),
    .A2(_3505_),
    .ZN(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7940_ (.A1(_3715_),
    .A2(_3357_),
    .B(_3731_),
    .ZN(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7941_ (.A1(net117),
    .A2(_3728_),
    .B1(_3729_),
    .B2(_3730_),
    .C(_3732_),
    .ZN(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7942_ (.I(_3733_),
    .Z(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7943_ (.A1(\reg_file.reg_storage[5][28] ),
    .A2(_3720_),
    .ZN(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7944_ (.A1(_3722_),
    .A2(_3734_),
    .B(_3735_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7945_ (.A1(_3588_),
    .A2(_2977_),
    .A3(_3029_),
    .B(_3713_),
    .ZN(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7946_ (.A1(_3360_),
    .A2(_3505_),
    .ZN(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7947_ (.A1(_3715_),
    .A2(_3366_),
    .B(_3737_),
    .ZN(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7948_ (.A1(net118),
    .A2(_3728_),
    .B1(_3729_),
    .B2(_3736_),
    .C(_3738_),
    .ZN(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7949_ (.I(_3739_),
    .Z(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7950_ (.A1(\reg_file.reg_storage[5][29] ),
    .A2(_3720_),
    .ZN(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7951_ (.A1(_3722_),
    .A2(_3740_),
    .B(_3741_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7952_ (.A1(_3712_),
    .A2(_3603_),
    .B(_3700_),
    .ZN(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7953_ (.A1(_1481_),
    .A2(_3505_),
    .ZN(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7954_ (.A1(_3715_),
    .A2(_3370_),
    .B(_3743_),
    .ZN(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7955_ (.A1(net120),
    .A2(_3728_),
    .B1(_3729_),
    .B2(_3742_),
    .C(_3744_),
    .ZN(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7956_ (.I(_3745_),
    .Z(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7957_ (.A1(\reg_file.reg_storage[5][30] ),
    .A2(_3399_),
    .ZN(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7958_ (.A1(_3722_),
    .A2(_3746_),
    .B(_3747_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7959_ (.A1(_3614_),
    .A2(_2977_),
    .A3(_3028_),
    .B(_3713_),
    .ZN(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _7960_ (.A1(_3702_),
    .A2(_3384_),
    .B1(_3496_),
    .B2(_1381_),
    .ZN(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7961_ (.A1(net211),
    .A2(_3728_),
    .B1(_3729_),
    .B2(_3748_),
    .C(_3749_),
    .ZN(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7962_ (.I(_3750_),
    .Z(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7963_ (.A1(\reg_file.reg_storage[5][31] ),
    .A2(_3399_),
    .ZN(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7964_ (.A1(_3422_),
    .A2(_3751_),
    .B(_3752_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _7965_ (.A1(_0975_),
    .A2(net2),
    .ZN(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _7966_ (.A1(_0880_),
    .A2(_3396_),
    .ZN(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7967_ (.A1(_3753_),
    .A2(_3754_),
    .ZN(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7968_ (.I(_3755_),
    .Z(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7969_ (.I(_3756_),
    .Z(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7970_ (.I(_3755_),
    .Z(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7971_ (.A1(\reg_file.reg_storage[3][0] ),
    .A2(_3758_),
    .ZN(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7972_ (.A1(_3421_),
    .A2(_3757_),
    .B(_3759_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7973_ (.I(_0975_),
    .Z(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _7974_ (.A1(_3389_),
    .A2(_3390_),
    .A3(_3394_),
    .ZN(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7975_ (.A1(_3760_),
    .A2(_3387_),
    .A3(_3761_),
    .ZN(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7976_ (.I(_3762_),
    .Z(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7977_ (.I(_3763_),
    .Z(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7978_ (.I(_3764_),
    .Z(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7979_ (.I(_3762_),
    .Z(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7980_ (.A1(\reg_file.reg_storage[3][1] ),
    .A2(_3766_),
    .ZN(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7981_ (.A1(_3443_),
    .A2(_3765_),
    .B(_3767_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7982_ (.I(_3762_),
    .Z(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7983_ (.I(_3768_),
    .Z(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7984_ (.I0(\reg_file.reg_storage[3][2] ),
    .I1(_3456_),
    .S(_3769_),
    .Z(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7985_ (.I(_3770_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7986_ (.I0(\reg_file.reg_storage[3][3] ),
    .I1(_3470_),
    .S(_3769_),
    .Z(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7987_ (.I(_3771_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7988_ (.A1(\reg_file.reg_storage[3][4] ),
    .A2(_3766_),
    .ZN(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7989_ (.A1(_3478_),
    .A2(_3765_),
    .B(_3772_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7990_ (.I0(\reg_file.reg_storage[3][5] ),
    .I1(_3491_),
    .S(_3769_),
    .Z(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7991_ (.I(_3773_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7992_ (.A1(\reg_file.reg_storage[3][6] ),
    .A2(_3766_),
    .ZN(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7993_ (.A1(_3502_),
    .A2(_3765_),
    .B(_3774_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7994_ (.I(_3763_),
    .Z(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7995_ (.I0(\reg_file.reg_storage[3][7] ),
    .I1(_3511_),
    .S(_3775_),
    .Z(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7996_ (.I(_3776_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7997_ (.I0(\reg_file.reg_storage[3][8] ),
    .I1(_3531_),
    .S(_3775_),
    .Z(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7998_ (.I(_3777_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7999_ (.I(_3763_),
    .Z(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8000_ (.A1(\reg_file.reg_storage[3][9] ),
    .A2(_3778_),
    .ZN(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8001_ (.A1(_3543_),
    .A2(_3765_),
    .B(_3779_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8002_ (.I0(\reg_file.reg_storage[3][10] ),
    .I1(_3557_),
    .S(_3775_),
    .Z(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8003_ (.I(_3780_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8004_ (.I0(\reg_file.reg_storage[3][11] ),
    .I1(_3568_),
    .S(_3775_),
    .Z(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8005_ (.I(_3781_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8006_ (.I0(\reg_file.reg_storage[3][12] ),
    .I1(_3585_),
    .S(_3768_),
    .Z(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8007_ (.I(_3782_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8008_ (.I0(\reg_file.reg_storage[3][13] ),
    .I1(_3598_),
    .S(_3768_),
    .Z(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8009_ (.I(_3783_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8010_ (.I(_3764_),
    .Z(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8011_ (.A1(\reg_file.reg_storage[3][14] ),
    .A2(_3778_),
    .ZN(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8012_ (.A1(_3611_),
    .A2(_3784_),
    .B(_3785_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8013_ (.I0(\reg_file.reg_storage[3][15] ),
    .I1(_3624_),
    .S(_3768_),
    .Z(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8014_ (.I(_3786_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8015_ (.A1(\reg_file.reg_storage[3][16] ),
    .A2(_3778_),
    .ZN(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8016_ (.A1(_3638_),
    .A2(_3784_),
    .B(_3787_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8017_ (.A1(\reg_file.reg_storage[3][17] ),
    .A2(_3778_),
    .ZN(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8018_ (.A1(_3649_),
    .A2(_3784_),
    .B(_3788_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8019_ (.I(_3763_),
    .Z(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8020_ (.A1(\reg_file.reg_storage[3][18] ),
    .A2(_3789_),
    .ZN(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8021_ (.A1(_3657_),
    .A2(_3784_),
    .B(_3790_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8022_ (.I(_3769_),
    .Z(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8023_ (.A1(\reg_file.reg_storage[3][19] ),
    .A2(_3789_),
    .ZN(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8024_ (.A1(_3667_),
    .A2(_3791_),
    .B(_3792_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8025_ (.A1(\reg_file.reg_storage[3][20] ),
    .A2(_3789_),
    .ZN(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8026_ (.A1(_3675_),
    .A2(_3791_),
    .B(_3793_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8027_ (.A1(\reg_file.reg_storage[3][21] ),
    .A2(_3789_),
    .ZN(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8028_ (.A1(_3682_),
    .A2(_3791_),
    .B(_3794_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8029_ (.A1(\reg_file.reg_storage[3][22] ),
    .A2(_3764_),
    .ZN(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8030_ (.A1(_3689_),
    .A2(_3791_),
    .B(_3795_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8031_ (.A1(\reg_file.reg_storage[3][23] ),
    .A2(_3764_),
    .ZN(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8032_ (.A1(_3696_),
    .A2(_3766_),
    .B(_3796_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8033_ (.A1(\reg_file.reg_storage[3][24] ),
    .A2(_3758_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8034_ (.A1(_3705_),
    .A2(_3757_),
    .B(_3797_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8035_ (.A1(\reg_file.reg_storage[3][25] ),
    .A2(_3758_),
    .ZN(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8036_ (.A1(_3710_),
    .A2(_3757_),
    .B(_3798_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8037_ (.I(_3755_),
    .Z(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8038_ (.A1(\reg_file.reg_storage[3][26] ),
    .A2(_3799_),
    .ZN(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8039_ (.A1(_3719_),
    .A2(_3757_),
    .B(_3800_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8040_ (.I(_3756_),
    .Z(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8041_ (.A1(\reg_file.reg_storage[3][27] ),
    .A2(_3799_),
    .ZN(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8042_ (.A1(_3726_),
    .A2(_3801_),
    .B(_3802_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8043_ (.A1(\reg_file.reg_storage[3][28] ),
    .A2(_3799_),
    .ZN(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8044_ (.A1(_3734_),
    .A2(_3801_),
    .B(_3803_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8045_ (.A1(\reg_file.reg_storage[3][29] ),
    .A2(_3799_),
    .ZN(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8046_ (.A1(_3740_),
    .A2(_3801_),
    .B(_3804_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8047_ (.A1(\reg_file.reg_storage[3][30] ),
    .A2(_3756_),
    .ZN(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8048_ (.A1(_3746_),
    .A2(_3801_),
    .B(_3805_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8049_ (.A1(\reg_file.reg_storage[3][31] ),
    .A2(_3756_),
    .ZN(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8050_ (.A1(_3751_),
    .A2(_3758_),
    .B(_3806_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8051_ (.I(net30),
    .ZN(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8052_ (.A1(_3389_),
    .A2(_3807_),
    .A3(_3394_),
    .Z(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8053_ (.I(_3808_),
    .Z(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8054_ (.A1(_3753_),
    .A2(_3809_),
    .ZN(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8055_ (.I(_3810_),
    .Z(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8056_ (.I(_3811_),
    .Z(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8057_ (.I(_3810_),
    .Z(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8058_ (.A1(\reg_file.reg_storage[2][0] ),
    .A2(_3813_),
    .ZN(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8059_ (.A1(_3421_),
    .A2(_3812_),
    .B(_3814_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8060_ (.A1(_3753_),
    .A2(_3808_),
    .Z(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8061_ (.I(_3815_),
    .Z(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8062_ (.I(_3816_),
    .Z(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8063_ (.I(_3817_),
    .Z(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8064_ (.I(_3815_),
    .Z(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8065_ (.A1(\reg_file.reg_storage[2][1] ),
    .A2(_3819_),
    .ZN(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8066_ (.A1(_3443_),
    .A2(_3818_),
    .B(_3820_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8067_ (.I(_3815_),
    .Z(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8068_ (.I(_3821_),
    .Z(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8069_ (.I0(\reg_file.reg_storage[2][2] ),
    .I1(_3456_),
    .S(_3822_),
    .Z(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8070_ (.I(_3823_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8071_ (.I0(\reg_file.reg_storage[2][3] ),
    .I1(_3470_),
    .S(_3822_),
    .Z(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8072_ (.I(_3824_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8073_ (.A1(\reg_file.reg_storage[2][4] ),
    .A2(_3819_),
    .ZN(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8074_ (.A1(_3478_),
    .A2(_3818_),
    .B(_3825_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8075_ (.I0(\reg_file.reg_storage[2][5] ),
    .I1(_3491_),
    .S(_3822_),
    .Z(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8076_ (.I(_3826_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8077_ (.A1(\reg_file.reg_storage[2][6] ),
    .A2(_3819_),
    .ZN(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8078_ (.A1(_3502_),
    .A2(_3818_),
    .B(_3827_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8079_ (.I(_3816_),
    .Z(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8080_ (.I0(\reg_file.reg_storage[2][7] ),
    .I1(_3511_),
    .S(_3828_),
    .Z(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8081_ (.I(_3829_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8082_ (.I0(\reg_file.reg_storage[2][8] ),
    .I1(_3531_),
    .S(_3828_),
    .Z(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8083_ (.I(_3830_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8084_ (.I(_3816_),
    .Z(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8085_ (.A1(\reg_file.reg_storage[2][9] ),
    .A2(_3831_),
    .ZN(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8086_ (.A1(_3543_),
    .A2(_3818_),
    .B(_3832_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8087_ (.I0(\reg_file.reg_storage[2][10] ),
    .I1(_3557_),
    .S(_3828_),
    .Z(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8088_ (.I(_3833_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8089_ (.I0(\reg_file.reg_storage[2][11] ),
    .I1(_3568_),
    .S(_3828_),
    .Z(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8090_ (.I(_3834_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8091_ (.I0(\reg_file.reg_storage[2][12] ),
    .I1(_3585_),
    .S(_3821_),
    .Z(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8092_ (.I(_3835_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8093_ (.I0(\reg_file.reg_storage[2][13] ),
    .I1(_3598_),
    .S(_3821_),
    .Z(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8094_ (.I(_3836_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8095_ (.I(_3817_),
    .Z(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8096_ (.A1(\reg_file.reg_storage[2][14] ),
    .A2(_3831_),
    .ZN(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8097_ (.A1(_3611_),
    .A2(_3837_),
    .B(_3838_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8098_ (.I0(\reg_file.reg_storage[2][15] ),
    .I1(_3624_),
    .S(_3821_),
    .Z(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8099_ (.I(_3839_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8100_ (.A1(\reg_file.reg_storage[2][16] ),
    .A2(_3831_),
    .ZN(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8101_ (.A1(_3638_),
    .A2(_3837_),
    .B(_3840_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8102_ (.A1(\reg_file.reg_storage[2][17] ),
    .A2(_3831_),
    .ZN(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8103_ (.A1(_3649_),
    .A2(_3837_),
    .B(_3841_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8104_ (.I(_3816_),
    .Z(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8105_ (.A1(\reg_file.reg_storage[2][18] ),
    .A2(_3842_),
    .ZN(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8106_ (.A1(_3657_),
    .A2(_3837_),
    .B(_3843_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8107_ (.I(_3822_),
    .Z(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8108_ (.A1(\reg_file.reg_storage[2][19] ),
    .A2(_3842_),
    .ZN(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8109_ (.A1(_3667_),
    .A2(_3844_),
    .B(_3845_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8110_ (.A1(\reg_file.reg_storage[2][20] ),
    .A2(_3842_),
    .ZN(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8111_ (.A1(_3675_),
    .A2(_3844_),
    .B(_3846_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8112_ (.A1(\reg_file.reg_storage[2][21] ),
    .A2(_3842_),
    .ZN(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8113_ (.A1(_3682_),
    .A2(_3844_),
    .B(_3847_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8114_ (.A1(\reg_file.reg_storage[2][22] ),
    .A2(_3817_),
    .ZN(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8115_ (.A1(_3689_),
    .A2(_3844_),
    .B(_3848_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8116_ (.A1(\reg_file.reg_storage[2][23] ),
    .A2(_3817_),
    .ZN(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8117_ (.A1(_3696_),
    .A2(_3819_),
    .B(_3849_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8118_ (.A1(\reg_file.reg_storage[2][24] ),
    .A2(_3813_),
    .ZN(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8119_ (.A1(_3705_),
    .A2(_3812_),
    .B(_3850_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8120_ (.A1(\reg_file.reg_storage[2][25] ),
    .A2(_3813_),
    .ZN(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8121_ (.A1(_3710_),
    .A2(_3812_),
    .B(_3851_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8122_ (.I(_3810_),
    .Z(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8123_ (.A1(\reg_file.reg_storage[2][26] ),
    .A2(_3852_),
    .ZN(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8124_ (.A1(_3719_),
    .A2(_3812_),
    .B(_3853_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8125_ (.I(_3811_),
    .Z(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8126_ (.A1(\reg_file.reg_storage[2][27] ),
    .A2(_3852_),
    .ZN(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8127_ (.A1(_3726_),
    .A2(_3854_),
    .B(_3855_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8128_ (.A1(\reg_file.reg_storage[2][28] ),
    .A2(_3852_),
    .ZN(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8129_ (.A1(_3734_),
    .A2(_3854_),
    .B(_3856_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8130_ (.A1(\reg_file.reg_storage[2][29] ),
    .A2(_3852_),
    .ZN(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8131_ (.A1(_3740_),
    .A2(_3854_),
    .B(_3857_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8132_ (.A1(\reg_file.reg_storage[2][30] ),
    .A2(_3811_),
    .ZN(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8133_ (.A1(_3746_),
    .A2(_3854_),
    .B(_3858_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8134_ (.A1(\reg_file.reg_storage[2][31] ),
    .A2(_3811_),
    .ZN(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8135_ (.A1(_3751_),
    .A2(_3813_),
    .B(_3859_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8136_ (.A1(_3388_),
    .A2(_3809_),
    .ZN(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8137_ (.I(_3860_),
    .Z(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8138_ (.I(_3861_),
    .Z(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8139_ (.I(_3860_),
    .Z(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8140_ (.A1(\reg_file.reg_storage[6][0] ),
    .A2(_3863_),
    .ZN(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8141_ (.A1(_3421_),
    .A2(_3862_),
    .B(_3864_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8142_ (.A1(_3389_),
    .A2(_3807_),
    .A3(_3395_),
    .ZN(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8143_ (.A1(_3424_),
    .A2(_3865_),
    .ZN(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8144_ (.I(_3866_),
    .Z(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8145_ (.I(_3867_),
    .Z(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8146_ (.I(_3868_),
    .Z(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8147_ (.I(_3866_),
    .Z(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8148_ (.A1(\reg_file.reg_storage[6][1] ),
    .A2(_3870_),
    .ZN(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8149_ (.A1(_3443_),
    .A2(_3869_),
    .B(_3871_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8150_ (.I(_3866_),
    .Z(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8151_ (.I(_3872_),
    .Z(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8152_ (.I0(\reg_file.reg_storage[6][2] ),
    .I1(_3456_),
    .S(_3873_),
    .Z(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8153_ (.I(_3874_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8154_ (.I0(\reg_file.reg_storage[6][3] ),
    .I1(_3470_),
    .S(_3873_),
    .Z(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8155_ (.I(_3875_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8156_ (.A1(\reg_file.reg_storage[6][4] ),
    .A2(_3870_),
    .ZN(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8157_ (.A1(_3478_),
    .A2(_3869_),
    .B(_3876_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8158_ (.I0(\reg_file.reg_storage[6][5] ),
    .I1(_3491_),
    .S(_3873_),
    .Z(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8159_ (.I(_3877_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8160_ (.A1(\reg_file.reg_storage[6][6] ),
    .A2(_3870_),
    .ZN(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8161_ (.A1(_3502_),
    .A2(_3869_),
    .B(_3878_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8162_ (.I(_3867_),
    .Z(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8163_ (.I0(\reg_file.reg_storage[6][7] ),
    .I1(_3511_),
    .S(_3879_),
    .Z(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8164_ (.I(_3880_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8165_ (.I0(\reg_file.reg_storage[6][8] ),
    .I1(_3531_),
    .S(_3879_),
    .Z(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8166_ (.I(_3881_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8167_ (.I(_3867_),
    .Z(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8168_ (.A1(\reg_file.reg_storage[6][9] ),
    .A2(_3882_),
    .ZN(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8169_ (.A1(_3543_),
    .A2(_3869_),
    .B(_3883_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8170_ (.I0(\reg_file.reg_storage[6][10] ),
    .I1(_3557_),
    .S(_3879_),
    .Z(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8171_ (.I(_3884_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8172_ (.I0(\reg_file.reg_storage[6][11] ),
    .I1(_3568_),
    .S(_3879_),
    .Z(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8173_ (.I(_3885_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8174_ (.I0(\reg_file.reg_storage[6][12] ),
    .I1(_3585_),
    .S(_3872_),
    .Z(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8175_ (.I(_3886_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8176_ (.I0(\reg_file.reg_storage[6][13] ),
    .I1(_3598_),
    .S(_3872_),
    .Z(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8177_ (.I(_3887_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8178_ (.I(_3868_),
    .Z(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8179_ (.A1(\reg_file.reg_storage[6][14] ),
    .A2(_3882_),
    .ZN(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8180_ (.A1(_3611_),
    .A2(_3888_),
    .B(_3889_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8181_ (.I0(\reg_file.reg_storage[6][15] ),
    .I1(_3624_),
    .S(_3872_),
    .Z(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8182_ (.I(_3890_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8183_ (.A1(\reg_file.reg_storage[6][16] ),
    .A2(_3882_),
    .ZN(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8184_ (.A1(_3638_),
    .A2(_3888_),
    .B(_3891_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8185_ (.A1(\reg_file.reg_storage[6][17] ),
    .A2(_3882_),
    .ZN(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8186_ (.A1(_3649_),
    .A2(_3888_),
    .B(_3892_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8187_ (.I(_3867_),
    .Z(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8188_ (.A1(\reg_file.reg_storage[6][18] ),
    .A2(_3893_),
    .ZN(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8189_ (.A1(_3657_),
    .A2(_3888_),
    .B(_3894_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8190_ (.I(_3873_),
    .Z(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8191_ (.A1(\reg_file.reg_storage[6][19] ),
    .A2(_3893_),
    .ZN(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8192_ (.A1(_3667_),
    .A2(_3895_),
    .B(_3896_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8193_ (.A1(\reg_file.reg_storage[6][20] ),
    .A2(_3893_),
    .ZN(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8194_ (.A1(_3675_),
    .A2(_3895_),
    .B(_3897_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8195_ (.A1(\reg_file.reg_storage[6][21] ),
    .A2(_3893_),
    .ZN(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8196_ (.A1(_3682_),
    .A2(_3895_),
    .B(_3898_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8197_ (.A1(\reg_file.reg_storage[6][22] ),
    .A2(_3868_),
    .ZN(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8198_ (.A1(_3689_),
    .A2(_3895_),
    .B(_3899_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8199_ (.A1(\reg_file.reg_storage[6][23] ),
    .A2(_3868_),
    .ZN(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8200_ (.A1(_3696_),
    .A2(_3870_),
    .B(_3900_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8201_ (.A1(\reg_file.reg_storage[6][24] ),
    .A2(_3863_),
    .ZN(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8202_ (.A1(_3705_),
    .A2(_3862_),
    .B(_3901_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8203_ (.A1(\reg_file.reg_storage[6][25] ),
    .A2(_3863_),
    .ZN(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8204_ (.A1(_3710_),
    .A2(_3862_),
    .B(_3902_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8205_ (.I(_3860_),
    .Z(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8206_ (.A1(\reg_file.reg_storage[6][26] ),
    .A2(_3903_),
    .ZN(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8207_ (.A1(_3719_),
    .A2(_3862_),
    .B(_3904_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8208_ (.I(_3861_),
    .Z(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8209_ (.A1(\reg_file.reg_storage[6][27] ),
    .A2(_3903_),
    .ZN(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8210_ (.A1(_3726_),
    .A2(_3905_),
    .B(_3906_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8211_ (.A1(\reg_file.reg_storage[6][28] ),
    .A2(_3903_),
    .ZN(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8212_ (.A1(_3734_),
    .A2(_3905_),
    .B(_3907_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8213_ (.A1(\reg_file.reg_storage[6][29] ),
    .A2(_3903_),
    .ZN(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8214_ (.A1(_3740_),
    .A2(_3905_),
    .B(_3908_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8215_ (.A1(\reg_file.reg_storage[6][30] ),
    .A2(_3861_),
    .ZN(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8216_ (.A1(_3746_),
    .A2(_3905_),
    .B(_3909_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8217_ (.A1(\reg_file.reg_storage[6][31] ),
    .A2(_3861_),
    .ZN(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8218_ (.A1(_3751_),
    .A2(_3863_),
    .B(_3910_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8219_ (.I(_3420_),
    .Z(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8220_ (.I(_3911_),
    .Z(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8221_ (.A1(_3388_),
    .A2(_3754_),
    .ZN(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8222_ (.I(_3913_),
    .Z(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8223_ (.I(_3914_),
    .Z(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8224_ (.I(_3913_),
    .Z(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8225_ (.A1(\reg_file.reg_storage[7][0] ),
    .A2(_3916_),
    .ZN(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8226_ (.A1(_3912_),
    .A2(_3915_),
    .B(_3917_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8227_ (.I(_3442_),
    .Z(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8228_ (.I(_3918_),
    .Z(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8229_ (.A1(_3424_),
    .A2(_3761_),
    .ZN(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8230_ (.I(_3920_),
    .Z(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8231_ (.I(_3921_),
    .Z(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8232_ (.I(_3922_),
    .Z(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8233_ (.I(_3920_),
    .Z(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8234_ (.A1(\reg_file.reg_storage[7][1] ),
    .A2(_3924_),
    .ZN(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8235_ (.A1(_3919_),
    .A2(_3923_),
    .B(_3925_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8236_ (.I(_3454_),
    .Z(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8237_ (.I(_3920_),
    .Z(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _8238_ (.I(_3927_),
    .Z(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8239_ (.I0(\reg_file.reg_storage[7][2] ),
    .I1(_3926_),
    .S(_3928_),
    .Z(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8240_ (.I(_3929_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8241_ (.I(_3468_),
    .Z(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8242_ (.I0(\reg_file.reg_storage[7][3] ),
    .I1(_3930_),
    .S(_3928_),
    .Z(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8243_ (.I(_3931_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8244_ (.I(_3477_),
    .Z(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8245_ (.I(_3932_),
    .Z(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8246_ (.A1(\reg_file.reg_storage[7][4] ),
    .A2(_3924_),
    .ZN(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8247_ (.A1(_3933_),
    .A2(_3923_),
    .B(_3934_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8248_ (.I(_3489_),
    .Z(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8249_ (.I0(\reg_file.reg_storage[7][5] ),
    .I1(_3935_),
    .S(_3928_),
    .Z(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8250_ (.I(_3936_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8251_ (.I(_3501_),
    .Z(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8252_ (.I(_3937_),
    .Z(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8253_ (.A1(\reg_file.reg_storage[7][6] ),
    .A2(_3924_),
    .ZN(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8254_ (.A1(_3938_),
    .A2(_3923_),
    .B(_3939_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8255_ (.I(_3509_),
    .Z(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8256_ (.I(_3921_),
    .Z(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8257_ (.I0(\reg_file.reg_storage[7][7] ),
    .I1(_3940_),
    .S(_3941_),
    .Z(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8258_ (.I(_3942_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8259_ (.I(_3529_),
    .Z(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8260_ (.I0(\reg_file.reg_storage[7][8] ),
    .I1(_3943_),
    .S(_3941_),
    .Z(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8261_ (.I(_3944_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8262_ (.I(_3542_),
    .Z(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8263_ (.I(_3945_),
    .Z(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8264_ (.I(_3921_),
    .Z(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8265_ (.A1(\reg_file.reg_storage[7][9] ),
    .A2(_3947_),
    .ZN(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8266_ (.A1(_3946_),
    .A2(_3923_),
    .B(_3948_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8267_ (.I(_3555_),
    .Z(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8268_ (.I0(\reg_file.reg_storage[7][10] ),
    .I1(_3949_),
    .S(_3941_),
    .Z(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8269_ (.I(_3950_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8270_ (.I(_3566_),
    .Z(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8271_ (.I0(\reg_file.reg_storage[7][11] ),
    .I1(_3951_),
    .S(_3941_),
    .Z(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8272_ (.I(_3952_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8273_ (.I(_3583_),
    .Z(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8274_ (.I0(\reg_file.reg_storage[7][12] ),
    .I1(_3953_),
    .S(_3927_),
    .Z(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8275_ (.I(_3954_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8276_ (.I(_3596_),
    .Z(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8277_ (.I0(\reg_file.reg_storage[7][13] ),
    .I1(_3955_),
    .S(_3927_),
    .Z(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8278_ (.I(_3956_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8279_ (.I(_3610_),
    .Z(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8280_ (.I(_3957_),
    .Z(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8281_ (.I(_3922_),
    .Z(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8282_ (.A1(\reg_file.reg_storage[7][14] ),
    .A2(_3947_),
    .ZN(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8283_ (.A1(_3958_),
    .A2(_3959_),
    .B(_3960_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8284_ (.I(_3622_),
    .Z(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8285_ (.I0(\reg_file.reg_storage[7][15] ),
    .I1(_3961_),
    .S(_3927_),
    .Z(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8286_ (.I(_3962_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8287_ (.I(_3637_),
    .Z(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8288_ (.I(_3963_),
    .Z(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8289_ (.A1(\reg_file.reg_storage[7][16] ),
    .A2(_3947_),
    .ZN(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8290_ (.A1(_3964_),
    .A2(_3959_),
    .B(_3965_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8291_ (.I(_3648_),
    .Z(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8292_ (.I(_3966_),
    .Z(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8293_ (.A1(\reg_file.reg_storage[7][17] ),
    .A2(_3947_),
    .ZN(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8294_ (.A1(_3967_),
    .A2(_3959_),
    .B(_3968_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8295_ (.I(_3656_),
    .Z(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8296_ (.I(_3969_),
    .Z(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8297_ (.I(_3921_),
    .Z(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8298_ (.A1(\reg_file.reg_storage[7][18] ),
    .A2(_3971_),
    .ZN(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8299_ (.A1(_3970_),
    .A2(_3959_),
    .B(_3972_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8300_ (.I(_3666_),
    .Z(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8301_ (.I(_3973_),
    .Z(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8302_ (.I(_3928_),
    .Z(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8303_ (.A1(\reg_file.reg_storage[7][19] ),
    .A2(_3971_),
    .ZN(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8304_ (.A1(_3974_),
    .A2(_3975_),
    .B(_3976_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8305_ (.I(_3674_),
    .Z(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8306_ (.I(_3977_),
    .Z(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8307_ (.A1(\reg_file.reg_storage[7][20] ),
    .A2(_3971_),
    .ZN(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8308_ (.A1(_3978_),
    .A2(_3975_),
    .B(_3979_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8309_ (.I(_3681_),
    .Z(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8310_ (.I(_3980_),
    .Z(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8311_ (.A1(\reg_file.reg_storage[7][21] ),
    .A2(_3971_),
    .ZN(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8312_ (.A1(_3981_),
    .A2(_3975_),
    .B(_3982_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8313_ (.I(_3688_),
    .Z(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8314_ (.I(_3983_),
    .Z(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8315_ (.A1(\reg_file.reg_storage[7][22] ),
    .A2(_3922_),
    .ZN(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8316_ (.A1(_3984_),
    .A2(_3975_),
    .B(_3985_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8317_ (.I(_3695_),
    .Z(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8318_ (.I(_3986_),
    .Z(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8319_ (.A1(\reg_file.reg_storage[7][23] ),
    .A2(_3922_),
    .ZN(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8320_ (.A1(_3987_),
    .A2(_3924_),
    .B(_3988_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8321_ (.I(_3704_),
    .Z(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8322_ (.I(_3989_),
    .Z(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8323_ (.A1(\reg_file.reg_storage[7][24] ),
    .A2(_3916_),
    .ZN(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8324_ (.A1(_3990_),
    .A2(_3915_),
    .B(_3991_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8325_ (.I(_3709_),
    .Z(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8326_ (.I(_3992_),
    .Z(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8327_ (.A1(\reg_file.reg_storage[7][25] ),
    .A2(_3916_),
    .ZN(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8328_ (.A1(_3993_),
    .A2(_3915_),
    .B(_3994_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8329_ (.I(_3718_),
    .Z(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8330_ (.I(_3995_),
    .Z(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8331_ (.I(_3913_),
    .Z(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8332_ (.A1(\reg_file.reg_storage[7][26] ),
    .A2(_3997_),
    .ZN(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8333_ (.A1(_3996_),
    .A2(_3915_),
    .B(_3998_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8334_ (.I(_3725_),
    .Z(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8335_ (.I(_3999_),
    .Z(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8336_ (.I(_3914_),
    .Z(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8337_ (.A1(\reg_file.reg_storage[7][27] ),
    .A2(_3997_),
    .ZN(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8338_ (.A1(_4000_),
    .A2(_4001_),
    .B(_4002_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8339_ (.I(_3733_),
    .Z(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8340_ (.I(_4003_),
    .Z(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8341_ (.A1(\reg_file.reg_storage[7][28] ),
    .A2(_3997_),
    .ZN(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8342_ (.A1(_4004_),
    .A2(_4001_),
    .B(_4005_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8343_ (.I(_3739_),
    .Z(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8344_ (.I(_4006_),
    .Z(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8345_ (.A1(\reg_file.reg_storage[7][29] ),
    .A2(_3997_),
    .ZN(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8346_ (.A1(_4007_),
    .A2(_4001_),
    .B(_4008_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8347_ (.I(_3745_),
    .Z(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8348_ (.I(_4009_),
    .Z(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8349_ (.A1(\reg_file.reg_storage[7][30] ),
    .A2(_3914_),
    .ZN(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8350_ (.A1(_4010_),
    .A2(_4001_),
    .B(_4011_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8351_ (.I(_3750_),
    .Z(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8352_ (.I(_4012_),
    .Z(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8353_ (.A1(\reg_file.reg_storage[7][31] ),
    .A2(_3914_),
    .ZN(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8354_ (.A1(_4013_),
    .A2(_3916_),
    .B(_4014_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _8355_ (.A1(_1236_),
    .A2(_1106_),
    .ZN(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8356_ (.A1(_3809_),
    .A2(_4015_),
    .ZN(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8357_ (.I(_4016_),
    .Z(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8358_ (.I(_4017_),
    .Z(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8359_ (.I(_4016_),
    .Z(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8360_ (.A1(\reg_file.reg_storage[14][0] ),
    .A2(_4019_),
    .ZN(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8361_ (.A1(_3912_),
    .A2(_4018_),
    .B(_4020_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8362_ (.A1(_3760_),
    .A2(net2),
    .ZN(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8363_ (.A1(_3865_),
    .A2(_4021_),
    .ZN(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8364_ (.I(_4022_),
    .Z(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8365_ (.I(_4023_),
    .Z(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8366_ (.I(_4024_),
    .Z(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8367_ (.I(_4022_),
    .Z(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8368_ (.A1(\reg_file.reg_storage[14][1] ),
    .A2(_4026_),
    .ZN(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8369_ (.A1(_3919_),
    .A2(_4025_),
    .B(_4027_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8370_ (.I(_4022_),
    .Z(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8371_ (.I(_4028_),
    .Z(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8372_ (.I0(\reg_file.reg_storage[14][2] ),
    .I1(_3926_),
    .S(_4029_),
    .Z(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8373_ (.I(_4030_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8374_ (.I0(\reg_file.reg_storage[14][3] ),
    .I1(_3930_),
    .S(_4029_),
    .Z(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8375_ (.I(_4031_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8376_ (.A1(\reg_file.reg_storage[14][4] ),
    .A2(_4026_),
    .ZN(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8377_ (.A1(_3933_),
    .A2(_4025_),
    .B(_4032_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8378_ (.I0(\reg_file.reg_storage[14][5] ),
    .I1(_3935_),
    .S(_4029_),
    .Z(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8379_ (.I(_4033_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8380_ (.A1(\reg_file.reg_storage[14][6] ),
    .A2(_4026_),
    .ZN(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8381_ (.A1(_3938_),
    .A2(_4025_),
    .B(_4034_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8382_ (.I(_4023_),
    .Z(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8383_ (.I0(\reg_file.reg_storage[14][7] ),
    .I1(_3940_),
    .S(_4035_),
    .Z(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8384_ (.I(_4036_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8385_ (.I0(\reg_file.reg_storage[14][8] ),
    .I1(_3943_),
    .S(_4035_),
    .Z(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8386_ (.I(_4037_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8387_ (.I(_4023_),
    .Z(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8388_ (.A1(\reg_file.reg_storage[14][9] ),
    .A2(_4038_),
    .ZN(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8389_ (.A1(_3946_),
    .A2(_4025_),
    .B(_4039_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8390_ (.I0(\reg_file.reg_storage[14][10] ),
    .I1(_3949_),
    .S(_4035_),
    .Z(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8391_ (.I(_4040_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8392_ (.I0(\reg_file.reg_storage[14][11] ),
    .I1(_3951_),
    .S(_4035_),
    .Z(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8393_ (.I(_4041_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8394_ (.I0(\reg_file.reg_storage[14][12] ),
    .I1(_3953_),
    .S(_4028_),
    .Z(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8395_ (.I(_4042_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8396_ (.I0(\reg_file.reg_storage[14][13] ),
    .I1(_3955_),
    .S(_4028_),
    .Z(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8397_ (.I(_4043_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8398_ (.I(_4024_),
    .Z(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8399_ (.A1(\reg_file.reg_storage[14][14] ),
    .A2(_4038_),
    .ZN(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8400_ (.A1(_3958_),
    .A2(_4044_),
    .B(_4045_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8401_ (.I0(\reg_file.reg_storage[14][15] ),
    .I1(_3961_),
    .S(_4028_),
    .Z(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8402_ (.I(_4046_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8403_ (.A1(\reg_file.reg_storage[14][16] ),
    .A2(_4038_),
    .ZN(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8404_ (.A1(_3964_),
    .A2(_4044_),
    .B(_4047_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8405_ (.A1(\reg_file.reg_storage[14][17] ),
    .A2(_4038_),
    .ZN(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8406_ (.A1(_3967_),
    .A2(_4044_),
    .B(_4048_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8407_ (.I(_4023_),
    .Z(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8408_ (.A1(\reg_file.reg_storage[14][18] ),
    .A2(_4049_),
    .ZN(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8409_ (.A1(_3970_),
    .A2(_4044_),
    .B(_4050_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8410_ (.I(_4029_),
    .Z(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8411_ (.A1(\reg_file.reg_storage[14][19] ),
    .A2(_4049_),
    .ZN(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8412_ (.A1(_3974_),
    .A2(_4051_),
    .B(_4052_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8413_ (.A1(\reg_file.reg_storage[14][20] ),
    .A2(_4049_),
    .ZN(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8414_ (.A1(_3978_),
    .A2(_4051_),
    .B(_4053_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8415_ (.A1(\reg_file.reg_storage[14][21] ),
    .A2(_4049_),
    .ZN(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8416_ (.A1(_3981_),
    .A2(_4051_),
    .B(_4054_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8417_ (.A1(\reg_file.reg_storage[14][22] ),
    .A2(_4024_),
    .ZN(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8418_ (.A1(_3984_),
    .A2(_4051_),
    .B(_4055_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8419_ (.A1(\reg_file.reg_storage[14][23] ),
    .A2(_4024_),
    .ZN(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8420_ (.A1(_3987_),
    .A2(_4026_),
    .B(_4056_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8421_ (.A1(\reg_file.reg_storage[14][24] ),
    .A2(_4019_),
    .ZN(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8422_ (.A1(_3990_),
    .A2(_4018_),
    .B(_4057_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8423_ (.A1(\reg_file.reg_storage[14][25] ),
    .A2(_4019_),
    .ZN(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8424_ (.A1(_3993_),
    .A2(_4018_),
    .B(_4058_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8425_ (.I(_4016_),
    .Z(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8426_ (.A1(\reg_file.reg_storage[14][26] ),
    .A2(_4059_),
    .ZN(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8427_ (.A1(_3996_),
    .A2(_4018_),
    .B(_4060_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8428_ (.I(_4017_),
    .Z(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8429_ (.A1(\reg_file.reg_storage[14][27] ),
    .A2(_4059_),
    .ZN(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8430_ (.A1(_4000_),
    .A2(_4061_),
    .B(_4062_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8431_ (.A1(\reg_file.reg_storage[14][28] ),
    .A2(_4059_),
    .ZN(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8432_ (.A1(_4004_),
    .A2(_4061_),
    .B(_4063_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8433_ (.A1(\reg_file.reg_storage[14][29] ),
    .A2(_4059_),
    .ZN(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8434_ (.A1(_4007_),
    .A2(_4061_),
    .B(_4064_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8435_ (.A1(\reg_file.reg_storage[14][30] ),
    .A2(_4017_),
    .ZN(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8436_ (.A1(_4010_),
    .A2(_4061_),
    .B(_4065_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8437_ (.A1(\reg_file.reg_storage[14][31] ),
    .A2(_4017_),
    .ZN(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8438_ (.A1(_4013_),
    .A2(_4019_),
    .B(_4066_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8439_ (.A1(_3397_),
    .A2(_4015_),
    .ZN(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8440_ (.I(_4067_),
    .Z(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8441_ (.I(_4068_),
    .Z(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8442_ (.I(_4067_),
    .Z(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8443_ (.A1(\reg_file.reg_storage[13][0] ),
    .A2(_4070_),
    .ZN(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8444_ (.A1(_3912_),
    .A2(_4069_),
    .B(_4071_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8445_ (.A1(_3425_),
    .A2(_4021_),
    .ZN(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8446_ (.I(_4072_),
    .Z(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8447_ (.I(_4073_),
    .Z(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8448_ (.I(_4074_),
    .Z(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8449_ (.I(_4072_),
    .Z(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8450_ (.A1(\reg_file.reg_storage[13][1] ),
    .A2(_4076_),
    .ZN(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8451_ (.A1(_3919_),
    .A2(_4075_),
    .B(_4077_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8452_ (.I(_4072_),
    .Z(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8453_ (.I(_4078_),
    .Z(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8454_ (.I0(\reg_file.reg_storage[13][2] ),
    .I1(_3926_),
    .S(_4079_),
    .Z(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8455_ (.I(_4080_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8456_ (.I0(\reg_file.reg_storage[13][3] ),
    .I1(_3930_),
    .S(_4079_),
    .Z(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8457_ (.I(_4081_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8458_ (.A1(\reg_file.reg_storage[13][4] ),
    .A2(_4076_),
    .ZN(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8459_ (.A1(_3933_),
    .A2(_4075_),
    .B(_4082_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8460_ (.I0(\reg_file.reg_storage[13][5] ),
    .I1(_3935_),
    .S(_4079_),
    .Z(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8461_ (.I(_4083_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8462_ (.A1(\reg_file.reg_storage[13][6] ),
    .A2(_4076_),
    .ZN(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8463_ (.A1(_3938_),
    .A2(_4075_),
    .B(_4084_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8464_ (.I(_4073_),
    .Z(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8465_ (.I0(\reg_file.reg_storage[13][7] ),
    .I1(_3940_),
    .S(_4085_),
    .Z(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8466_ (.I(_4086_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8467_ (.I0(\reg_file.reg_storage[13][8] ),
    .I1(_3943_),
    .S(_4085_),
    .Z(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8468_ (.I(_4087_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8469_ (.I(_4073_),
    .Z(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8470_ (.A1(\reg_file.reg_storage[13][9] ),
    .A2(_4088_),
    .ZN(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8471_ (.A1(_3946_),
    .A2(_4075_),
    .B(_4089_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8472_ (.I0(\reg_file.reg_storage[13][10] ),
    .I1(_3949_),
    .S(_4085_),
    .Z(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8473_ (.I(_4090_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8474_ (.I0(\reg_file.reg_storage[13][11] ),
    .I1(_3951_),
    .S(_4085_),
    .Z(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8475_ (.I(_4091_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8476_ (.I0(\reg_file.reg_storage[13][12] ),
    .I1(_3953_),
    .S(_4078_),
    .Z(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8477_ (.I(_4092_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8478_ (.I0(\reg_file.reg_storage[13][13] ),
    .I1(_3955_),
    .S(_4078_),
    .Z(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8479_ (.I(_4093_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8480_ (.I(_4074_),
    .Z(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8481_ (.A1(\reg_file.reg_storage[13][14] ),
    .A2(_4088_),
    .ZN(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8482_ (.A1(_3958_),
    .A2(_4094_),
    .B(_4095_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8483_ (.I0(\reg_file.reg_storage[13][15] ),
    .I1(_3961_),
    .S(_4078_),
    .Z(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8484_ (.I(_4096_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8485_ (.A1(\reg_file.reg_storage[13][16] ),
    .A2(_4088_),
    .ZN(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8486_ (.A1(_3964_),
    .A2(_4094_),
    .B(_4097_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8487_ (.A1(\reg_file.reg_storage[13][17] ),
    .A2(_4088_),
    .ZN(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8488_ (.A1(_3967_),
    .A2(_4094_),
    .B(_4098_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8489_ (.I(_4073_),
    .Z(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8490_ (.A1(\reg_file.reg_storage[13][18] ),
    .A2(_4099_),
    .ZN(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8491_ (.A1(_3970_),
    .A2(_4094_),
    .B(_4100_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8492_ (.I(_4079_),
    .Z(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8493_ (.A1(\reg_file.reg_storage[13][19] ),
    .A2(_4099_),
    .ZN(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8494_ (.A1(_3974_),
    .A2(_4101_),
    .B(_4102_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8495_ (.A1(\reg_file.reg_storage[13][20] ),
    .A2(_4099_),
    .ZN(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8496_ (.A1(_3978_),
    .A2(_4101_),
    .B(_4103_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8497_ (.A1(\reg_file.reg_storage[13][21] ),
    .A2(_4099_),
    .ZN(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8498_ (.A1(_3981_),
    .A2(_4101_),
    .B(_4104_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8499_ (.A1(\reg_file.reg_storage[13][22] ),
    .A2(_4074_),
    .ZN(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8500_ (.A1(_3984_),
    .A2(_4101_),
    .B(_4105_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8501_ (.A1(\reg_file.reg_storage[13][23] ),
    .A2(_4074_),
    .ZN(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8502_ (.A1(_3987_),
    .A2(_4076_),
    .B(_4106_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8503_ (.A1(\reg_file.reg_storage[13][24] ),
    .A2(_4070_),
    .ZN(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8504_ (.A1(_3990_),
    .A2(_4069_),
    .B(_4107_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8505_ (.A1(\reg_file.reg_storage[13][25] ),
    .A2(_4070_),
    .ZN(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8506_ (.A1(_3993_),
    .A2(_4069_),
    .B(_4108_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8507_ (.I(_4067_),
    .Z(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8508_ (.A1(\reg_file.reg_storage[13][26] ),
    .A2(_4109_),
    .ZN(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8509_ (.A1(_3996_),
    .A2(_4069_),
    .B(_4110_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8510_ (.I(_4068_),
    .Z(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8511_ (.A1(\reg_file.reg_storage[13][27] ),
    .A2(_4109_),
    .ZN(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8512_ (.A1(_4000_),
    .A2(_4111_),
    .B(_4112_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8513_ (.A1(\reg_file.reg_storage[13][28] ),
    .A2(_4109_),
    .ZN(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8514_ (.A1(_4004_),
    .A2(_4111_),
    .B(_4113_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8515_ (.A1(\reg_file.reg_storage[13][29] ),
    .A2(_4109_),
    .ZN(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8516_ (.A1(_4007_),
    .A2(_4111_),
    .B(_4114_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8517_ (.A1(\reg_file.reg_storage[13][30] ),
    .A2(_4068_),
    .ZN(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8518_ (.A1(_4010_),
    .A2(_4111_),
    .B(_4115_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8519_ (.A1(\reg_file.reg_storage[13][31] ),
    .A2(_4068_),
    .ZN(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8520_ (.A1(_4013_),
    .A2(_4070_),
    .B(_4116_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8521_ (.A1(net31),
    .A2(_3390_),
    .ZN(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _8522_ (.A1(_3395_),
    .A2(_4117_),
    .Z(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8523_ (.A1(_4015_),
    .A2(_4118_),
    .ZN(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8524_ (.I(_4119_),
    .Z(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8525_ (.I(_4120_),
    .Z(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8526_ (.I(_4119_),
    .Z(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8527_ (.A1(\reg_file.reg_storage[12][0] ),
    .A2(_4122_),
    .ZN(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8528_ (.A1(_3912_),
    .A2(_4121_),
    .B(_4123_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _8529_ (.A1(_3395_),
    .A2(_4117_),
    .ZN(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8530_ (.A1(_4021_),
    .A2(_4124_),
    .ZN(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8531_ (.I(_4125_),
    .Z(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8532_ (.I(_4126_),
    .Z(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8533_ (.I(_4127_),
    .Z(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8534_ (.I(_4125_),
    .Z(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8535_ (.A1(\reg_file.reg_storage[12][1] ),
    .A2(_4129_),
    .ZN(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8536_ (.A1(_3919_),
    .A2(_4128_),
    .B(_4130_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8537_ (.I(_4125_),
    .Z(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8538_ (.I(_4131_),
    .Z(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8539_ (.I0(\reg_file.reg_storage[12][2] ),
    .I1(_3926_),
    .S(_4132_),
    .Z(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8540_ (.I(_4133_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8541_ (.I0(\reg_file.reg_storage[12][3] ),
    .I1(_3930_),
    .S(_4132_),
    .Z(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8542_ (.I(_4134_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8543_ (.A1(\reg_file.reg_storage[12][4] ),
    .A2(_4129_),
    .ZN(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8544_ (.A1(_3933_),
    .A2(_4128_),
    .B(_4135_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8545_ (.I0(\reg_file.reg_storage[12][5] ),
    .I1(_3935_),
    .S(_4132_),
    .Z(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8546_ (.I(_4136_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8547_ (.A1(\reg_file.reg_storage[12][6] ),
    .A2(_4129_),
    .ZN(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8548_ (.A1(_3938_),
    .A2(_4128_),
    .B(_4137_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8549_ (.I(_4126_),
    .Z(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8550_ (.I0(\reg_file.reg_storage[12][7] ),
    .I1(_3940_),
    .S(_4138_),
    .Z(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8551_ (.I(_4139_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8552_ (.I0(\reg_file.reg_storage[12][8] ),
    .I1(_3943_),
    .S(_4138_),
    .Z(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8553_ (.I(_4140_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8554_ (.I(_4126_),
    .Z(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8555_ (.A1(\reg_file.reg_storage[12][9] ),
    .A2(_4141_),
    .ZN(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8556_ (.A1(_3946_),
    .A2(_4128_),
    .B(_4142_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8557_ (.I0(\reg_file.reg_storage[12][10] ),
    .I1(_3949_),
    .S(_4138_),
    .Z(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8558_ (.I(_4143_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8559_ (.I0(\reg_file.reg_storage[12][11] ),
    .I1(_3951_),
    .S(_4138_),
    .Z(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8560_ (.I(_4144_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8561_ (.I0(\reg_file.reg_storage[12][12] ),
    .I1(_3953_),
    .S(_4131_),
    .Z(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8562_ (.I(_4145_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8563_ (.I0(\reg_file.reg_storage[12][13] ),
    .I1(_3955_),
    .S(_4131_),
    .Z(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8564_ (.I(_4146_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8565_ (.I(_4127_),
    .Z(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8566_ (.A1(\reg_file.reg_storage[12][14] ),
    .A2(_4141_),
    .ZN(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8567_ (.A1(_3958_),
    .A2(_4147_),
    .B(_4148_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8568_ (.I0(\reg_file.reg_storage[12][15] ),
    .I1(_3961_),
    .S(_4131_),
    .Z(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8569_ (.I(_4149_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8570_ (.A1(\reg_file.reg_storage[12][16] ),
    .A2(_4141_),
    .ZN(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8571_ (.A1(_3964_),
    .A2(_4147_),
    .B(_4150_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8572_ (.A1(\reg_file.reg_storage[12][17] ),
    .A2(_4141_),
    .ZN(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8573_ (.A1(_3967_),
    .A2(_4147_),
    .B(_4151_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8574_ (.I(_4126_),
    .Z(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8575_ (.A1(\reg_file.reg_storage[12][18] ),
    .A2(_4152_),
    .ZN(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8576_ (.A1(_3970_),
    .A2(_4147_),
    .B(_4153_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8577_ (.I(_4132_),
    .Z(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8578_ (.A1(\reg_file.reg_storage[12][19] ),
    .A2(_4152_),
    .ZN(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8579_ (.A1(_3974_),
    .A2(_4154_),
    .B(_4155_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8580_ (.A1(\reg_file.reg_storage[12][20] ),
    .A2(_4152_),
    .ZN(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8581_ (.A1(_3978_),
    .A2(_4154_),
    .B(_4156_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8582_ (.A1(\reg_file.reg_storage[12][21] ),
    .A2(_4152_),
    .ZN(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8583_ (.A1(_3981_),
    .A2(_4154_),
    .B(_4157_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8584_ (.A1(\reg_file.reg_storage[12][22] ),
    .A2(_4127_),
    .ZN(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8585_ (.A1(_3984_),
    .A2(_4154_),
    .B(_4158_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8586_ (.A1(\reg_file.reg_storage[12][23] ),
    .A2(_4127_),
    .ZN(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8587_ (.A1(_3987_),
    .A2(_4129_),
    .B(_4159_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8588_ (.A1(\reg_file.reg_storage[12][24] ),
    .A2(_4122_),
    .ZN(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8589_ (.A1(_3990_),
    .A2(_4121_),
    .B(_4160_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8590_ (.A1(\reg_file.reg_storage[12][25] ),
    .A2(_4122_),
    .ZN(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8591_ (.A1(_3993_),
    .A2(_4121_),
    .B(_4161_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8592_ (.I(_4119_),
    .Z(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8593_ (.A1(\reg_file.reg_storage[12][26] ),
    .A2(_4162_),
    .ZN(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8594_ (.A1(_3996_),
    .A2(_4121_),
    .B(_4163_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8595_ (.I(_4120_),
    .Z(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8596_ (.A1(\reg_file.reg_storage[12][27] ),
    .A2(_4162_),
    .ZN(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8597_ (.A1(_4000_),
    .A2(_4164_),
    .B(_4165_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8598_ (.A1(\reg_file.reg_storage[12][28] ),
    .A2(_4162_),
    .ZN(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8599_ (.A1(_4004_),
    .A2(_4164_),
    .B(_4166_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8600_ (.A1(\reg_file.reg_storage[12][29] ),
    .A2(_4162_),
    .ZN(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8601_ (.A1(_4007_),
    .A2(_4164_),
    .B(_4167_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8602_ (.A1(\reg_file.reg_storage[12][30] ),
    .A2(_4120_),
    .ZN(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8603_ (.A1(_4010_),
    .A2(_4164_),
    .B(_4168_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8604_ (.A1(\reg_file.reg_storage[12][31] ),
    .A2(_4120_),
    .ZN(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8605_ (.A1(_4013_),
    .A2(_4122_),
    .B(_4169_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8606_ (.I(_3420_),
    .Z(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _8607_ (.A1(_3760_),
    .A2(_1106_),
    .ZN(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8608_ (.A1(_4118_),
    .A2(_4171_),
    .ZN(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8609_ (.I(_4172_),
    .Z(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8610_ (.I(_4173_),
    .Z(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8611_ (.I(_4172_),
    .Z(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8612_ (.A1(\reg_file.reg_storage[8][0] ),
    .A2(_4175_),
    .ZN(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8613_ (.A1(_4170_),
    .A2(_4174_),
    .B(_4176_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8614_ (.I(_3442_),
    .Z(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _8615_ (.A1(_1236_),
    .A2(_3387_),
    .ZN(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8616_ (.A1(_4124_),
    .A2(_4178_),
    .ZN(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8617_ (.I(_4179_),
    .Z(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8618_ (.I(_4180_),
    .Z(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8619_ (.I(_4181_),
    .Z(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8620_ (.I(_4179_),
    .Z(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8621_ (.A1(\reg_file.reg_storage[8][1] ),
    .A2(_4183_),
    .ZN(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8622_ (.A1(_4177_),
    .A2(_4182_),
    .B(_4184_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8623_ (.I(_3454_),
    .Z(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8624_ (.I(_4179_),
    .Z(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8625_ (.I(_4186_),
    .Z(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8626_ (.I0(\reg_file.reg_storage[8][2] ),
    .I1(_4185_),
    .S(_4187_),
    .Z(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8627_ (.I(_4188_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8628_ (.I(_3468_),
    .Z(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8629_ (.I0(\reg_file.reg_storage[8][3] ),
    .I1(_4189_),
    .S(_4187_),
    .Z(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8630_ (.I(_4190_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8631_ (.I(_3477_),
    .Z(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8632_ (.A1(\reg_file.reg_storage[8][4] ),
    .A2(_4183_),
    .ZN(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8633_ (.A1(_4191_),
    .A2(_4182_),
    .B(_4192_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8634_ (.I(_3489_),
    .Z(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8635_ (.I0(\reg_file.reg_storage[8][5] ),
    .I1(_4193_),
    .S(_4187_),
    .Z(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8636_ (.I(_4194_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8637_ (.I(_3501_),
    .Z(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8638_ (.A1(\reg_file.reg_storage[8][6] ),
    .A2(_4183_),
    .ZN(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8639_ (.A1(_4195_),
    .A2(_4182_),
    .B(_4196_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8640_ (.I(_3509_),
    .Z(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8641_ (.I(_4180_),
    .Z(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8642_ (.I0(\reg_file.reg_storage[8][7] ),
    .I1(_4197_),
    .S(_4198_),
    .Z(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8643_ (.I(_4199_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8644_ (.I(_3529_),
    .Z(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8645_ (.I0(\reg_file.reg_storage[8][8] ),
    .I1(_4200_),
    .S(_4198_),
    .Z(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8646_ (.I(_4201_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8647_ (.I(_3542_),
    .Z(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8648_ (.I(_4180_),
    .Z(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8649_ (.A1(\reg_file.reg_storage[8][9] ),
    .A2(_4203_),
    .ZN(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8650_ (.A1(_4202_),
    .A2(_4182_),
    .B(_4204_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8651_ (.I(_3555_),
    .Z(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8652_ (.I0(\reg_file.reg_storage[8][10] ),
    .I1(_4205_),
    .S(_4198_),
    .Z(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8653_ (.I(_4206_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8654_ (.I(_3566_),
    .Z(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8655_ (.I0(\reg_file.reg_storage[8][11] ),
    .I1(_4207_),
    .S(_4198_),
    .Z(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8656_ (.I(_4208_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8657_ (.I(_3583_),
    .Z(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8658_ (.I0(\reg_file.reg_storage[8][12] ),
    .I1(_4209_),
    .S(_4186_),
    .Z(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8659_ (.I(_4210_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8660_ (.I(_3596_),
    .Z(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8661_ (.I0(\reg_file.reg_storage[8][13] ),
    .I1(_4211_),
    .S(_4186_),
    .Z(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8662_ (.I(_4212_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8663_ (.I(_3610_),
    .Z(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8664_ (.I(_4181_),
    .Z(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8665_ (.A1(\reg_file.reg_storage[8][14] ),
    .A2(_4203_),
    .ZN(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8666_ (.A1(_4213_),
    .A2(_4214_),
    .B(_4215_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8667_ (.I(_3622_),
    .Z(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8668_ (.I0(\reg_file.reg_storage[8][15] ),
    .I1(_4216_),
    .S(_4186_),
    .Z(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8669_ (.I(_4217_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8670_ (.I(_3637_),
    .Z(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8671_ (.A1(\reg_file.reg_storage[8][16] ),
    .A2(_4203_),
    .ZN(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8672_ (.A1(_4218_),
    .A2(_4214_),
    .B(_4219_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8673_ (.I(_3648_),
    .Z(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8674_ (.A1(\reg_file.reg_storage[8][17] ),
    .A2(_4203_),
    .ZN(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8675_ (.A1(_4220_),
    .A2(_4214_),
    .B(_4221_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8676_ (.I(_3656_),
    .Z(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8677_ (.I(_4180_),
    .Z(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8678_ (.A1(\reg_file.reg_storage[8][18] ),
    .A2(_4223_),
    .ZN(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8679_ (.A1(_4222_),
    .A2(_4214_),
    .B(_4224_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8680_ (.I(_3666_),
    .Z(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8681_ (.I(_4187_),
    .Z(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8682_ (.A1(\reg_file.reg_storage[8][19] ),
    .A2(_4223_),
    .ZN(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8683_ (.A1(_4225_),
    .A2(_4226_),
    .B(_4227_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8684_ (.I(_3674_),
    .Z(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8685_ (.A1(\reg_file.reg_storage[8][20] ),
    .A2(_4223_),
    .ZN(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8686_ (.A1(_4228_),
    .A2(_4226_),
    .B(_4229_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8687_ (.I(_3681_),
    .Z(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8688_ (.A1(\reg_file.reg_storage[8][21] ),
    .A2(_4223_),
    .ZN(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8689_ (.A1(_4230_),
    .A2(_4226_),
    .B(_4231_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8690_ (.I(_3688_),
    .Z(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8691_ (.A1(\reg_file.reg_storage[8][22] ),
    .A2(_4181_),
    .ZN(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8692_ (.A1(_4232_),
    .A2(_4226_),
    .B(_4233_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8693_ (.I(_3695_),
    .Z(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8694_ (.A1(\reg_file.reg_storage[8][23] ),
    .A2(_4181_),
    .ZN(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8695_ (.A1(_4234_),
    .A2(_4183_),
    .B(_4235_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8696_ (.I(_3704_),
    .Z(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8697_ (.A1(\reg_file.reg_storage[8][24] ),
    .A2(_4175_),
    .ZN(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8698_ (.A1(_4236_),
    .A2(_4174_),
    .B(_4237_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8699_ (.I(_3709_),
    .Z(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8700_ (.A1(\reg_file.reg_storage[8][25] ),
    .A2(_4175_),
    .ZN(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8701_ (.A1(_4238_),
    .A2(_4174_),
    .B(_4239_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8702_ (.I(_3718_),
    .Z(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8703_ (.I(_4172_),
    .Z(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8704_ (.A1(\reg_file.reg_storage[8][26] ),
    .A2(_4241_),
    .ZN(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8705_ (.A1(_4240_),
    .A2(_4174_),
    .B(_4242_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8706_ (.I(_3725_),
    .Z(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8707_ (.I(_4173_),
    .Z(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8708_ (.A1(\reg_file.reg_storage[8][27] ),
    .A2(_4241_),
    .ZN(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8709_ (.A1(_4243_),
    .A2(_4244_),
    .B(_4245_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8710_ (.I(_3733_),
    .Z(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8711_ (.A1(\reg_file.reg_storage[8][28] ),
    .A2(_4241_),
    .ZN(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8712_ (.A1(_4246_),
    .A2(_4244_),
    .B(_4247_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8713_ (.I(_3739_),
    .Z(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8714_ (.A1(\reg_file.reg_storage[8][29] ),
    .A2(_4241_),
    .ZN(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8715_ (.A1(_4248_),
    .A2(_4244_),
    .B(_4249_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8716_ (.I(_3745_),
    .Z(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8717_ (.A1(\reg_file.reg_storage[8][30] ),
    .A2(_4173_),
    .ZN(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8718_ (.A1(_4250_),
    .A2(_4244_),
    .B(_4251_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8719_ (.I(_3750_),
    .Z(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8720_ (.A1(\reg_file.reg_storage[8][31] ),
    .A2(_4173_),
    .ZN(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8721_ (.A1(_4252_),
    .A2(_4175_),
    .B(_4253_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8722_ (.A1(_3754_),
    .A2(_4171_),
    .ZN(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8723_ (.I(_4254_),
    .Z(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8724_ (.I(_4255_),
    .Z(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8725_ (.I(_4254_),
    .Z(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8726_ (.A1(\reg_file.reg_storage[11][0] ),
    .A2(_4257_),
    .ZN(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8727_ (.A1(_4170_),
    .A2(_4256_),
    .B(_4258_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8728_ (.A1(_3761_),
    .A2(_4178_),
    .ZN(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8729_ (.I(_4259_),
    .Z(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8730_ (.I(_4260_),
    .Z(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8731_ (.I(_4261_),
    .Z(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8732_ (.I(_4259_),
    .Z(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8733_ (.A1(\reg_file.reg_storage[11][1] ),
    .A2(_4263_),
    .ZN(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8734_ (.A1(_4177_),
    .A2(_4262_),
    .B(_4264_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8735_ (.I(_4259_),
    .Z(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8736_ (.I(_4265_),
    .Z(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8737_ (.I0(\reg_file.reg_storage[11][2] ),
    .I1(_4185_),
    .S(_4266_),
    .Z(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8738_ (.I(_4267_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8739_ (.I0(\reg_file.reg_storage[11][3] ),
    .I1(_4189_),
    .S(_4266_),
    .Z(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8740_ (.I(_4268_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8741_ (.A1(\reg_file.reg_storage[11][4] ),
    .A2(_4263_),
    .ZN(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8742_ (.A1(_4191_),
    .A2(_4262_),
    .B(_4269_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8743_ (.I0(\reg_file.reg_storage[11][5] ),
    .I1(_4193_),
    .S(_4266_),
    .Z(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8744_ (.I(_4270_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8745_ (.A1(\reg_file.reg_storage[11][6] ),
    .A2(_4263_),
    .ZN(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8746_ (.A1(_4195_),
    .A2(_4262_),
    .B(_4271_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8747_ (.I(_4260_),
    .Z(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8748_ (.I0(\reg_file.reg_storage[11][7] ),
    .I1(_4197_),
    .S(_4272_),
    .Z(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8749_ (.I(_4273_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8750_ (.I0(\reg_file.reg_storage[11][8] ),
    .I1(_4200_),
    .S(_4272_),
    .Z(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8751_ (.I(_4274_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8752_ (.I(_4260_),
    .Z(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8753_ (.A1(\reg_file.reg_storage[11][9] ),
    .A2(_4275_),
    .ZN(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8754_ (.A1(_4202_),
    .A2(_4262_),
    .B(_4276_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8755_ (.I0(\reg_file.reg_storage[11][10] ),
    .I1(_4205_),
    .S(_4272_),
    .Z(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8756_ (.I(_4277_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8757_ (.I0(\reg_file.reg_storage[11][11] ),
    .I1(_4207_),
    .S(_4272_),
    .Z(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8758_ (.I(_4278_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8759_ (.I0(\reg_file.reg_storage[11][12] ),
    .I1(_4209_),
    .S(_4265_),
    .Z(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8760_ (.I(_4279_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8761_ (.I0(\reg_file.reg_storage[11][13] ),
    .I1(_4211_),
    .S(_4265_),
    .Z(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8762_ (.I(_4280_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8763_ (.I(_4261_),
    .Z(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8764_ (.A1(\reg_file.reg_storage[11][14] ),
    .A2(_4275_),
    .ZN(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8765_ (.A1(_4213_),
    .A2(_4281_),
    .B(_4282_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8766_ (.I0(\reg_file.reg_storage[11][15] ),
    .I1(_4216_),
    .S(_4265_),
    .Z(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8767_ (.I(_4283_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8768_ (.A1(\reg_file.reg_storage[11][16] ),
    .A2(_4275_),
    .ZN(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8769_ (.A1(_4218_),
    .A2(_4281_),
    .B(_4284_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8770_ (.A1(\reg_file.reg_storage[11][17] ),
    .A2(_4275_),
    .ZN(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8771_ (.A1(_4220_),
    .A2(_4281_),
    .B(_4285_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8772_ (.I(_4260_),
    .Z(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8773_ (.A1(\reg_file.reg_storage[11][18] ),
    .A2(_4286_),
    .ZN(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8774_ (.A1(_4222_),
    .A2(_4281_),
    .B(_4287_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8775_ (.I(_4266_),
    .Z(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8776_ (.A1(\reg_file.reg_storage[11][19] ),
    .A2(_4286_),
    .ZN(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8777_ (.A1(_4225_),
    .A2(_4288_),
    .B(_4289_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8778_ (.A1(\reg_file.reg_storage[11][20] ),
    .A2(_4286_),
    .ZN(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8779_ (.A1(_4228_),
    .A2(_4288_),
    .B(_4290_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8780_ (.A1(\reg_file.reg_storage[11][21] ),
    .A2(_4286_),
    .ZN(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8781_ (.A1(_4230_),
    .A2(_4288_),
    .B(_4291_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8782_ (.A1(\reg_file.reg_storage[11][22] ),
    .A2(_4261_),
    .ZN(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8783_ (.A1(_4232_),
    .A2(_4288_),
    .B(_4292_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8784_ (.A1(\reg_file.reg_storage[11][23] ),
    .A2(_4261_),
    .ZN(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8785_ (.A1(_4234_),
    .A2(_4263_),
    .B(_4293_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8786_ (.A1(\reg_file.reg_storage[11][24] ),
    .A2(_4257_),
    .ZN(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8787_ (.A1(_4236_),
    .A2(_4256_),
    .B(_4294_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8788_ (.A1(\reg_file.reg_storage[11][25] ),
    .A2(_4257_),
    .ZN(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8789_ (.A1(_4238_),
    .A2(_4256_),
    .B(_4295_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8790_ (.I(_4254_),
    .Z(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8791_ (.A1(\reg_file.reg_storage[11][26] ),
    .A2(_4296_),
    .ZN(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8792_ (.A1(_4240_),
    .A2(_4256_),
    .B(_4297_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8793_ (.I(_4255_),
    .Z(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8794_ (.A1(\reg_file.reg_storage[11][27] ),
    .A2(_4296_),
    .ZN(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8795_ (.A1(_4243_),
    .A2(_4298_),
    .B(_4299_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8796_ (.A1(\reg_file.reg_storage[11][28] ),
    .A2(_4296_),
    .ZN(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8797_ (.A1(_4246_),
    .A2(_4298_),
    .B(_4300_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8798_ (.A1(\reg_file.reg_storage[11][29] ),
    .A2(_4296_),
    .ZN(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8799_ (.A1(_4248_),
    .A2(_4298_),
    .B(_4301_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8800_ (.A1(\reg_file.reg_storage[11][30] ),
    .A2(_4255_),
    .ZN(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8801_ (.A1(_4250_),
    .A2(_4298_),
    .B(_4302_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8802_ (.A1(\reg_file.reg_storage[11][31] ),
    .A2(_4255_),
    .ZN(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8803_ (.A1(_4252_),
    .A2(_4257_),
    .B(_4303_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8804_ (.A1(_3809_),
    .A2(_4171_),
    .ZN(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8805_ (.I(_4304_),
    .Z(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8806_ (.I(_4305_),
    .Z(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8807_ (.I(_4304_),
    .Z(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8808_ (.A1(\reg_file.reg_storage[10][0] ),
    .A2(_4307_),
    .ZN(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8809_ (.A1(_4170_),
    .A2(_4306_),
    .B(_4308_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8810_ (.A1(_3865_),
    .A2(_4178_),
    .ZN(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8811_ (.I(_4309_),
    .Z(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8812_ (.I(_4310_),
    .Z(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8813_ (.I(_4311_),
    .Z(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8814_ (.I(_4309_),
    .Z(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8815_ (.A1(\reg_file.reg_storage[10][1] ),
    .A2(_4313_),
    .ZN(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8816_ (.A1(_4177_),
    .A2(_4312_),
    .B(_4314_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8817_ (.I(_4309_),
    .Z(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8818_ (.I(_4315_),
    .Z(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8819_ (.I0(\reg_file.reg_storage[10][2] ),
    .I1(_4185_),
    .S(_4316_),
    .Z(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8820_ (.I(_4317_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8821_ (.I0(\reg_file.reg_storage[10][3] ),
    .I1(_4189_),
    .S(_4316_),
    .Z(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8822_ (.I(_4318_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8823_ (.A1(\reg_file.reg_storage[10][4] ),
    .A2(_4313_),
    .ZN(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8824_ (.A1(_4191_),
    .A2(_4312_),
    .B(_4319_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8825_ (.I0(\reg_file.reg_storage[10][5] ),
    .I1(_4193_),
    .S(_4316_),
    .Z(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8826_ (.I(_4320_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8827_ (.A1(\reg_file.reg_storage[10][6] ),
    .A2(_4313_),
    .ZN(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8828_ (.A1(_4195_),
    .A2(_4312_),
    .B(_4321_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8829_ (.I(_4310_),
    .Z(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8830_ (.I0(\reg_file.reg_storage[10][7] ),
    .I1(_4197_),
    .S(_4322_),
    .Z(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8831_ (.I(_4323_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8832_ (.I0(\reg_file.reg_storage[10][8] ),
    .I1(_4200_),
    .S(_4322_),
    .Z(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8833_ (.I(_4324_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8834_ (.I(_4310_),
    .Z(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8835_ (.A1(\reg_file.reg_storage[10][9] ),
    .A2(_4325_),
    .ZN(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8836_ (.A1(_4202_),
    .A2(_4312_),
    .B(_4326_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8837_ (.I0(\reg_file.reg_storage[10][10] ),
    .I1(_4205_),
    .S(_4322_),
    .Z(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8838_ (.I(_4327_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8839_ (.I0(\reg_file.reg_storage[10][11] ),
    .I1(_4207_),
    .S(_4322_),
    .Z(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8840_ (.I(_4328_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8841_ (.I0(\reg_file.reg_storage[10][12] ),
    .I1(_4209_),
    .S(_4315_),
    .Z(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8842_ (.I(_4329_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8843_ (.I0(\reg_file.reg_storage[10][13] ),
    .I1(_4211_),
    .S(_4315_),
    .Z(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8844_ (.I(_4330_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8845_ (.I(_4311_),
    .Z(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8846_ (.A1(\reg_file.reg_storage[10][14] ),
    .A2(_4325_),
    .ZN(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8847_ (.A1(_4213_),
    .A2(_4331_),
    .B(_4332_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8848_ (.I0(\reg_file.reg_storage[10][15] ),
    .I1(_4216_),
    .S(_4315_),
    .Z(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8849_ (.I(_4333_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8850_ (.A1(\reg_file.reg_storage[10][16] ),
    .A2(_4325_),
    .ZN(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8851_ (.A1(_4218_),
    .A2(_4331_),
    .B(_4334_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8852_ (.A1(\reg_file.reg_storage[10][17] ),
    .A2(_4325_),
    .ZN(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8853_ (.A1(_4220_),
    .A2(_4331_),
    .B(_4335_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8854_ (.I(_4310_),
    .Z(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8855_ (.A1(\reg_file.reg_storage[10][18] ),
    .A2(_4336_),
    .ZN(_4337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8856_ (.A1(_4222_),
    .A2(_4331_),
    .B(_4337_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8857_ (.I(_4316_),
    .Z(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8858_ (.A1(\reg_file.reg_storage[10][19] ),
    .A2(_4336_),
    .ZN(_4339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8859_ (.A1(_4225_),
    .A2(_4338_),
    .B(_4339_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8860_ (.A1(\reg_file.reg_storage[10][20] ),
    .A2(_4336_),
    .ZN(_4340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8861_ (.A1(_4228_),
    .A2(_4338_),
    .B(_4340_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8862_ (.A1(\reg_file.reg_storage[10][21] ),
    .A2(_4336_),
    .ZN(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8863_ (.A1(_4230_),
    .A2(_4338_),
    .B(_4341_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8864_ (.A1(\reg_file.reg_storage[10][22] ),
    .A2(_4311_),
    .ZN(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8865_ (.A1(_4232_),
    .A2(_4338_),
    .B(_4342_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8866_ (.A1(\reg_file.reg_storage[10][23] ),
    .A2(_4311_),
    .ZN(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8867_ (.A1(_4234_),
    .A2(_4313_),
    .B(_4343_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8868_ (.A1(\reg_file.reg_storage[10][24] ),
    .A2(_4307_),
    .ZN(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8869_ (.A1(_4236_),
    .A2(_4306_),
    .B(_4344_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8870_ (.A1(\reg_file.reg_storage[10][25] ),
    .A2(_4307_),
    .ZN(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8871_ (.A1(_4238_),
    .A2(_4306_),
    .B(_4345_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8872_ (.I(_4304_),
    .Z(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8873_ (.A1(\reg_file.reg_storage[10][26] ),
    .A2(_4346_),
    .ZN(_4347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8874_ (.A1(_4240_),
    .A2(_4306_),
    .B(_4347_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8875_ (.I(_4305_),
    .Z(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8876_ (.A1(\reg_file.reg_storage[10][27] ),
    .A2(_4346_),
    .ZN(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8877_ (.A1(_4243_),
    .A2(_4348_),
    .B(_4349_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8878_ (.A1(\reg_file.reg_storage[10][28] ),
    .A2(_4346_),
    .ZN(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8879_ (.A1(_4246_),
    .A2(_4348_),
    .B(_4350_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8880_ (.A1(\reg_file.reg_storage[10][29] ),
    .A2(_4346_),
    .ZN(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8881_ (.A1(_4248_),
    .A2(_4348_),
    .B(_4351_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8882_ (.A1(\reg_file.reg_storage[10][30] ),
    .A2(_4305_),
    .ZN(_4352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8883_ (.A1(_4250_),
    .A2(_4348_),
    .B(_4352_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8884_ (.A1(\reg_file.reg_storage[10][31] ),
    .A2(_4305_),
    .ZN(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8885_ (.A1(_4252_),
    .A2(_4307_),
    .B(_4353_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8886_ (.A1(_3397_),
    .A2(_4171_),
    .ZN(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8887_ (.I(_4354_),
    .Z(_4355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8888_ (.I(_4355_),
    .Z(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8889_ (.I(_4354_),
    .Z(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8890_ (.A1(\reg_file.reg_storage[9][0] ),
    .A2(_4357_),
    .ZN(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8891_ (.A1(_4170_),
    .A2(_4356_),
    .B(_4358_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8892_ (.A1(_3425_),
    .A2(_4178_),
    .ZN(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8893_ (.I(_4359_),
    .Z(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8894_ (.I(_4360_),
    .Z(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8895_ (.I(_4361_),
    .Z(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8896_ (.I(_4359_),
    .Z(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8897_ (.A1(\reg_file.reg_storage[9][1] ),
    .A2(_4363_),
    .ZN(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8898_ (.A1(_4177_),
    .A2(_4362_),
    .B(_4364_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8899_ (.I(_4359_),
    .Z(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _8900_ (.I(_4365_),
    .Z(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8901_ (.I0(\reg_file.reg_storage[9][2] ),
    .I1(_4185_),
    .S(_4366_),
    .Z(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8902_ (.I(_4367_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8903_ (.I0(\reg_file.reg_storage[9][3] ),
    .I1(_4189_),
    .S(_4366_),
    .Z(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8904_ (.I(_4368_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8905_ (.A1(\reg_file.reg_storage[9][4] ),
    .A2(_4363_),
    .ZN(_4369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8906_ (.A1(_4191_),
    .A2(_4362_),
    .B(_4369_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8907_ (.I0(\reg_file.reg_storage[9][5] ),
    .I1(_4193_),
    .S(_4366_),
    .Z(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8908_ (.I(_4370_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8909_ (.A1(\reg_file.reg_storage[9][6] ),
    .A2(_4363_),
    .ZN(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8910_ (.A1(_4195_),
    .A2(_4362_),
    .B(_4371_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8911_ (.I(_4360_),
    .Z(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8912_ (.I0(\reg_file.reg_storage[9][7] ),
    .I1(_4197_),
    .S(_4372_),
    .Z(_4373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8913_ (.I(_4373_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8914_ (.I0(\reg_file.reg_storage[9][8] ),
    .I1(_4200_),
    .S(_4372_),
    .Z(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8915_ (.I(_4374_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8916_ (.I(_4360_),
    .Z(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8917_ (.A1(\reg_file.reg_storage[9][9] ),
    .A2(_4375_),
    .ZN(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8918_ (.A1(_4202_),
    .A2(_4362_),
    .B(_4376_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8919_ (.I0(\reg_file.reg_storage[9][10] ),
    .I1(_4205_),
    .S(_4372_),
    .Z(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8920_ (.I(_4377_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8921_ (.I0(\reg_file.reg_storage[9][11] ),
    .I1(_4207_),
    .S(_4372_),
    .Z(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8922_ (.I(_4378_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8923_ (.I0(\reg_file.reg_storage[9][12] ),
    .I1(_4209_),
    .S(_4365_),
    .Z(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8924_ (.I(_4379_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8925_ (.I0(\reg_file.reg_storage[9][13] ),
    .I1(_4211_),
    .S(_4365_),
    .Z(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8926_ (.I(_4380_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8927_ (.I(_4361_),
    .Z(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8928_ (.A1(\reg_file.reg_storage[9][14] ),
    .A2(_4375_),
    .ZN(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8929_ (.A1(_4213_),
    .A2(_4381_),
    .B(_4382_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8930_ (.I0(\reg_file.reg_storage[9][15] ),
    .I1(_4216_),
    .S(_4365_),
    .Z(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8931_ (.I(_4383_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8932_ (.A1(\reg_file.reg_storage[9][16] ),
    .A2(_4375_),
    .ZN(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8933_ (.A1(_4218_),
    .A2(_4381_),
    .B(_4384_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8934_ (.A1(\reg_file.reg_storage[9][17] ),
    .A2(_4375_),
    .ZN(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8935_ (.A1(_4220_),
    .A2(_4381_),
    .B(_4385_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8936_ (.I(_4360_),
    .Z(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8937_ (.A1(\reg_file.reg_storage[9][18] ),
    .A2(_4386_),
    .ZN(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8938_ (.A1(_4222_),
    .A2(_4381_),
    .B(_4387_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8939_ (.I(_4366_),
    .Z(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8940_ (.A1(\reg_file.reg_storage[9][19] ),
    .A2(_4386_),
    .ZN(_4389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8941_ (.A1(_4225_),
    .A2(_4388_),
    .B(_4389_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8942_ (.A1(\reg_file.reg_storage[9][20] ),
    .A2(_4386_),
    .ZN(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8943_ (.A1(_4228_),
    .A2(_4388_),
    .B(_4390_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8944_ (.A1(\reg_file.reg_storage[9][21] ),
    .A2(_4386_),
    .ZN(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8945_ (.A1(_4230_),
    .A2(_4388_),
    .B(_4391_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8946_ (.A1(\reg_file.reg_storage[9][22] ),
    .A2(_4361_),
    .ZN(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8947_ (.A1(_4232_),
    .A2(_4388_),
    .B(_4392_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8948_ (.A1(\reg_file.reg_storage[9][23] ),
    .A2(_4361_),
    .ZN(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8949_ (.A1(_4234_),
    .A2(_4363_),
    .B(_4393_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8950_ (.A1(\reg_file.reg_storage[9][24] ),
    .A2(_4357_),
    .ZN(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8951_ (.A1(_4236_),
    .A2(_4356_),
    .B(_4394_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8952_ (.A1(\reg_file.reg_storage[9][25] ),
    .A2(_4357_),
    .ZN(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8953_ (.A1(_4238_),
    .A2(_4356_),
    .B(_4395_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8954_ (.I(_4354_),
    .Z(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8955_ (.A1(\reg_file.reg_storage[9][26] ),
    .A2(_4396_),
    .ZN(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8956_ (.A1(_4240_),
    .A2(_4356_),
    .B(_4397_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8957_ (.I(_4355_),
    .Z(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8958_ (.A1(\reg_file.reg_storage[9][27] ),
    .A2(_4396_),
    .ZN(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8959_ (.A1(_4243_),
    .A2(_4398_),
    .B(_4399_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8960_ (.A1(\reg_file.reg_storage[9][28] ),
    .A2(_4396_),
    .ZN(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8961_ (.A1(_4246_),
    .A2(_4398_),
    .B(_4400_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8962_ (.A1(\reg_file.reg_storage[9][29] ),
    .A2(_4396_),
    .ZN(_4401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8963_ (.A1(_4248_),
    .A2(_4398_),
    .B(_4401_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8964_ (.A1(\reg_file.reg_storage[9][30] ),
    .A2(_4355_),
    .ZN(_4402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8965_ (.A1(_4250_),
    .A2(_4398_),
    .B(_4402_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8966_ (.A1(\reg_file.reg_storage[9][31] ),
    .A2(_4355_),
    .ZN(_4403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8967_ (.A1(_4252_),
    .A2(_4357_),
    .B(_4403_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8968_ (.A1(_3397_),
    .A2(_3753_),
    .ZN(_4404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8969_ (.I(_4404_),
    .Z(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8970_ (.I(_4405_),
    .Z(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8971_ (.I(_4404_),
    .Z(_4407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8972_ (.A1(\reg_file.reg_storage[1][0] ),
    .A2(_4407_),
    .ZN(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8973_ (.A1(_3911_),
    .A2(_4406_),
    .B(_4408_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8974_ (.A1(_3760_),
    .A2(_3387_),
    .A3(_3425_),
    .ZN(_4409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8975_ (.I(_4409_),
    .Z(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8976_ (.I(_4410_),
    .Z(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8977_ (.I(_4409_),
    .Z(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8978_ (.A1(\reg_file.reg_storage[1][1] ),
    .A2(_4412_),
    .ZN(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8979_ (.A1(_3918_),
    .A2(_4411_),
    .B(_4413_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8980_ (.I(_4409_),
    .Z(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8981_ (.I(_4414_),
    .Z(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8982_ (.I0(\reg_file.reg_storage[1][2] ),
    .I1(_3455_),
    .S(_4415_),
    .Z(_4416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8983_ (.I(_4416_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8984_ (.I0(\reg_file.reg_storage[1][3] ),
    .I1(_3469_),
    .S(_4415_),
    .Z(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8985_ (.I(_4417_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8986_ (.A1(\reg_file.reg_storage[1][4] ),
    .A2(_4412_),
    .ZN(_4418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8987_ (.A1(_3932_),
    .A2(_4411_),
    .B(_4418_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8988_ (.I0(\reg_file.reg_storage[1][5] ),
    .I1(_3490_),
    .S(_4415_),
    .Z(_4419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8989_ (.I(_4419_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8990_ (.A1(\reg_file.reg_storage[1][6] ),
    .A2(_4412_),
    .ZN(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8991_ (.A1(_3937_),
    .A2(_4411_),
    .B(_4420_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8992_ (.I(_4414_),
    .Z(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8993_ (.I0(\reg_file.reg_storage[1][7] ),
    .I1(_3510_),
    .S(_4421_),
    .Z(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8994_ (.I(_4422_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8995_ (.I0(\reg_file.reg_storage[1][8] ),
    .I1(_3530_),
    .S(_4421_),
    .Z(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8996_ (.I(_4423_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8997_ (.I(_4414_),
    .Z(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8998_ (.A1(\reg_file.reg_storage[1][9] ),
    .A2(_4424_),
    .ZN(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8999_ (.A1(_3945_),
    .A2(_4411_),
    .B(_4425_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9000_ (.A1(_3556_),
    .A2(_4405_),
    .ZN(_4426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9001_ (.A1(_1197_),
    .A2(_4406_),
    .B(_4426_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9002_ (.I0(\reg_file.reg_storage[1][11] ),
    .I1(_3567_),
    .S(_4421_),
    .Z(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9003_ (.I(_4427_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9004_ (.I0(\reg_file.reg_storage[1][12] ),
    .I1(_3584_),
    .S(_4421_),
    .Z(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9005_ (.I(_4428_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9006_ (.I0(\reg_file.reg_storage[1][13] ),
    .I1(_3597_),
    .S(_4414_),
    .Z(_4429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9007_ (.I(_4429_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _9008_ (.I(_4410_),
    .Z(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9009_ (.A1(\reg_file.reg_storage[1][14] ),
    .A2(_4424_),
    .ZN(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9010_ (.A1(_3957_),
    .A2(_4430_),
    .B(_4431_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9011_ (.A1(_3623_),
    .A2(_4405_),
    .ZN(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9012_ (.A1(_1167_),
    .A2(_4406_),
    .B(_4432_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9013_ (.A1(\reg_file.reg_storage[1][16] ),
    .A2(_4424_),
    .ZN(_4433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9014_ (.A1(_3963_),
    .A2(_4430_),
    .B(_4433_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9015_ (.A1(\reg_file.reg_storage[1][17] ),
    .A2(_4424_),
    .ZN(_4434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9016_ (.A1(_3966_),
    .A2(_4430_),
    .B(_4434_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9017_ (.I(_4409_),
    .Z(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9018_ (.A1(\reg_file.reg_storage[1][18] ),
    .A2(_4435_),
    .ZN(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9019_ (.A1(_3969_),
    .A2(_4430_),
    .B(_4436_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9020_ (.I(_4415_),
    .Z(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9021_ (.A1(\reg_file.reg_storage[1][19] ),
    .A2(_4435_),
    .ZN(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9022_ (.A1(_3973_),
    .A2(_4437_),
    .B(_4438_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9023_ (.A1(\reg_file.reg_storage[1][20] ),
    .A2(_4435_),
    .ZN(_4439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9024_ (.A1(_3977_),
    .A2(_4437_),
    .B(_4439_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9025_ (.A1(\reg_file.reg_storage[1][21] ),
    .A2(_4435_),
    .ZN(_4440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9026_ (.A1(_3980_),
    .A2(_4437_),
    .B(_4440_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9027_ (.A1(\reg_file.reg_storage[1][22] ),
    .A2(_4410_),
    .ZN(_4441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9028_ (.A1(_3983_),
    .A2(_4437_),
    .B(_4441_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9029_ (.A1(\reg_file.reg_storage[1][23] ),
    .A2(_4410_),
    .ZN(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9030_ (.A1(_3986_),
    .A2(_4412_),
    .B(_4442_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _9031_ (.I(_4404_),
    .Z(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9032_ (.A1(\reg_file.reg_storage[1][24] ),
    .A2(_4443_),
    .ZN(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9033_ (.A1(_3989_),
    .A2(_4406_),
    .B(_4444_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _9034_ (.I(_4405_),
    .Z(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9035_ (.A1(\reg_file.reg_storage[1][25] ),
    .A2(_4443_),
    .ZN(_4446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9036_ (.A1(_3992_),
    .A2(_4445_),
    .B(_4446_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9037_ (.A1(\reg_file.reg_storage[1][26] ),
    .A2(_4443_),
    .ZN(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9038_ (.A1(_3995_),
    .A2(_4445_),
    .B(_4447_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9039_ (.A1(\reg_file.reg_storage[1][27] ),
    .A2(_4443_),
    .ZN(_4448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9040_ (.A1(_3999_),
    .A2(_4445_),
    .B(_4448_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _9041_ (.I(_4404_),
    .Z(_4449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9042_ (.A1(\reg_file.reg_storage[1][28] ),
    .A2(_4449_),
    .ZN(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9043_ (.A1(_4003_),
    .A2(_4445_),
    .B(_4450_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9044_ (.A1(\reg_file.reg_storage[1][29] ),
    .A2(_4449_),
    .ZN(_4451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9045_ (.A1(_4006_),
    .A2(_4407_),
    .B(_4451_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9046_ (.A1(\reg_file.reg_storage[1][30] ),
    .A2(_4449_),
    .ZN(_4452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9047_ (.A1(_4009_),
    .A2(_4407_),
    .B(_4452_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9048_ (.A1(\reg_file.reg_storage[1][31] ),
    .A2(_4449_),
    .ZN(_4453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9049_ (.A1(_4012_),
    .A2(_4407_),
    .B(_4453_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9050_ (.A1(_3388_),
    .A2(_4118_),
    .ZN(_4454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _9051_ (.I(_4454_),
    .Z(_4455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9052_ (.I(_4455_),
    .Z(_4456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9053_ (.I(_4454_),
    .Z(_4457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9054_ (.A1(\reg_file.reg_storage[4][0] ),
    .A2(_4457_),
    .ZN(_4458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9055_ (.A1(_3911_),
    .A2(_4456_),
    .B(_4458_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _9056_ (.A1(_3424_),
    .A2(_4124_),
    .ZN(_4459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9057_ (.I(_4459_),
    .Z(_4460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _9058_ (.I(_4460_),
    .Z(_4461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9059_ (.I(_4461_),
    .Z(_4462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9060_ (.I(_4459_),
    .Z(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9061_ (.A1(\reg_file.reg_storage[4][1] ),
    .A2(_4463_),
    .ZN(_4464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9062_ (.A1(_3918_),
    .A2(_4462_),
    .B(_4464_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _9063_ (.I(_4459_),
    .Z(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _9064_ (.I(_4465_),
    .Z(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9065_ (.I0(\reg_file.reg_storage[4][2] ),
    .I1(_3455_),
    .S(_4466_),
    .Z(_4467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9066_ (.I(_4467_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9067_ (.I0(\reg_file.reg_storage[4][3] ),
    .I1(_3469_),
    .S(_4466_),
    .Z(_4468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9068_ (.I(_4468_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9069_ (.A1(\reg_file.reg_storage[4][4] ),
    .A2(_4463_),
    .ZN(_4469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9070_ (.A1(_3932_),
    .A2(_4462_),
    .B(_4469_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9071_ (.I0(\reg_file.reg_storage[4][5] ),
    .I1(_3490_),
    .S(_4466_),
    .Z(_4470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9072_ (.I(_4470_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9073_ (.A1(\reg_file.reg_storage[4][6] ),
    .A2(_4463_),
    .ZN(_4471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9074_ (.A1(_3937_),
    .A2(_4462_),
    .B(_4471_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _9075_ (.I(_4460_),
    .Z(_4472_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9076_ (.I0(\reg_file.reg_storage[4][7] ),
    .I1(_3510_),
    .S(_4472_),
    .Z(_4473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9077_ (.I(_4473_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9078_ (.I0(\reg_file.reg_storage[4][8] ),
    .I1(_3530_),
    .S(_4472_),
    .Z(_4474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9079_ (.I(_4474_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9080_ (.I(_4460_),
    .Z(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9081_ (.A1(\reg_file.reg_storage[4][9] ),
    .A2(_4475_),
    .ZN(_4476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9082_ (.A1(_3945_),
    .A2(_4462_),
    .B(_4476_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9083_ (.I0(\reg_file.reg_storage[4][10] ),
    .I1(_3556_),
    .S(_4472_),
    .Z(_4477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9084_ (.I(_4477_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9085_ (.I0(\reg_file.reg_storage[4][11] ),
    .I1(_3567_),
    .S(_4472_),
    .Z(_4478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9086_ (.I(_4478_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9087_ (.I0(\reg_file.reg_storage[4][12] ),
    .I1(_3584_),
    .S(_4465_),
    .Z(_4479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9088_ (.I(_4479_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9089_ (.I0(\reg_file.reg_storage[4][13] ),
    .I1(_3597_),
    .S(_4465_),
    .Z(_4480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9090_ (.I(_4480_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _9091_ (.I(_4461_),
    .Z(_4481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9092_ (.A1(\reg_file.reg_storage[4][14] ),
    .A2(_4475_),
    .ZN(_4482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9093_ (.A1(_3957_),
    .A2(_4481_),
    .B(_4482_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9094_ (.I0(\reg_file.reg_storage[4][15] ),
    .I1(_3623_),
    .S(_4465_),
    .Z(_4483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9095_ (.I(_4483_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9096_ (.A1(\reg_file.reg_storage[4][16] ),
    .A2(_4475_),
    .ZN(_4484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9097_ (.A1(_3963_),
    .A2(_4481_),
    .B(_4484_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9098_ (.A1(\reg_file.reg_storage[4][17] ),
    .A2(_4475_),
    .ZN(_4485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9099_ (.A1(_3966_),
    .A2(_4481_),
    .B(_4485_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9100_ (.I(_4460_),
    .Z(_4486_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9101_ (.A1(\reg_file.reg_storage[4][18] ),
    .A2(_4486_),
    .ZN(_4487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9102_ (.A1(_3969_),
    .A2(_4481_),
    .B(_4487_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _9103_ (.I(_4466_),
    .Z(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9104_ (.A1(\reg_file.reg_storage[4][19] ),
    .A2(_4486_),
    .ZN(_4489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9105_ (.A1(_3973_),
    .A2(_4488_),
    .B(_4489_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9106_ (.A1(\reg_file.reg_storage[4][20] ),
    .A2(_4486_),
    .ZN(_4490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9107_ (.A1(_3977_),
    .A2(_4488_),
    .B(_4490_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9108_ (.A1(\reg_file.reg_storage[4][21] ),
    .A2(_4486_),
    .ZN(_4491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9109_ (.A1(_3980_),
    .A2(_4488_),
    .B(_4491_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9110_ (.A1(\reg_file.reg_storage[4][22] ),
    .A2(_4461_),
    .ZN(_4492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9111_ (.A1(_3983_),
    .A2(_4488_),
    .B(_4492_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9112_ (.A1(\reg_file.reg_storage[4][23] ),
    .A2(_4461_),
    .ZN(_4493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9113_ (.A1(_3986_),
    .A2(_4463_),
    .B(_4493_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9114_ (.A1(\reg_file.reg_storage[4][24] ),
    .A2(_4457_),
    .ZN(_4494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9115_ (.A1(_3989_),
    .A2(_4456_),
    .B(_4494_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9116_ (.A1(\reg_file.reg_storage[4][25] ),
    .A2(_4457_),
    .ZN(_4495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9117_ (.A1(_3992_),
    .A2(_4456_),
    .B(_4495_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _9118_ (.I(_4454_),
    .Z(_4496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9119_ (.A1(\reg_file.reg_storage[4][26] ),
    .A2(_4496_),
    .ZN(_4497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9120_ (.A1(_3995_),
    .A2(_4456_),
    .B(_4497_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9121_ (.I(_4455_),
    .Z(_4498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9122_ (.A1(\reg_file.reg_storage[4][27] ),
    .A2(_4496_),
    .ZN(_4499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9123_ (.A1(_3999_),
    .A2(_4498_),
    .B(_4499_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9124_ (.A1(\reg_file.reg_storage[4][28] ),
    .A2(_4496_),
    .ZN(_4500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9125_ (.A1(_4003_),
    .A2(_4498_),
    .B(_4500_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9126_ (.A1(\reg_file.reg_storage[4][29] ),
    .A2(_4496_),
    .ZN(_4501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9127_ (.A1(_4006_),
    .A2(_4498_),
    .B(_4501_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9128_ (.A1(\reg_file.reg_storage[4][30] ),
    .A2(_4455_),
    .ZN(_4502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9129_ (.A1(_4009_),
    .A2(_4498_),
    .B(_4502_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9130_ (.A1(\reg_file.reg_storage[4][31] ),
    .A2(_4455_),
    .ZN(_4503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9131_ (.A1(_4012_),
    .A2(_4457_),
    .B(_4503_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9132_ (.A1(_3754_),
    .A2(_4015_),
    .ZN(_4504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9133_ (.I(_4504_),
    .Z(_4505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _9134_ (.I(_4505_),
    .Z(_4506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _9135_ (.I(_4504_),
    .Z(_4507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9136_ (.A1(\reg_file.reg_storage[15][0] ),
    .A2(_4507_),
    .ZN(_4508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9137_ (.A1(_3911_),
    .A2(_4506_),
    .B(_4508_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9138_ (.A1(_3761_),
    .A2(_4021_),
    .ZN(_4509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _9139_ (.I(_4509_),
    .Z(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9140_ (.I(_4510_),
    .Z(_4511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9141_ (.I(_4511_),
    .Z(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9142_ (.I(_4509_),
    .Z(_4513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9143_ (.A1(\reg_file.reg_storage[15][1] ),
    .A2(_4513_),
    .ZN(_4514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9144_ (.A1(_3918_),
    .A2(_4512_),
    .B(_4514_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _9145_ (.I(_4509_),
    .Z(_4515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _9146_ (.I(_4515_),
    .Z(_4516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9147_ (.I0(\reg_file.reg_storage[15][2] ),
    .I1(_3455_),
    .S(_4516_),
    .Z(_4517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9148_ (.I(_4517_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9149_ (.I0(\reg_file.reg_storage[15][3] ),
    .I1(_3469_),
    .S(_4516_),
    .Z(_4518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9150_ (.I(_4518_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9151_ (.A1(\reg_file.reg_storage[15][4] ),
    .A2(_4513_),
    .ZN(_4519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9152_ (.A1(_3932_),
    .A2(_4512_),
    .B(_4519_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9153_ (.I0(\reg_file.reg_storage[15][5] ),
    .I1(_3490_),
    .S(_4516_),
    .Z(_4520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9154_ (.I(_4520_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9155_ (.A1(\reg_file.reg_storage[15][6] ),
    .A2(_4513_),
    .ZN(_4521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9156_ (.A1(_3937_),
    .A2(_4512_),
    .B(_4521_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _9157_ (.I(_4510_),
    .Z(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9158_ (.I0(\reg_file.reg_storage[15][7] ),
    .I1(_3510_),
    .S(_4522_),
    .Z(_4523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9159_ (.I(_4523_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9160_ (.I0(\reg_file.reg_storage[15][8] ),
    .I1(_3530_),
    .S(_4522_),
    .Z(_4524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9161_ (.I(_4524_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _9162_ (.I(_4510_),
    .Z(_4525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9163_ (.A1(\reg_file.reg_storage[15][9] ),
    .A2(_4525_),
    .ZN(_4526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9164_ (.A1(_3945_),
    .A2(_4512_),
    .B(_4526_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9165_ (.I0(\reg_file.reg_storage[15][10] ),
    .I1(_3556_),
    .S(_4522_),
    .Z(_4527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9166_ (.I(_4527_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9167_ (.I0(\reg_file.reg_storage[15][11] ),
    .I1(_3567_),
    .S(_4522_),
    .Z(_4528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9168_ (.I(_4528_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9169_ (.I0(\reg_file.reg_storage[15][12] ),
    .I1(_3584_),
    .S(_4515_),
    .Z(_4529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9170_ (.I(_4529_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9171_ (.I0(\reg_file.reg_storage[15][13] ),
    .I1(_3597_),
    .S(_4515_),
    .Z(_4530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9172_ (.I(_4530_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9173_ (.I(_4511_),
    .Z(_4531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9174_ (.A1(\reg_file.reg_storage[15][14] ),
    .A2(_4525_),
    .ZN(_4532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9175_ (.A1(_3957_),
    .A2(_4531_),
    .B(_4532_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _9176_ (.I0(\reg_file.reg_storage[15][15] ),
    .I1(_3623_),
    .S(_4515_),
    .Z(_4533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9177_ (.I(_4533_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9178_ (.A1(\reg_file.reg_storage[15][16] ),
    .A2(_4525_),
    .ZN(_4534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9179_ (.A1(_3963_),
    .A2(_4531_),
    .B(_4534_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9180_ (.A1(\reg_file.reg_storage[15][17] ),
    .A2(_4525_),
    .ZN(_4535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9181_ (.A1(_3966_),
    .A2(_4531_),
    .B(_4535_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9182_ (.I(_4510_),
    .Z(_4536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9183_ (.A1(\reg_file.reg_storage[15][18] ),
    .A2(_4536_),
    .ZN(_4537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9184_ (.A1(_3969_),
    .A2(_4531_),
    .B(_4537_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _9185_ (.I(_4516_),
    .Z(_4538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9186_ (.A1(\reg_file.reg_storage[15][19] ),
    .A2(_4536_),
    .ZN(_4539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9187_ (.A1(_3973_),
    .A2(_4538_),
    .B(_4539_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9188_ (.A1(\reg_file.reg_storage[15][20] ),
    .A2(_4536_),
    .ZN(_4540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9189_ (.A1(_3977_),
    .A2(_4538_),
    .B(_4540_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9190_ (.A1(\reg_file.reg_storage[15][21] ),
    .A2(_4536_),
    .ZN(_4541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9191_ (.A1(_3980_),
    .A2(_4538_),
    .B(_4541_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9192_ (.A1(\reg_file.reg_storage[15][22] ),
    .A2(_4511_),
    .ZN(_4542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9193_ (.A1(_3983_),
    .A2(_4538_),
    .B(_4542_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9194_ (.A1(\reg_file.reg_storage[15][23] ),
    .A2(_4511_),
    .ZN(_4543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9195_ (.A1(_3986_),
    .A2(_4513_),
    .B(_4543_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9196_ (.A1(\reg_file.reg_storage[15][24] ),
    .A2(_4507_),
    .ZN(_4544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9197_ (.A1(_3989_),
    .A2(_4506_),
    .B(_4544_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9198_ (.A1(\reg_file.reg_storage[15][25] ),
    .A2(_4507_),
    .ZN(_4545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9199_ (.A1(_3992_),
    .A2(_4506_),
    .B(_4545_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _9200_ (.I(_4504_),
    .Z(_4546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9201_ (.A1(\reg_file.reg_storage[15][26] ),
    .A2(_4546_),
    .ZN(_4547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9202_ (.A1(_3995_),
    .A2(_4506_),
    .B(_4547_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _9203_ (.I(_4505_),
    .Z(_4548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9204_ (.A1(\reg_file.reg_storage[15][27] ),
    .A2(_4546_),
    .ZN(_4549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9205_ (.A1(_3999_),
    .A2(_4548_),
    .B(_4549_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9206_ (.A1(\reg_file.reg_storage[15][28] ),
    .A2(_4546_),
    .ZN(_4550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9207_ (.A1(_4003_),
    .A2(_4548_),
    .B(_4550_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9208_ (.A1(\reg_file.reg_storage[15][29] ),
    .A2(_4546_),
    .ZN(_4551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9209_ (.A1(_4006_),
    .A2(_4548_),
    .B(_4551_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9210_ (.A1(\reg_file.reg_storage[15][30] ),
    .A2(_4505_),
    .ZN(_4552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9211_ (.A1(_4009_),
    .A2(_4548_),
    .B(_4552_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9212_ (.A1(\reg_file.reg_storage[15][31] ),
    .A2(_4505_),
    .ZN(_4553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9213_ (.A1(_4012_),
    .A2(_4507_),
    .B(_4553_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9214_ (.D(_0000_),
    .CLK(clknet_leaf_112_clk),
    .Q(\reg_file.reg_storage[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9215_ (.D(_0001_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9216_ (.D(_0002_),
    .CLK(clknet_leaf_129_clk),
    .Q(\reg_file.reg_storage[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9217_ (.D(_0003_),
    .CLK(clknet_leaf_126_clk),
    .Q(\reg_file.reg_storage[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9218_ (.D(_0004_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9219_ (.D(_0005_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9220_ (.D(_0006_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9221_ (.D(_0007_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9222_ (.D(_0008_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9223_ (.D(_0009_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9224_ (.D(_0010_),
    .CLK(clknet_4_10_0_clk),
    .Q(\reg_file.reg_storage[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9225_ (.D(_0011_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9226_ (.D(_0012_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9227_ (.D(_0013_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9228_ (.D(_0014_),
    .CLK(clknet_leaf_61_clk),
    .Q(\reg_file.reg_storage[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9229_ (.D(_0015_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9230_ (.D(_0016_),
    .CLK(clknet_leaf_60_clk),
    .Q(\reg_file.reg_storage[5][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9231_ (.D(_0017_),
    .CLK(clknet_4_10_0_clk),
    .Q(\reg_file.reg_storage[5][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9232_ (.D(_0018_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[5][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9233_ (.D(_0019_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[5][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9234_ (.D(_0020_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[5][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9235_ (.D(_0021_),
    .CLK(clknet_leaf_78_clk),
    .Q(\reg_file.reg_storage[5][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9236_ (.D(_0022_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[5][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9237_ (.D(_0023_),
    .CLK(clknet_leaf_119_clk),
    .Q(\reg_file.reg_storage[5][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9238_ (.D(_0024_),
    .CLK(clknet_leaf_112_clk),
    .Q(\reg_file.reg_storage[5][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9239_ (.D(_0025_),
    .CLK(clknet_leaf_114_clk),
    .Q(\reg_file.reg_storage[5][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9240_ (.D(_0026_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[5][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9241_ (.D(_0027_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[5][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9242_ (.D(_0028_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[5][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9243_ (.D(_0029_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[5][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9244_ (.D(_0030_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[5][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9245_ (.D(_0031_),
    .CLK(clknet_leaf_114_clk),
    .Q(\reg_file.reg_storage[5][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9246_ (.D(_0032_),
    .CLK(clknet_leaf_116_clk),
    .Q(\reg_file.reg_storage[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9247_ (.D(_0033_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9248_ (.D(_0034_),
    .CLK(clknet_leaf_132_clk),
    .Q(\reg_file.reg_storage[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9249_ (.D(_0035_),
    .CLK(clknet_leaf_130_clk),
    .Q(\reg_file.reg_storage[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9250_ (.D(_0036_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9251_ (.D(_0037_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9252_ (.D(_0038_),
    .CLK(clknet_4_7_0_clk),
    .Q(\reg_file.reg_storage[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9253_ (.D(_0039_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9254_ (.D(_0040_),
    .CLK(clknet_leaf_42_clk),
    .Q(\reg_file.reg_storage[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9255_ (.D(_0041_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9256_ (.D(_0042_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9257_ (.D(_0043_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9258_ (.D(_0044_),
    .CLK(clknet_leaf_14_clk),
    .Q(\reg_file.reg_storage[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9259_ (.D(_0045_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9260_ (.D(_0046_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9261_ (.D(_0047_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9262_ (.D(_0048_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[3][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9263_ (.D(_0049_),
    .CLK(clknet_leaf_58_clk),
    .Q(\reg_file.reg_storage[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9264_ (.D(_0050_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[3][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9265_ (.D(_0051_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9266_ (.D(_0052_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9267_ (.D(_0053_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9268_ (.D(_0054_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9269_ (.D(_0055_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[3][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9270_ (.D(_0056_),
    .CLK(clknet_leaf_116_clk),
    .Q(\reg_file.reg_storage[3][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9271_ (.D(_0057_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[3][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9272_ (.D(_0058_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[3][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9273_ (.D(_0059_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[3][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9274_ (.D(_0060_),
    .CLK(clknet_leaf_86_clk),
    .Q(\reg_file.reg_storage[3][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9275_ (.D(_0061_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[3][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9276_ (.D(_0062_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[3][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9277_ (.D(_0063_),
    .CLK(clknet_leaf_78_clk),
    .Q(\reg_file.reg_storage[3][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9278_ (.D(_0064_),
    .CLK(clknet_leaf_116_clk),
    .Q(\reg_file.reg_storage[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9279_ (.D(_0065_),
    .CLK(clknet_leaf_121_clk),
    .Q(\reg_file.reg_storage[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9280_ (.D(_0066_),
    .CLK(clknet_leaf_132_clk),
    .Q(\reg_file.reg_storage[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9281_ (.D(_0067_),
    .CLK(clknet_4_5_0_clk),
    .Q(\reg_file.reg_storage[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9282_ (.D(_0068_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9283_ (.D(_0069_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9284_ (.D(_0070_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9285_ (.D(_0071_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9286_ (.D(_0072_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9287_ (.D(_0073_),
    .CLK(clknet_4_3_0_clk),
    .Q(\reg_file.reg_storage[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9288_ (.D(_0074_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9289_ (.D(_0075_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9290_ (.D(_0076_),
    .CLK(clknet_leaf_15_clk),
    .Q(\reg_file.reg_storage[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9291_ (.D(_0077_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9292_ (.D(_0078_),
    .CLK(clknet_leaf_58_clk),
    .Q(\reg_file.reg_storage[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9293_ (.D(_0079_),
    .CLK(clknet_leaf_15_clk),
    .Q(\reg_file.reg_storage[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9294_ (.D(_0080_),
    .CLK(clknet_4_11_0_clk),
    .Q(\reg_file.reg_storage[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9295_ (.D(_0081_),
    .CLK(clknet_leaf_58_clk),
    .Q(\reg_file.reg_storage[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9296_ (.D(_0082_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9297_ (.D(_0083_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9298_ (.D(_0084_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9299_ (.D(_0085_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9300_ (.D(_0086_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9301_ (.D(_0087_),
    .CLK(clknet_leaf_24_clk),
    .Q(\reg_file.reg_storage[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9302_ (.D(_0088_),
    .CLK(clknet_leaf_116_clk),
    .Q(\reg_file.reg_storage[2][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9303_ (.D(_0089_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[2][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9304_ (.D(_0090_),
    .CLK(clknet_leaf_82_clk),
    .Q(\reg_file.reg_storage[2][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9305_ (.D(_0091_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[2][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9306_ (.D(_0092_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[2][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9307_ (.D(_0093_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[2][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9308_ (.D(_0094_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[2][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9309_ (.D(_0095_),
    .CLK(clknet_4_12_0_clk),
    .Q(\reg_file.reg_storage[2][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9310_ (.D(_0096_),
    .CLK(clknet_leaf_112_clk),
    .Q(\reg_file.reg_storage[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9311_ (.D(_0097_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9312_ (.D(_0098_),
    .CLK(clknet_leaf_133_clk),
    .Q(\reg_file.reg_storage[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9313_ (.D(_0099_),
    .CLK(clknet_leaf_130_clk),
    .Q(\reg_file.reg_storage[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9314_ (.D(_0100_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9315_ (.D(_0101_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9316_ (.D(_0102_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9317_ (.D(_0103_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9318_ (.D(_0104_),
    .CLK(clknet_leaf_42_clk),
    .Q(\reg_file.reg_storage[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9319_ (.D(_0105_),
    .CLK(clknet_leaf_34_clk),
    .Q(\reg_file.reg_storage[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9320_ (.D(_0106_),
    .CLK(clknet_leaf_49_clk),
    .Q(\reg_file.reg_storage[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9321_ (.D(_0107_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9322_ (.D(_0108_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9323_ (.D(_0109_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9324_ (.D(_0110_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9325_ (.D(_0111_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9326_ (.D(_0112_),
    .CLK(clknet_leaf_57_clk),
    .Q(\reg_file.reg_storage[6][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9327_ (.D(_0113_),
    .CLK(clknet_leaf_57_clk),
    .Q(\reg_file.reg_storage[6][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9328_ (.D(_0114_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[6][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9329_ (.D(_0115_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[6][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9330_ (.D(_0116_),
    .CLK(clknet_4_9_0_clk),
    .Q(\reg_file.reg_storage[6][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9331_ (.D(_0117_),
    .CLK(clknet_leaf_74_clk),
    .Q(\reg_file.reg_storage[6][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9332_ (.D(_0118_),
    .CLK(clknet_leaf_24_clk),
    .Q(\reg_file.reg_storage[6][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9333_ (.D(_0119_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9334_ (.D(_0120_),
    .CLK(clknet_leaf_114_clk),
    .Q(\reg_file.reg_storage[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9335_ (.D(_0121_),
    .CLK(clknet_leaf_114_clk),
    .Q(\reg_file.reg_storage[6][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9336_ (.D(_0122_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9337_ (.D(_0123_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[6][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9338_ (.D(_0124_),
    .CLK(clknet_leaf_95_clk),
    .Q(\reg_file.reg_storage[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9339_ (.D(_0125_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[6][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9340_ (.D(_0126_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[6][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9341_ (.D(_0127_),
    .CLK(clknet_leaf_115_clk),
    .Q(\reg_file.reg_storage[6][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9342_ (.D(_0128_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9343_ (.D(_0129_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9344_ (.D(_0130_),
    .CLK(clknet_leaf_134_clk),
    .Q(\reg_file.reg_storage[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9345_ (.D(_0131_),
    .CLK(clknet_leaf_130_clk),
    .Q(\reg_file.reg_storage[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9346_ (.D(_0132_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9347_ (.D(_0133_),
    .CLK(clknet_leaf_136_clk),
    .Q(\reg_file.reg_storage[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9348_ (.D(_0134_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9349_ (.D(_0135_),
    .CLK(clknet_leaf_40_clk),
    .Q(\reg_file.reg_storage[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9350_ (.D(_0136_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9351_ (.D(_0137_),
    .CLK(clknet_leaf_34_clk),
    .Q(\reg_file.reg_storage[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9352_ (.D(_0138_),
    .CLK(clknet_leaf_49_clk),
    .Q(\reg_file.reg_storage[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9353_ (.D(_0139_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9354_ (.D(_0140_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9355_ (.D(_0141_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9356_ (.D(_0142_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9357_ (.D(_0143_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9358_ (.D(_0144_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[7][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9359_ (.D(_0145_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[7][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9360_ (.D(_0146_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[7][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9361_ (.D(_0147_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[7][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9362_ (.D(_0148_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9363_ (.D(_0149_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9364_ (.D(_0150_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9365_ (.D(_0151_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9366_ (.D(_0152_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9367_ (.D(_0153_),
    .CLK(clknet_leaf_91_clk),
    .Q(\reg_file.reg_storage[7][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9368_ (.D(_0154_),
    .CLK(clknet_leaf_95_clk),
    .Q(\reg_file.reg_storage[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9369_ (.D(_0155_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[7][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9370_ (.D(_0156_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9371_ (.D(_0157_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[7][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9372_ (.D(_0158_),
    .CLK(clknet_leaf_90_clk),
    .Q(\reg_file.reg_storage[7][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9373_ (.D(_0159_),
    .CLK(clknet_leaf_91_clk),
    .Q(\reg_file.reg_storage[7][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9374_ (.D(_0160_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9375_ (.D(_0161_),
    .CLK(clknet_leaf_4_clk),
    .Q(\reg_file.reg_storage[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9376_ (.D(_0162_),
    .CLK(clknet_leaf_134_clk),
    .Q(\reg_file.reg_storage[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9377_ (.D(_0163_),
    .CLK(clknet_leaf_132_clk),
    .Q(\reg_file.reg_storage[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9378_ (.D(_0164_),
    .CLK(clknet_leaf_4_clk),
    .Q(\reg_file.reg_storage[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9379_ (.D(_0165_),
    .CLK(clknet_leaf_136_clk),
    .Q(\reg_file.reg_storage[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9380_ (.D(_0166_),
    .CLK(clknet_leaf_15_clk),
    .Q(\reg_file.reg_storage[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9381_ (.D(_0167_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9382_ (.D(_0168_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9383_ (.D(_0169_),
    .CLK(clknet_4_2_0_clk),
    .Q(\reg_file.reg_storage[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9384_ (.D(_0170_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9385_ (.D(_0171_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9386_ (.D(_0172_),
    .CLK(clknet_leaf_8_clk),
    .Q(\reg_file.reg_storage[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9387_ (.D(_0173_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9388_ (.D(_0174_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9389_ (.D(_0175_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9390_ (.D(_0176_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[14][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9391_ (.D(_0177_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[14][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9392_ (.D(_0178_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[14][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9393_ (.D(_0179_),
    .CLK(clknet_leaf_31_clk),
    .Q(\reg_file.reg_storage[14][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9394_ (.D(_0180_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[14][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9395_ (.D(_0181_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[14][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9396_ (.D(_0182_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[14][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9397_ (.D(_0183_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[14][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9398_ (.D(_0184_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9399_ (.D(_0185_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9400_ (.D(_0186_),
    .CLK(clknet_leaf_90_clk),
    .Q(\reg_file.reg_storage[14][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9401_ (.D(_0187_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9402_ (.D(_0188_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[14][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9403_ (.D(_0189_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[14][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9404_ (.D(_0190_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[14][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9405_ (.D(_0191_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[14][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9406_ (.D(_0192_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9407_ (.D(_0193_),
    .CLK(clknet_leaf_4_clk),
    .Q(\reg_file.reg_storage[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9408_ (.D(_0194_),
    .CLK(clknet_leaf_134_clk),
    .Q(\reg_file.reg_storage[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9409_ (.D(_0195_),
    .CLK(clknet_leaf_132_clk),
    .Q(\reg_file.reg_storage[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9410_ (.D(_0196_),
    .CLK(clknet_leaf_4_clk),
    .Q(\reg_file.reg_storage[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9411_ (.D(_0197_),
    .CLK(clknet_leaf_135_clk),
    .Q(\reg_file.reg_storage[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9412_ (.D(_0198_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9413_ (.D(_0199_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9414_ (.D(_0200_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9415_ (.D(_0201_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9416_ (.D(_0202_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9417_ (.D(_0203_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9418_ (.D(_0204_),
    .CLK(clknet_leaf_8_clk),
    .Q(\reg_file.reg_storage[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9419_ (.D(_0205_),
    .CLK(clknet_leaf_2_clk),
    .Q(\reg_file.reg_storage[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9420_ (.D(_0206_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9421_ (.D(_0207_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9422_ (.D(_0208_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[13][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9423_ (.D(_0209_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[13][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9424_ (.D(_0210_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[13][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9425_ (.D(_0211_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[13][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9426_ (.D(_0212_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[13][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9427_ (.D(_0213_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[13][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9428_ (.D(_0214_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[13][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9429_ (.D(_0215_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[13][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9430_ (.D(_0216_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9431_ (.D(_0217_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[13][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9432_ (.D(_0218_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9433_ (.D(_0219_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9434_ (.D(_0220_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[13][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9435_ (.D(_0221_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[13][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9436_ (.D(_0222_),
    .CLK(clknet_leaf_90_clk),
    .Q(\reg_file.reg_storage[13][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9437_ (.D(_0223_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[13][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9438_ (.D(_0224_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9439_ (.D(_0225_),
    .CLK(clknet_leaf_131_clk),
    .Q(\reg_file.reg_storage[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9440_ (.D(_0226_),
    .CLK(clknet_leaf_134_clk),
    .Q(\reg_file.reg_storage[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9441_ (.D(_0227_),
    .CLK(clknet_leaf_133_clk),
    .Q(\reg_file.reg_storage[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9442_ (.D(_0228_),
    .CLK(clknet_leaf_131_clk),
    .Q(\reg_file.reg_storage[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9443_ (.D(_0229_),
    .CLK(clknet_leaf_136_clk),
    .Q(\reg_file.reg_storage[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9444_ (.D(_0230_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9445_ (.D(_0231_),
    .CLK(clknet_leaf_40_clk),
    .Q(\reg_file.reg_storage[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9446_ (.D(_0232_),
    .CLK(clknet_leaf_42_clk),
    .Q(\reg_file.reg_storage[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9447_ (.D(_0233_),
    .CLK(clknet_leaf_34_clk),
    .Q(\reg_file.reg_storage[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9448_ (.D(_0234_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9449_ (.D(_0235_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9450_ (.D(_0236_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9451_ (.D(_0237_),
    .CLK(clknet_leaf_2_clk),
    .Q(\reg_file.reg_storage[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9452_ (.D(_0238_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9453_ (.D(_0239_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9454_ (.D(_0240_),
    .CLK(clknet_leaf_57_clk),
    .Q(\reg_file.reg_storage[12][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9455_ (.D(_0241_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[12][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9456_ (.D(_0242_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[12][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9457_ (.D(_0243_),
    .CLK(clknet_leaf_31_clk),
    .Q(\reg_file.reg_storage[12][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9458_ (.D(_0244_),
    .CLK(clknet_leaf_74_clk),
    .Q(\reg_file.reg_storage[12][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9459_ (.D(_0245_),
    .CLK(clknet_leaf_74_clk),
    .Q(\reg_file.reg_storage[12][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9460_ (.D(_0246_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[12][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9461_ (.D(_0247_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[12][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9462_ (.D(_0248_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[12][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9463_ (.D(_0249_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[12][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9464_ (.D(_0250_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[12][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9465_ (.D(_0251_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[12][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9466_ (.D(_0252_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[12][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9467_ (.D(_0253_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[12][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9468_ (.D(_0254_),
    .CLK(clknet_leaf_90_clk),
    .Q(\reg_file.reg_storage[12][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9469_ (.D(_0255_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[12][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9470_ (.D(_0256_),
    .CLK(clknet_leaf_109_clk),
    .Q(\reg_file.reg_storage[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9471_ (.D(_0257_),
    .CLK(clknet_leaf_120_clk),
    .Q(\reg_file.reg_storage[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9472_ (.D(_0258_),
    .CLK(clknet_leaf_127_clk),
    .Q(\reg_file.reg_storage[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9473_ (.D(_0259_),
    .CLK(clknet_leaf_126_clk),
    .Q(\reg_file.reg_storage[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9474_ (.D(_0260_),
    .CLK(clknet_leaf_120_clk),
    .Q(\reg_file.reg_storage[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9475_ (.D(_0261_),
    .CLK(clknet_leaf_135_clk),
    .Q(\reg_file.reg_storage[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9476_ (.D(_0262_),
    .CLK(clknet_leaf_120_clk),
    .Q(\reg_file.reg_storage[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9477_ (.D(_0263_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9478_ (.D(_0264_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9479_ (.D(_0265_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9480_ (.D(_0266_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9481_ (.D(_0267_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9482_ (.D(_0268_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9483_ (.D(_0269_),
    .CLK(clknet_leaf_2_clk),
    .Q(\reg_file.reg_storage[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9484_ (.D(_0270_),
    .CLK(clknet_leaf_65_clk),
    .Q(\reg_file.reg_storage[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9485_ (.D(_0271_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9486_ (.D(_0272_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[8][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9487_ (.D(_0273_),
    .CLK(clknet_leaf_64_clk),
    .Q(\reg_file.reg_storage[8][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9488_ (.D(_0274_),
    .CLK(clknet_leaf_68_clk),
    .Q(\reg_file.reg_storage[8][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9489_ (.D(_0275_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[8][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9490_ (.D(_0276_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[8][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9491_ (.D(_0277_),
    .CLK(clknet_leaf_77_clk),
    .Q(\reg_file.reg_storage[8][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9492_ (.D(_0278_),
    .CLK(clknet_leaf_117_clk),
    .Q(\reg_file.reg_storage[8][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9493_ (.D(_0279_),
    .CLK(clknet_leaf_119_clk),
    .Q(\reg_file.reg_storage[8][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9494_ (.D(_0280_),
    .CLK(clknet_leaf_108_clk),
    .Q(\reg_file.reg_storage[8][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9495_ (.D(_0281_),
    .CLK(clknet_leaf_108_clk),
    .Q(\reg_file.reg_storage[8][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9496_ (.D(_0282_),
    .CLK(clknet_leaf_106_clk),
    .Q(\reg_file.reg_storage[8][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9497_ (.D(_0283_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[8][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9498_ (.D(_0284_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[8][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9499_ (.D(_0285_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[8][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9500_ (.D(_0286_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[8][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9501_ (.D(_0287_),
    .CLK(clknet_leaf_107_clk),
    .Q(\reg_file.reg_storage[8][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9502_ (.D(_0288_),
    .CLK(clknet_leaf_109_clk),
    .Q(\reg_file.reg_storage[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9503_ (.D(_0289_),
    .CLK(clknet_leaf_123_clk),
    .Q(\reg_file.reg_storage[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9504_ (.D(_0290_),
    .CLK(clknet_leaf_128_clk),
    .Q(\reg_file.reg_storage[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9505_ (.D(_0291_),
    .CLK(clknet_leaf_127_clk),
    .Q(\reg_file.reg_storage[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9506_ (.D(_0292_),
    .CLK(clknet_leaf_121_clk),
    .Q(\reg_file.reg_storage[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9507_ (.D(_0293_),
    .CLK(clknet_leaf_135_clk),
    .Q(\reg_file.reg_storage[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9508_ (.D(_0294_),
    .CLK(clknet_leaf_121_clk),
    .Q(\reg_file.reg_storage[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9509_ (.D(_0295_),
    .CLK(clknet_leaf_40_clk),
    .Q(\reg_file.reg_storage[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9510_ (.D(_0296_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9511_ (.D(_0297_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9512_ (.D(_0298_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9513_ (.D(_0299_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9514_ (.D(_0300_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9515_ (.D(_0301_),
    .CLK(clknet_leaf_1_clk),
    .Q(\reg_file.reg_storage[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9516_ (.D(_0302_),
    .CLK(clknet_leaf_64_clk),
    .Q(\reg_file.reg_storage[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9517_ (.D(_0303_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9518_ (.D(_0304_),
    .CLK(clknet_leaf_60_clk),
    .Q(\reg_file.reg_storage[11][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9519_ (.D(_0305_),
    .CLK(clknet_leaf_64_clk),
    .Q(\reg_file.reg_storage[11][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9520_ (.D(_0306_),
    .CLK(clknet_leaf_68_clk),
    .Q(\reg_file.reg_storage[11][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9521_ (.D(_0307_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[11][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9522_ (.D(_0308_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[11][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9523_ (.D(_0309_),
    .CLK(clknet_leaf_76_clk),
    .Q(\reg_file.reg_storage[11][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9524_ (.D(_0310_),
    .CLK(clknet_leaf_24_clk),
    .Q(\reg_file.reg_storage[11][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9525_ (.D(_0311_),
    .CLK(clknet_leaf_119_clk),
    .Q(\reg_file.reg_storage[11][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9526_ (.D(_0312_),
    .CLK(clknet_leaf_109_clk),
    .Q(\reg_file.reg_storage[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9527_ (.D(_0313_),
    .CLK(clknet_leaf_108_clk),
    .Q(\reg_file.reg_storage[11][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9528_ (.D(_0314_),
    .CLK(clknet_leaf_106_clk),
    .Q(\reg_file.reg_storage[11][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9529_ (.D(_0315_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[11][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9530_ (.D(_0316_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[11][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9531_ (.D(_0317_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[11][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9532_ (.D(_0318_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[11][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9533_ (.D(_0319_),
    .CLK(clknet_leaf_108_clk),
    .Q(\reg_file.reg_storage[11][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9534_ (.D(_0320_),
    .CLK(clknet_4_13_0_clk),
    .Q(\reg_file.reg_storage[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9535_ (.D(_0321_),
    .CLK(clknet_leaf_123_clk),
    .Q(\reg_file.reg_storage[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9536_ (.D(_0322_),
    .CLK(clknet_leaf_128_clk),
    .Q(\reg_file.reg_storage[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9537_ (.D(_0323_),
    .CLK(clknet_leaf_127_clk),
    .Q(\reg_file.reg_storage[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9538_ (.D(_0324_),
    .CLK(clknet_leaf_121_clk),
    .Q(\reg_file.reg_storage[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9539_ (.D(_0325_),
    .CLK(clknet_4_4_0_clk),
    .Q(\reg_file.reg_storage[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9540_ (.D(_0326_),
    .CLK(clknet_leaf_121_clk),
    .Q(\reg_file.reg_storage[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9541_ (.D(_0327_),
    .CLK(clknet_leaf_40_clk),
    .Q(\reg_file.reg_storage[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9542_ (.D(_0328_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9543_ (.D(_0329_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9544_ (.D(_0330_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9545_ (.D(_0331_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9546_ (.D(_0332_),
    .CLK(clknet_leaf_2_clk),
    .Q(\reg_file.reg_storage[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9547_ (.D(_0333_),
    .CLK(clknet_leaf_1_clk),
    .Q(\reg_file.reg_storage[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9548_ (.D(_0334_),
    .CLK(clknet_leaf_65_clk),
    .Q(\reg_file.reg_storage[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9549_ (.D(_0335_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9550_ (.D(_0336_),
    .CLK(clknet_leaf_60_clk),
    .Q(\reg_file.reg_storage[10][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9551_ (.D(_0337_),
    .CLK(clknet_leaf_64_clk),
    .Q(\reg_file.reg_storage[10][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9552_ (.D(_0338_),
    .CLK(clknet_leaf_68_clk),
    .Q(\reg_file.reg_storage[10][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9553_ (.D(_0339_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[10][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9554_ (.D(_0340_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[10][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9555_ (.D(_0341_),
    .CLK(clknet_leaf_76_clk),
    .Q(\reg_file.reg_storage[10][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9556_ (.D(_0342_),
    .CLK(clknet_leaf_118_clk),
    .Q(\reg_file.reg_storage[10][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9557_ (.D(_0343_),
    .CLK(clknet_leaf_119_clk),
    .Q(\reg_file.reg_storage[10][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9558_ (.D(_0344_),
    .CLK(clknet_leaf_113_clk),
    .Q(\reg_file.reg_storage[10][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9559_ (.D(_0345_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[10][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9560_ (.D(_0346_),
    .CLK(clknet_leaf_106_clk),
    .Q(\reg_file.reg_storage[10][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9561_ (.D(_0347_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[10][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9562_ (.D(_0348_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[10][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9563_ (.D(_0349_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[10][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9564_ (.D(_0350_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[10][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9565_ (.D(_0351_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[10][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9566_ (.D(_0352_),
    .CLK(clknet_leaf_110_clk),
    .Q(\reg_file.reg_storage[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9567_ (.D(_0353_),
    .CLK(clknet_leaf_123_clk),
    .Q(\reg_file.reg_storage[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9568_ (.D(_0354_),
    .CLK(clknet_leaf_127_clk),
    .Q(\reg_file.reg_storage[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9569_ (.D(_0355_),
    .CLK(clknet_4_5_0_clk),
    .Q(\reg_file.reg_storage[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9570_ (.D(_0356_),
    .CLK(clknet_leaf_120_clk),
    .Q(\reg_file.reg_storage[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9571_ (.D(_0357_),
    .CLK(clknet_leaf_134_clk),
    .Q(\reg_file.reg_storage[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9572_ (.D(_0358_),
    .CLK(clknet_leaf_119_clk),
    .Q(\reg_file.reg_storage[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9573_ (.D(_0359_),
    .CLK(clknet_4_2_0_clk),
    .Q(\reg_file.reg_storage[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9574_ (.D(_0360_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9575_ (.D(_0361_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9576_ (.D(_0362_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9577_ (.D(_0363_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9578_ (.D(_0364_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9579_ (.D(_0365_),
    .CLK(clknet_leaf_1_clk),
    .Q(\reg_file.reg_storage[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9580_ (.D(_0366_),
    .CLK(clknet_leaf_65_clk),
    .Q(\reg_file.reg_storage[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9581_ (.D(_0367_),
    .CLK(clknet_leaf_14_clk),
    .Q(\reg_file.reg_storage[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9582_ (.D(_0368_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[9][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9583_ (.D(_0369_),
    .CLK(clknet_leaf_64_clk),
    .Q(\reg_file.reg_storage[9][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9584_ (.D(_0370_),
    .CLK(clknet_leaf_68_clk),
    .Q(\reg_file.reg_storage[9][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9585_ (.D(_0371_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[9][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9586_ (.D(_0372_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[9][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9587_ (.D(_0373_),
    .CLK(clknet_leaf_77_clk),
    .Q(\reg_file.reg_storage[9][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9588_ (.D(_0374_),
    .CLK(clknet_leaf_117_clk),
    .Q(\reg_file.reg_storage[9][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9589_ (.D(_0375_),
    .CLK(clknet_leaf_119_clk),
    .Q(\reg_file.reg_storage[9][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9590_ (.D(_0376_),
    .CLK(clknet_leaf_110_clk),
    .Q(\reg_file.reg_storage[9][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9591_ (.D(_0377_),
    .CLK(clknet_leaf_107_clk),
    .Q(\reg_file.reg_storage[9][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9592_ (.D(_0378_),
    .CLK(clknet_leaf_107_clk),
    .Q(\reg_file.reg_storage[9][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9593_ (.D(_0379_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[9][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9594_ (.D(_0380_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[9][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9595_ (.D(_0381_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[9][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9596_ (.D(_0382_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[9][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9597_ (.D(_0383_),
    .CLK(clknet_leaf_107_clk),
    .Q(\reg_file.reg_storage[9][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9598_ (.D(_0384_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9599_ (.D(_0385_),
    .CLK(clknet_4_7_0_clk),
    .Q(\reg_file.reg_storage[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9600_ (.D(_0386_),
    .CLK(clknet_leaf_129_clk),
    .Q(\reg_file.reg_storage[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9601_ (.D(_0387_),
    .CLK(clknet_leaf_126_clk),
    .Q(\reg_file.reg_storage[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9602_ (.D(_0388_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9603_ (.D(_0389_),
    .CLK(clknet_leaf_136_clk),
    .Q(\reg_file.reg_storage[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9604_ (.D(_0390_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9605_ (.D(_0391_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9606_ (.D(_0392_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9607_ (.D(_0393_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9608_ (.D(_0394_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9609_ (.D(_0395_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9610_ (.D(_0396_),
    .CLK(clknet_4_0_0_clk),
    .Q(\reg_file.reg_storage[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9611_ (.D(_0397_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9612_ (.D(_0398_),
    .CLK(clknet_leaf_63_clk),
    .Q(\reg_file.reg_storage[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9613_ (.D(_0399_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9614_ (.D(_0400_),
    .CLK(clknet_leaf_62_clk),
    .Q(\reg_file.reg_storage[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9615_ (.D(_0401_),
    .CLK(clknet_leaf_63_clk),
    .Q(\reg_file.reg_storage[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9616_ (.D(_0402_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9617_ (.D(_0403_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9618_ (.D(_0404_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9619_ (.D(_0405_),
    .CLK(clknet_leaf_76_clk),
    .Q(\reg_file.reg_storage[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9620_ (.D(_0406_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9621_ (.D(_0407_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9622_ (.D(_0408_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[1][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9623_ (.D(_0409_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[1][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9624_ (.D(_0410_),
    .CLK(clknet_leaf_82_clk),
    .Q(\reg_file.reg_storage[1][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9625_ (.D(_0411_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[1][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9626_ (.D(_0412_),
    .CLK(clknet_4_14_0_clk),
    .Q(\reg_file.reg_storage[1][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9627_ (.D(_0413_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[1][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9628_ (.D(_0414_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[1][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9629_ (.D(_0415_),
    .CLK(clknet_leaf_82_clk),
    .Q(\reg_file.reg_storage[1][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9630_ (.D(_0416_),
    .CLK(clknet_leaf_112_clk),
    .Q(\reg_file.reg_storage[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9631_ (.D(_0417_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9632_ (.D(_0418_),
    .CLK(clknet_leaf_129_clk),
    .Q(\reg_file.reg_storage[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9633_ (.D(_0419_),
    .CLK(clknet_leaf_126_clk),
    .Q(\reg_file.reg_storage[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9634_ (.D(_0420_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9635_ (.D(_0421_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9636_ (.D(_0422_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9637_ (.D(_0423_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9638_ (.D(_0424_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9639_ (.D(_0425_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9640_ (.D(_0426_),
    .CLK(clknet_leaf_58_clk),
    .Q(\reg_file.reg_storage[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9641_ (.D(_0427_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9642_ (.D(_0428_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9643_ (.D(_0429_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9644_ (.D(_0430_),
    .CLK(clknet_leaf_62_clk),
    .Q(\reg_file.reg_storage[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9645_ (.D(_0431_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9646_ (.D(_0432_),
    .CLK(clknet_leaf_61_clk),
    .Q(\reg_file.reg_storage[4][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9647_ (.D(_0433_),
    .CLK(clknet_leaf_62_clk),
    .Q(\reg_file.reg_storage[4][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9648_ (.D(_0434_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[4][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9649_ (.D(_0435_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[4][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9650_ (.D(_0436_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[4][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9651_ (.D(_0437_),
    .CLK(clknet_leaf_78_clk),
    .Q(\reg_file.reg_storage[4][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9652_ (.D(_0438_),
    .CLK(clknet_leaf_24_clk),
    .Q(\reg_file.reg_storage[4][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9653_ (.D(_0439_),
    .CLK(clknet_leaf_118_clk),
    .Q(\reg_file.reg_storage[4][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9654_ (.D(_0440_),
    .CLK(clknet_leaf_113_clk),
    .Q(\reg_file.reg_storage[4][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9655_ (.D(_0441_),
    .CLK(clknet_leaf_115_clk),
    .Q(\reg_file.reg_storage[4][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9656_ (.D(_0442_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[4][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9657_ (.D(_0443_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[4][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9658_ (.D(_0444_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[4][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9659_ (.D(_0445_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[4][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9660_ (.D(_0446_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[4][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9661_ (.D(_0447_),
    .CLK(clknet_leaf_115_clk),
    .Q(\reg_file.reg_storage[4][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9662_ (.D(_0448_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9663_ (.D(_0449_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9664_ (.D(_0450_),
    .CLK(clknet_leaf_133_clk),
    .Q(\reg_file.reg_storage[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9665_ (.D(_0451_),
    .CLK(clknet_leaf_133_clk),
    .Q(\reg_file.reg_storage[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9666_ (.D(_0452_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9667_ (.D(_0453_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9668_ (.D(_0454_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9669_ (.D(_0455_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9670_ (.D(_0456_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9671_ (.D(_0457_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9672_ (.D(_0458_),
    .CLK(clknet_leaf_49_clk),
    .Q(\reg_file.reg_storage[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9673_ (.D(_0459_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9674_ (.D(_0460_),
    .CLK(clknet_leaf_8_clk),
    .Q(\reg_file.reg_storage[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9675_ (.D(_0461_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9676_ (.D(_0462_),
    .CLK(clknet_leaf_62_clk),
    .Q(\reg_file.reg_storage[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9677_ (.D(_0463_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9678_ (.D(_0464_),
    .CLK(clknet_leaf_62_clk),
    .Q(\reg_file.reg_storage[15][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9679_ (.D(_0465_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[15][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9680_ (.D(_0466_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[15][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9681_ (.D(_0467_),
    .CLK(clknet_leaf_31_clk),
    .Q(\reg_file.reg_storage[15][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9682_ (.D(_0468_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[15][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9683_ (.D(_0469_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[15][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9684_ (.D(_0470_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[15][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9685_ (.D(_0471_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[15][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9686_ (.D(_0472_),
    .CLK(clknet_leaf_86_clk),
    .Q(\reg_file.reg_storage[15][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9687_ (.D(_0473_),
    .CLK(clknet_leaf_92_clk),
    .Q(\reg_file.reg_storage[15][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9688_ (.D(_0474_),
    .CLK(clknet_leaf_92_clk),
    .Q(\reg_file.reg_storage[15][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9689_ (.D(_0475_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[15][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9690_ (.D(_0476_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[15][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9691_ (.D(_0477_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[15][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9692_ (.D(_0478_),
    .CLK(clknet_leaf_91_clk),
    .Q(\reg_file.reg_storage[15][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9693_ (.D(_0479_),
    .CLK(clknet_leaf_92_clk),
    .Q(\reg_file.reg_storage[15][31] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_116_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_leaf_117_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_leaf_118_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_leaf_119_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_leaf_120_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_leaf_121_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_123_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_126_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_128_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_129_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_130_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_131_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_131_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_132_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_133_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_133_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_134_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_135_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_136_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_136_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1 (.I(inst[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(inst[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(inst[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input12 (.I(inst[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input13 (.I(inst[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input14 (.I(inst[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(inst[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input16 (.I(inst[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input17 (.I(inst[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input18 (.I(inst[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input19 (.I(inst[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input2 (.I(inst[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input20 (.I(inst[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input21 (.I(inst[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input22 (.I(inst[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input23 (.I(inst[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input24 (.I(inst[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input25 (.I(inst[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input26 (.I(inst[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input27 (.I(inst[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input28 (.I(inst[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input29 (.I(inst[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input3 (.I(inst[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input30 (.I(inst[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input31 (.I(inst[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input32 (.I(inst[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(mem_ld_dat[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(mem_ld_dat[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(mem_ld_dat[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(mem_ld_dat[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(mem_ld_dat[13]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(mem_ld_dat[14]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(mem_ld_dat[15]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input4 (.I(inst[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(mem_ld_dat[16]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input41 (.I(mem_ld_dat[17]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(mem_ld_dat[18]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input43 (.I(mem_ld_dat[19]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(mem_ld_dat[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input45 (.I(mem_ld_dat[20]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input46 (.I(mem_ld_dat[21]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input47 (.I(mem_ld_dat[22]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input48 (.I(mem_ld_dat[23]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input49 (.I(mem_ld_dat[24]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input5 (.I(inst[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input50 (.I(mem_ld_dat[25]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(mem_ld_dat[26]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(mem_ld_dat[27]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(mem_ld_dat[28]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(mem_ld_dat[29]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(mem_ld_dat[2]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input56 (.I(mem_ld_dat[30]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(mem_ld_dat[31]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(mem_ld_dat[3]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input59 (.I(mem_ld_dat[4]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input6 (.I(inst[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input60 (.I(mem_ld_dat[5]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input61 (.I(mem_ld_dat[6]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input62 (.I(mem_ld_dat[7]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input63 (.I(mem_ld_dat[8]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input64 (.I(mem_ld_dat[9]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input65 (.I(pc[0]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input66 (.I(pc[10]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input67 (.I(pc[11]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(pc[12]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input69 (.I(pc[13]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(inst[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input70 (.I(pc[14]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input71 (.I(pc[15]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input72 (.I(pc[16]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input73 (.I(pc[17]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input74 (.I(pc[18]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input75 (.I(pc[19]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input76 (.I(pc[1]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input77 (.I(pc[20]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input78 (.I(pc[21]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input79 (.I(pc[22]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input8 (.I(inst[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input80 (.I(pc[23]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input81 (.I(pc[24]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input82 (.I(pc[25]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input83 (.I(pc[26]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input84 (.I(pc[27]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input85 (.I(pc[28]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input86 (.I(pc[29]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input87 (.I(pc[2]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input88 (.I(pc[30]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input89 (.I(pc[31]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input9 (.I(inst[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input90 (.I(pc[3]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input91 (.I(pc[4]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input92 (.I(pc[5]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input93 (.I(pc[6]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input94 (.I(pc[7]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input95 (.I(pc[8]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input96 (.I(pc[9]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 load_slew1 (.I(_2413_),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output100 (.I(net100),
    .Z(mem_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output101 (.I(net101),
    .Z(mem_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output102 (.I(net102),
    .Z(mem_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output103 (.I(net103),
    .Z(mem_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output104 (.I(net104),
    .Z(mem_addr[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output105 (.I(net105),
    .Z(mem_addr[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output106 (.I(net106),
    .Z(mem_addr[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output107 (.I(net107),
    .Z(mem_addr[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output108 (.I(net108),
    .Z(mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output109 (.I(net109),
    .Z(mem_addr[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output110 (.I(net110),
    .Z(mem_addr[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output111 (.I(net111),
    .Z(mem_addr[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output112 (.I(net112),
    .Z(mem_addr[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output113 (.I(net113),
    .Z(mem_addr[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output114 (.I(net114),
    .Z(mem_addr[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output115 (.I(net115),
    .Z(mem_addr[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output116 (.I(net116),
    .Z(mem_addr[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output117 (.I(net117),
    .Z(mem_addr[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output118 (.I(net118),
    .Z(mem_addr[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output119 (.I(net119),
    .Z(mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output120 (.I(net120),
    .Z(mem_addr[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output121 (.I(net211),
    .Z(mem_addr[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output122 (.I(net122),
    .Z(mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output123 (.I(net123),
    .Z(mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output124 (.I(net124),
    .Z(mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output125 (.I(net125),
    .Z(mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output126 (.I(net126),
    .Z(mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output127 (.I(net127),
    .Z(mem_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output128 (.I(net128),
    .Z(mem_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output129 (.I(net129),
    .Z(mem_ld_en));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output130 (.I(net130),
    .Z(mem_ld_mask[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output131 (.I(net131),
    .Z(mem_ld_mask[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output132 (.I(net132),
    .Z(mem_ld_mask[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output133 (.I(net133),
    .Z(mem_ld_mask[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output134 (.I(net134),
    .Z(mem_st_dat[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output135 (.I(net135),
    .Z(mem_st_dat[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output136 (.I(net136),
    .Z(mem_st_dat[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output137 (.I(net137),
    .Z(mem_st_dat[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output138 (.I(net138),
    .Z(mem_st_dat[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output139 (.I(net139),
    .Z(mem_st_dat[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output140 (.I(net140),
    .Z(mem_st_dat[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output141 (.I(net141),
    .Z(mem_st_dat[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output142 (.I(net142),
    .Z(mem_st_dat[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output143 (.I(net143),
    .Z(mem_st_dat[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output144 (.I(net144),
    .Z(mem_st_dat[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output145 (.I(net145),
    .Z(mem_st_dat[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output146 (.I(net146),
    .Z(mem_st_dat[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output147 (.I(net147),
    .Z(mem_st_dat[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output148 (.I(net148),
    .Z(mem_st_dat[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output149 (.I(net149),
    .Z(mem_st_dat[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output150 (.I(net150),
    .Z(mem_st_dat[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output151 (.I(net151),
    .Z(mem_st_dat[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output152 (.I(net152),
    .Z(mem_st_dat[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output153 (.I(net153),
    .Z(mem_st_dat[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output154 (.I(net154),
    .Z(mem_st_dat[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output155 (.I(net155),
    .Z(mem_st_dat[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output156 (.I(net156),
    .Z(mem_st_dat[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output157 (.I(net157),
    .Z(mem_st_dat[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output158 (.I(net158),
    .Z(mem_st_dat[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output159 (.I(net159),
    .Z(mem_st_dat[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output160 (.I(net160),
    .Z(mem_st_dat[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output161 (.I(net161),
    .Z(mem_st_dat[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output162 (.I(net162),
    .Z(mem_st_dat[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output163 (.I(net163),
    .Z(mem_st_dat[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output164 (.I(net164),
    .Z(mem_st_dat[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output165 (.I(net165),
    .Z(mem_st_dat[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output166 (.I(net166),
    .Z(mem_st_en));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output167 (.I(net167),
    .Z(mem_st_mask[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output168 (.I(net168),
    .Z(mem_st_mask[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output169 (.I(net169),
    .Z(mem_st_mask[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output170 (.I(net170),
    .Z(mem_st_mask[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output171 (.I(net171),
    .Z(pc_next[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output172 (.I(net172),
    .Z(pc_next[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output173 (.I(net173),
    .Z(pc_next[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output174 (.I(net174),
    .Z(pc_next[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output175 (.I(net175),
    .Z(pc_next[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output176 (.I(net176),
    .Z(pc_next[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output177 (.I(net177),
    .Z(pc_next[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output178 (.I(net178),
    .Z(pc_next[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output179 (.I(net179),
    .Z(pc_next[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output180 (.I(net180),
    .Z(pc_next[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output181 (.I(net181),
    .Z(pc_next[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output182 (.I(net182),
    .Z(pc_next[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output183 (.I(net183),
    .Z(pc_next[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output184 (.I(net184),
    .Z(pc_next[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output185 (.I(net185),
    .Z(pc_next[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output186 (.I(net186),
    .Z(pc_next[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output187 (.I(net187),
    .Z(pc_next[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output188 (.I(net188),
    .Z(pc_next[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output189 (.I(net189),
    .Z(pc_next[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output190 (.I(net190),
    .Z(pc_next[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output191 (.I(net191),
    .Z(pc_next[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output192 (.I(net192),
    .Z(pc_next[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output193 (.I(net193),
    .Z(pc_next[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output194 (.I(net194),
    .Z(pc_next[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output195 (.I(net195),
    .Z(pc_next[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output196 (.I(net196),
    .Z(pc_next[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output197 (.I(net197),
    .Z(pc_next[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output198 (.I(net198),
    .Z(pc_next[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output199 (.I(net199),
    .Z(pc_next[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output200 (.I(net200),
    .Z(pc_next[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output201 (.I(net201),
    .Z(pc_next[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output202 (.I(net202),
    .Z(pc_next[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output97 (.I(net97),
    .Z(mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output98 (.I(net98),
    .Z(mem_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output99 (.I(net99),
    .Z(mem_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer1 (.I(_1509_),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer10 (.I(_1752_),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer11 (.I(_2934_),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer12 (.I(_0656_),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer13 (.I(_0675_),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer14 (.I(net232),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer15 (.I(_0522_),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer16 (.I(_1439_),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer17 (.I(_1493_),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer18 (.I(_0564_),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer19 (.I(_1618_),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer2 (.I(_1509_),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer20 (.I(_1506_),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer21 (.I(_1733_),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer22 (.I(_1631_),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer23 (.I(_0883_),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer24 (.I(net226),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer25 (.I(_1598_),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer26 (.I(_0498_),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer27 (.I(_0610_),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer28 (.I(_0511_),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer29 (.I(_2317_),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer3 (.I(net210),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer30 (.I(_1519_),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer31 (.I(_2886_),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer32 (.I(_0739_),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer33 (.I(_1496_),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer34 (.I(_1648_),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer35 (.I(net238),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer36 (.I(net239),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer4 (.I(_2400_),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(_2400_),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer6 (.I(_2400_),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer7 (.I(net209),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer8 (.I(net121),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer9 (.I(_1742_),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire203 (.I(_2088_),
    .Z(net203));
endmodule

