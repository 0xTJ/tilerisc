magic
tech gf180mcuD
magscale 1 10
timestamp 1699637960
<< metal1 >>
rect 1344 36874 78624 36908
rect 1344 36822 10874 36874
rect 10926 36822 10978 36874
rect 11030 36822 11082 36874
rect 11134 36822 30194 36874
rect 30246 36822 30298 36874
rect 30350 36822 30402 36874
rect 30454 36822 49514 36874
rect 49566 36822 49618 36874
rect 49670 36822 49722 36874
rect 49774 36822 68834 36874
rect 68886 36822 68938 36874
rect 68990 36822 69042 36874
rect 69094 36822 78624 36874
rect 1344 36788 78624 36822
rect 43934 36706 43986 36718
rect 43934 36642 43986 36654
rect 47630 36706 47682 36718
rect 47630 36642 47682 36654
rect 56030 36706 56082 36718
rect 71822 36706 71874 36718
rect 64082 36654 64094 36706
rect 64146 36654 64158 36706
rect 56030 36642 56082 36654
rect 71822 36642 71874 36654
rect 75070 36706 75122 36718
rect 75070 36642 75122 36654
rect 1934 36594 1986 36606
rect 1934 36530 1986 36542
rect 6526 36594 6578 36606
rect 6526 36530 6578 36542
rect 8878 36594 8930 36606
rect 8878 36530 8930 36542
rect 11454 36594 11506 36606
rect 11454 36530 11506 36542
rect 13918 36594 13970 36606
rect 13918 36530 13970 36542
rect 16382 36594 16434 36606
rect 16382 36530 16434 36542
rect 18846 36594 18898 36606
rect 18846 36530 18898 36542
rect 19630 36594 19682 36606
rect 19630 36530 19682 36542
rect 21310 36594 21362 36606
rect 21310 36530 21362 36542
rect 22094 36594 22146 36606
rect 22094 36530 22146 36542
rect 23662 36594 23714 36606
rect 23662 36530 23714 36542
rect 26350 36594 26402 36606
rect 26350 36530 26402 36542
rect 31166 36594 31218 36606
rect 31166 36530 31218 36542
rect 31614 36594 31666 36606
rect 31614 36530 31666 36542
rect 34862 36594 34914 36606
rect 34862 36530 34914 36542
rect 35534 36594 35586 36606
rect 35534 36530 35586 36542
rect 38446 36594 38498 36606
rect 41010 36542 41022 36594
rect 41074 36542 41086 36594
rect 38446 36530 38498 36542
rect 6750 36482 6802 36494
rect 3938 36430 3950 36482
rect 4002 36430 4014 36482
rect 6750 36418 6802 36430
rect 9326 36482 9378 36494
rect 9326 36418 9378 36430
rect 11678 36482 11730 36494
rect 11678 36418 11730 36430
rect 14142 36482 14194 36494
rect 19070 36482 19122 36494
rect 17042 36430 17054 36482
rect 17106 36430 17118 36482
rect 14142 36418 14194 36430
rect 19070 36418 19122 36430
rect 21534 36482 21586 36494
rect 21534 36418 21586 36430
rect 24558 36482 24610 36494
rect 24558 36418 24610 36430
rect 25118 36482 25170 36494
rect 25118 36418 25170 36430
rect 27358 36482 27410 36494
rect 32846 36482 32898 36494
rect 29138 36430 29150 36482
rect 29202 36430 29214 36482
rect 30706 36430 30718 36482
rect 30770 36430 30782 36482
rect 27358 36418 27410 36430
rect 32846 36418 32898 36430
rect 33854 36482 33906 36494
rect 33854 36418 33906 36430
rect 34414 36482 34466 36494
rect 38670 36482 38722 36494
rect 36530 36430 36542 36482
rect 36594 36430 36606 36482
rect 34414 36418 34466 36430
rect 38670 36418 38722 36430
rect 39230 36482 39282 36494
rect 43026 36430 43038 36482
rect 43090 36430 43102 36482
rect 46274 36430 46286 36482
rect 46338 36430 46350 36482
rect 49858 36430 49870 36482
rect 49922 36430 49934 36482
rect 53666 36430 53678 36482
rect 53730 36430 53742 36482
rect 55010 36430 55022 36482
rect 55074 36430 55086 36482
rect 58930 36430 58942 36482
rect 58994 36430 59006 36482
rect 62626 36430 62638 36482
rect 62690 36430 62702 36482
rect 66546 36430 66558 36482
rect 66610 36430 66622 36482
rect 70802 36430 70814 36482
rect 70866 36430 70878 36482
rect 74050 36430 74062 36482
rect 74114 36430 74126 36482
rect 39230 36418 39282 36430
rect 7310 36370 7362 36382
rect 7310 36306 7362 36318
rect 9886 36370 9938 36382
rect 9886 36306 9938 36318
rect 12238 36370 12290 36382
rect 24110 36370 24162 36382
rect 14466 36318 14478 36370
rect 14530 36318 14542 36370
rect 12238 36306 12290 36318
rect 24110 36306 24162 36318
rect 27022 36370 27074 36382
rect 27022 36306 27074 36318
rect 29822 36370 29874 36382
rect 29822 36306 29874 36318
rect 30382 36370 30434 36382
rect 30382 36306 30434 36318
rect 32510 36370 32562 36382
rect 52098 36318 52110 36370
rect 52162 36318 52174 36370
rect 60610 36318 60622 36370
rect 60674 36318 60686 36370
rect 32510 36306 32562 36318
rect 17726 36258 17778 36270
rect 17266 36206 17278 36258
rect 17330 36206 17342 36258
rect 17726 36194 17778 36206
rect 25902 36258 25954 36270
rect 27694 36258 27746 36270
rect 26674 36206 26686 36258
rect 26738 36206 26750 36258
rect 25902 36194 25954 36206
rect 27694 36194 27746 36206
rect 28702 36258 28754 36270
rect 30494 36258 30546 36270
rect 28914 36206 28926 36258
rect 28978 36206 28990 36258
rect 28702 36194 28754 36206
rect 30494 36194 30546 36206
rect 32174 36258 32226 36270
rect 40014 36258 40066 36270
rect 33170 36206 33182 36258
rect 33234 36206 33246 36258
rect 36306 36206 36318 36258
rect 36370 36206 36382 36258
rect 32174 36194 32226 36206
rect 40014 36194 40066 36206
rect 46846 36258 46898 36270
rect 46846 36194 46898 36206
rect 50430 36258 50482 36270
rect 50430 36194 50482 36206
rect 65886 36258 65938 36270
rect 65886 36194 65938 36206
rect 67454 36258 67506 36270
rect 67454 36194 67506 36206
rect 70478 36258 70530 36270
rect 70478 36194 70530 36206
rect 1344 36090 78784 36124
rect 1344 36038 20534 36090
rect 20586 36038 20638 36090
rect 20690 36038 20742 36090
rect 20794 36038 39854 36090
rect 39906 36038 39958 36090
rect 40010 36038 40062 36090
rect 40114 36038 59174 36090
rect 59226 36038 59278 36090
rect 59330 36038 59382 36090
rect 59434 36038 78494 36090
rect 78546 36038 78598 36090
rect 78650 36038 78702 36090
rect 78754 36038 78784 36090
rect 1344 36004 78784 36038
rect 3278 35922 3330 35934
rect 3278 35858 3330 35870
rect 4622 35922 4674 35934
rect 4622 35858 4674 35870
rect 24782 35922 24834 35934
rect 30382 35922 30434 35934
rect 28242 35870 28254 35922
rect 28306 35870 28318 35922
rect 24782 35858 24834 35870
rect 30382 35858 30434 35870
rect 65438 35922 65490 35934
rect 65438 35858 65490 35870
rect 76638 35922 76690 35934
rect 76638 35858 76690 35870
rect 17726 35810 17778 35822
rect 38222 35810 38274 35822
rect 28802 35758 28814 35810
rect 28866 35758 28878 35810
rect 37202 35758 37214 35810
rect 37266 35758 37278 35810
rect 17726 35746 17778 35758
rect 38222 35746 38274 35758
rect 48190 35810 48242 35822
rect 48190 35746 48242 35758
rect 48974 35810 49026 35822
rect 48974 35746 49026 35758
rect 50654 35810 50706 35822
rect 50654 35746 50706 35758
rect 54574 35810 54626 35822
rect 54574 35746 54626 35758
rect 63870 35810 63922 35822
rect 63870 35746 63922 35758
rect 67342 35810 67394 35822
rect 67342 35746 67394 35758
rect 71262 35810 71314 35822
rect 71262 35746 71314 35758
rect 17614 35698 17666 35710
rect 29038 35698 29090 35710
rect 4274 35646 4286 35698
rect 4338 35646 4350 35698
rect 10322 35646 10334 35698
rect 10386 35646 10398 35698
rect 13794 35646 13806 35698
rect 13858 35646 13870 35698
rect 19282 35646 19294 35698
rect 19346 35646 19358 35698
rect 25330 35646 25342 35698
rect 25394 35646 25406 35698
rect 17614 35634 17666 35646
rect 29038 35634 29090 35646
rect 29486 35698 29538 35710
rect 32398 35698 32450 35710
rect 30146 35646 30158 35698
rect 30210 35646 30222 35698
rect 31266 35646 31278 35698
rect 31330 35646 31342 35698
rect 29486 35634 29538 35646
rect 32398 35634 32450 35646
rect 33294 35698 33346 35710
rect 47630 35698 47682 35710
rect 36866 35646 36878 35698
rect 36930 35646 36942 35698
rect 38770 35646 38782 35698
rect 38834 35646 38846 35698
rect 45042 35646 45054 35698
rect 45106 35646 45118 35698
rect 46274 35646 46286 35698
rect 46338 35646 46350 35698
rect 33294 35634 33346 35646
rect 47630 35634 47682 35646
rect 47966 35698 48018 35710
rect 47966 35634 48018 35646
rect 48862 35698 48914 35710
rect 48862 35634 48914 35646
rect 49086 35698 49138 35710
rect 49086 35634 49138 35646
rect 50430 35698 50482 35710
rect 50430 35634 50482 35646
rect 50990 35698 51042 35710
rect 54910 35698 54962 35710
rect 67678 35698 67730 35710
rect 71598 35698 71650 35710
rect 51314 35646 51326 35698
rect 51378 35646 51390 35698
rect 60946 35646 60958 35698
rect 61010 35646 61022 35698
rect 64418 35646 64430 35698
rect 64482 35646 64494 35698
rect 68338 35646 68350 35698
rect 68402 35646 68414 35698
rect 73154 35646 73166 35698
rect 73218 35646 73230 35698
rect 76066 35646 76078 35698
rect 76130 35646 76142 35698
rect 50990 35634 51042 35646
rect 54910 35634 54962 35646
rect 67678 35634 67730 35646
rect 71598 35634 71650 35646
rect 5182 35586 5234 35598
rect 16606 35586 16658 35598
rect 10994 35534 11006 35586
rect 11058 35534 11070 35586
rect 13234 35534 13246 35586
rect 13298 35534 13310 35586
rect 14466 35534 14478 35586
rect 14530 35534 14542 35586
rect 5182 35522 5234 35534
rect 16606 35522 16658 35534
rect 18286 35586 18338 35598
rect 18286 35522 18338 35534
rect 19070 35586 19122 35598
rect 23662 35586 23714 35598
rect 28702 35586 28754 35598
rect 20066 35534 20078 35586
rect 20130 35534 20142 35586
rect 22306 35534 22318 35586
rect 22370 35534 22382 35586
rect 26002 35534 26014 35586
rect 26066 35534 26078 35586
rect 19070 35522 19122 35534
rect 23662 35522 23714 35534
rect 28702 35522 28754 35534
rect 30830 35586 30882 35598
rect 33070 35586 33122 35598
rect 31938 35534 31950 35586
rect 32002 35534 32014 35586
rect 30830 35522 30882 35534
rect 33070 35522 33122 35534
rect 35422 35586 35474 35598
rect 37774 35586 37826 35598
rect 39902 35586 39954 35598
rect 36530 35534 36542 35586
rect 36594 35534 36606 35586
rect 39106 35534 39118 35586
rect 39170 35534 39182 35586
rect 35422 35522 35474 35534
rect 37774 35522 37826 35534
rect 39902 35522 39954 35534
rect 42142 35586 42194 35598
rect 46958 35586 47010 35598
rect 44258 35534 44270 35586
rect 44322 35534 44334 35586
rect 45602 35534 45614 35586
rect 45666 35534 45678 35586
rect 42142 35522 42194 35534
rect 46958 35522 47010 35534
rect 47742 35586 47794 35598
rect 55358 35586 55410 35598
rect 69358 35586 69410 35598
rect 52098 35534 52110 35586
rect 52162 35534 52174 35586
rect 54226 35534 54238 35586
rect 54290 35534 54302 35586
rect 58034 35534 58046 35586
rect 58098 35534 58110 35586
rect 60274 35534 60286 35586
rect 60338 35534 60350 35586
rect 47742 35522 47794 35534
rect 55358 35522 55410 35534
rect 69358 35522 69410 35534
rect 72494 35586 72546 35598
rect 72494 35522 72546 35534
rect 75070 35586 75122 35598
rect 75070 35522 75122 35534
rect 17726 35474 17778 35486
rect 17726 35410 17778 35422
rect 29710 35474 29762 35486
rect 29710 35410 29762 35422
rect 30494 35474 30546 35486
rect 30494 35410 30546 35422
rect 33518 35474 33570 35486
rect 33518 35410 33570 35422
rect 33966 35474 34018 35486
rect 33966 35410 34018 35422
rect 37886 35474 37938 35486
rect 37886 35410 37938 35422
rect 40014 35474 40066 35486
rect 45490 35422 45502 35474
rect 45554 35422 45566 35474
rect 49522 35422 49534 35474
rect 49586 35422 49598 35474
rect 40014 35410 40066 35422
rect 1344 35306 78624 35340
rect 1344 35254 10874 35306
rect 10926 35254 10978 35306
rect 11030 35254 11082 35306
rect 11134 35254 30194 35306
rect 30246 35254 30298 35306
rect 30350 35254 30402 35306
rect 30454 35254 49514 35306
rect 49566 35254 49618 35306
rect 49670 35254 49722 35306
rect 49774 35254 68834 35306
rect 68886 35254 68938 35306
rect 68990 35254 69042 35306
rect 69094 35254 78624 35306
rect 1344 35220 78624 35254
rect 2942 35138 2994 35150
rect 2942 35074 2994 35086
rect 25454 35138 25506 35150
rect 44382 35138 44434 35150
rect 40562 35086 40574 35138
rect 40626 35086 40638 35138
rect 25454 35074 25506 35086
rect 44382 35074 44434 35086
rect 3502 35026 3554 35038
rect 3502 34962 3554 34974
rect 4398 35026 4450 35038
rect 4398 34962 4450 34974
rect 13582 35026 13634 35038
rect 13582 34962 13634 34974
rect 14254 35026 14306 35038
rect 14254 34962 14306 34974
rect 14702 35026 14754 35038
rect 18398 35026 18450 35038
rect 17714 34974 17726 35026
rect 17778 34974 17790 35026
rect 14702 34962 14754 34974
rect 18398 34962 18450 34974
rect 18958 35026 19010 35038
rect 43038 35026 43090 35038
rect 33506 34974 33518 35026
rect 33570 34974 33582 35026
rect 18958 34962 19010 34974
rect 43038 34962 43090 34974
rect 44942 35026 44994 35038
rect 44942 34962 44994 34974
rect 45390 35026 45442 35038
rect 45390 34962 45442 34974
rect 46398 35026 46450 35038
rect 53902 35026 53954 35038
rect 68574 35026 68626 35038
rect 73726 35026 73778 35038
rect 52098 34974 52110 35026
rect 52162 34974 52174 35026
rect 57250 34974 57262 35026
rect 57314 34974 57326 35026
rect 67666 34974 67678 35026
rect 67730 34974 67742 35026
rect 73042 34974 73054 35026
rect 73106 34974 73118 35026
rect 46398 34962 46450 34974
rect 53902 34962 53954 34974
rect 68574 34962 68626 34974
rect 73726 34962 73778 34974
rect 1822 34914 1874 34926
rect 1822 34850 1874 34862
rect 2382 34914 2434 34926
rect 2382 34850 2434 34862
rect 15374 34914 15426 34926
rect 15374 34850 15426 34862
rect 16270 34914 16322 34926
rect 16270 34850 16322 34862
rect 16494 34914 16546 34926
rect 16494 34850 16546 34862
rect 17054 34914 17106 34926
rect 26798 34914 26850 34926
rect 29486 34914 29538 34926
rect 30830 34914 30882 34926
rect 18050 34862 18062 34914
rect 18114 34862 18126 34914
rect 21522 34862 21534 34914
rect 21586 34862 21598 34914
rect 26562 34862 26574 34914
rect 26626 34862 26638 34914
rect 28354 34862 28366 34914
rect 28418 34862 28430 34914
rect 30034 34862 30046 34914
rect 30098 34862 30110 34914
rect 17054 34850 17106 34862
rect 26798 34850 26850 34862
rect 29486 34850 29538 34862
rect 30830 34850 30882 34862
rect 31166 34914 31218 34926
rect 34526 34914 34578 34926
rect 35870 34914 35922 34926
rect 37326 34914 37378 34926
rect 40350 34914 40402 34926
rect 43710 34914 43762 34926
rect 32834 34862 32846 34914
rect 32898 34862 32910 34914
rect 33842 34862 33854 34914
rect 33906 34862 33918 34914
rect 34738 34862 34750 34914
rect 34802 34862 34814 34914
rect 36194 34862 36206 34914
rect 36258 34862 36270 34914
rect 37762 34862 37774 34914
rect 37826 34862 37838 34914
rect 38434 34862 38446 34914
rect 38498 34862 38510 34914
rect 39330 34862 39342 34914
rect 39394 34862 39406 34914
rect 40562 34862 40574 34914
rect 40626 34862 40638 34914
rect 31166 34850 31218 34862
rect 34526 34850 34578 34862
rect 35870 34850 35922 34862
rect 37326 34850 37378 34862
rect 40350 34850 40402 34862
rect 43710 34850 43762 34862
rect 45614 34914 45666 34926
rect 45938 34862 45950 34914
rect 46002 34862 46014 34914
rect 47618 34862 47630 34914
rect 47682 34862 47694 34914
rect 47954 34862 47966 34914
rect 48018 34862 48030 34914
rect 49186 34862 49198 34914
rect 49250 34862 49262 34914
rect 54338 34862 54350 34914
rect 54402 34862 54414 34914
rect 60610 34862 60622 34914
rect 60674 34862 60686 34914
rect 64754 34862 64766 34914
rect 64818 34862 64830 34914
rect 70130 34862 70142 34914
rect 70194 34862 70206 34914
rect 45614 34850 45666 34862
rect 3054 34802 3106 34814
rect 3054 34738 3106 34750
rect 15710 34802 15762 34814
rect 25342 34802 25394 34814
rect 22194 34750 22206 34802
rect 22258 34750 22270 34802
rect 15710 34738 15762 34750
rect 25342 34738 25394 34750
rect 25902 34802 25954 34814
rect 25902 34738 25954 34750
rect 27358 34802 27410 34814
rect 27358 34738 27410 34750
rect 27470 34802 27522 34814
rect 27470 34738 27522 34750
rect 29710 34802 29762 34814
rect 29710 34738 29762 34750
rect 34302 34802 34354 34814
rect 42590 34802 42642 34814
rect 38546 34750 38558 34802
rect 38610 34750 38622 34802
rect 34302 34738 34354 34750
rect 42590 34738 42642 34750
rect 43486 34802 43538 34814
rect 43486 34738 43538 34750
rect 44046 34802 44098 34814
rect 44046 34738 44098 34750
rect 44270 34802 44322 34814
rect 44270 34738 44322 34750
rect 45726 34802 45778 34814
rect 57598 34802 57650 34814
rect 46946 34750 46958 34802
rect 47010 34750 47022 34802
rect 49970 34750 49982 34802
rect 50034 34750 50046 34802
rect 55122 34750 55134 34802
rect 55186 34750 55198 34802
rect 45726 34738 45778 34750
rect 57598 34738 57650 34750
rect 57934 34802 57986 34814
rect 61282 34750 61294 34802
rect 61346 34750 61358 34802
rect 65538 34750 65550 34802
rect 65602 34750 65614 34802
rect 70914 34750 70926 34802
rect 70978 34750 70990 34802
rect 57934 34738 57986 34750
rect 4734 34690 4786 34702
rect 4734 34626 4786 34638
rect 15598 34690 15650 34702
rect 15598 34626 15650 34638
rect 15934 34690 15986 34702
rect 25006 34690 25058 34702
rect 24434 34638 24446 34690
rect 24498 34638 24510 34690
rect 15934 34626 15986 34638
rect 25006 34626 25058 34638
rect 27134 34690 27186 34702
rect 27134 34626 27186 34638
rect 28030 34690 28082 34702
rect 29598 34690 29650 34702
rect 28578 34638 28590 34690
rect 28642 34638 28654 34690
rect 28030 34626 28082 34638
rect 29598 34626 29650 34638
rect 35758 34690 35810 34702
rect 35758 34626 35810 34638
rect 36430 34690 36482 34702
rect 36430 34626 36482 34638
rect 36542 34690 36594 34702
rect 41134 34690 41186 34702
rect 39330 34638 39342 34690
rect 39394 34638 39406 34690
rect 36542 34626 36594 34638
rect 41134 34626 41186 34638
rect 54014 34690 54066 34702
rect 75406 34690 75458 34702
rect 63522 34638 63534 34690
rect 63586 34638 63598 34690
rect 54014 34626 54066 34638
rect 75406 34626 75458 34638
rect 76302 34690 76354 34702
rect 76302 34626 76354 34638
rect 1344 34522 78784 34556
rect 1344 34470 20534 34522
rect 20586 34470 20638 34522
rect 20690 34470 20742 34522
rect 20794 34470 39854 34522
rect 39906 34470 39958 34522
rect 40010 34470 40062 34522
rect 40114 34470 59174 34522
rect 59226 34470 59278 34522
rect 59330 34470 59382 34522
rect 59434 34470 78494 34522
rect 78546 34470 78598 34522
rect 78650 34470 78702 34522
rect 78754 34470 78784 34522
rect 1344 34436 78784 34470
rect 16942 34354 16994 34366
rect 13906 34302 13918 34354
rect 13970 34302 13982 34354
rect 16942 34290 16994 34302
rect 20414 34354 20466 34366
rect 20414 34290 20466 34302
rect 24222 34354 24274 34366
rect 24222 34290 24274 34302
rect 26350 34354 26402 34366
rect 26350 34290 26402 34302
rect 27134 34354 27186 34366
rect 27134 34290 27186 34302
rect 27694 34354 27746 34366
rect 33070 34354 33122 34366
rect 29362 34302 29374 34354
rect 29426 34302 29438 34354
rect 27694 34290 27746 34302
rect 33070 34290 33122 34302
rect 33294 34354 33346 34366
rect 33294 34290 33346 34302
rect 41246 34354 41298 34366
rect 41246 34290 41298 34302
rect 41918 34354 41970 34366
rect 41918 34290 41970 34302
rect 44158 34354 44210 34366
rect 55582 34354 55634 34366
rect 65326 34354 65378 34366
rect 48066 34302 48078 34354
rect 48130 34302 48142 34354
rect 58146 34302 58158 34354
rect 58210 34302 58222 34354
rect 44158 34290 44210 34302
rect 55582 34290 55634 34302
rect 65326 34290 65378 34302
rect 24446 34242 24498 34254
rect 43486 34242 43538 34254
rect 28802 34190 28814 34242
rect 28866 34190 28878 34242
rect 24446 34178 24498 34190
rect 43486 34178 43538 34190
rect 44718 34242 44770 34254
rect 60062 34242 60114 34254
rect 70030 34242 70082 34254
rect 45826 34190 45838 34242
rect 45890 34190 45902 34242
rect 58818 34190 58830 34242
rect 58882 34190 58894 34242
rect 66434 34190 66446 34242
rect 66498 34190 66510 34242
rect 71026 34190 71038 34242
rect 71090 34190 71102 34242
rect 71362 34190 71374 34242
rect 71426 34190 71438 34242
rect 44718 34178 44770 34190
rect 60062 34178 60114 34190
rect 70030 34178 70082 34190
rect 20526 34130 20578 34142
rect 23886 34130 23938 34142
rect 4274 34078 4286 34130
rect 4338 34078 4350 34130
rect 10994 34078 11006 34130
rect 11058 34078 11070 34130
rect 14802 34078 14814 34130
rect 14866 34078 14878 34130
rect 15362 34078 15374 34130
rect 15426 34078 15438 34130
rect 17826 34078 17838 34130
rect 17890 34078 17902 34130
rect 18274 34078 18286 34130
rect 18338 34078 18350 34130
rect 22978 34078 22990 34130
rect 23042 34078 23054 34130
rect 23426 34078 23438 34130
rect 23490 34078 23502 34130
rect 20526 34066 20578 34078
rect 23886 34066 23938 34078
rect 24110 34130 24162 34142
rect 24110 34066 24162 34078
rect 25902 34130 25954 34142
rect 25902 34066 25954 34078
rect 26798 34130 26850 34142
rect 33182 34130 33234 34142
rect 28914 34078 28926 34130
rect 28978 34078 28990 34130
rect 29474 34078 29486 34130
rect 29538 34078 29550 34130
rect 29810 34078 29822 34130
rect 29874 34078 29886 34130
rect 32050 34078 32062 34130
rect 32114 34078 32126 34130
rect 26798 34066 26850 34078
rect 33182 34066 33234 34078
rect 33742 34130 33794 34142
rect 40798 34130 40850 34142
rect 33954 34078 33966 34130
rect 34018 34078 34030 34130
rect 34290 34078 34302 34130
rect 34354 34078 34366 34130
rect 36530 34078 36542 34130
rect 36594 34078 36606 34130
rect 36978 34078 36990 34130
rect 37042 34078 37054 34130
rect 40114 34078 40126 34130
rect 40178 34078 40190 34130
rect 33742 34066 33794 34078
rect 40798 34066 40850 34078
rect 41470 34130 41522 34142
rect 41470 34066 41522 34078
rect 41694 34130 41746 34142
rect 41694 34066 41746 34078
rect 42030 34130 42082 34142
rect 42030 34066 42082 34078
rect 44382 34130 44434 34142
rect 54126 34130 54178 34142
rect 60398 34130 60450 34142
rect 69694 34130 69746 34142
rect 45154 34078 45166 34130
rect 45218 34078 45230 34130
rect 49410 34078 49422 34130
rect 49474 34078 49486 34130
rect 53666 34078 53678 34130
rect 53730 34078 53742 34130
rect 54450 34078 54462 34130
rect 54514 34078 54526 34130
rect 57250 34078 57262 34130
rect 57314 34078 57326 34130
rect 58034 34078 58046 34130
rect 58098 34078 58110 34130
rect 59042 34078 59054 34130
rect 59106 34078 59118 34130
rect 60722 34078 60734 34130
rect 60786 34078 60798 34130
rect 65090 34078 65102 34130
rect 65154 34078 65166 34130
rect 65650 34078 65662 34130
rect 65714 34078 65726 34130
rect 44382 34066 44434 34078
rect 54126 34066 54178 34078
rect 60398 34066 60450 34078
rect 69694 34066 69746 34078
rect 70478 34130 70530 34142
rect 70478 34066 70530 34078
rect 70814 34130 70866 34142
rect 73154 34078 73166 34130
rect 73218 34078 73230 34130
rect 75618 34078 75630 34130
rect 75682 34078 75694 34130
rect 70814 34066 70866 34078
rect 4846 34018 4898 34030
rect 18510 34018 18562 34030
rect 11666 33966 11678 34018
rect 11730 33966 11742 34018
rect 15922 33966 15934 34018
rect 15986 33966 15998 34018
rect 4846 33954 4898 33966
rect 18510 33954 18562 33966
rect 19518 34018 19570 34030
rect 25342 34018 25394 34030
rect 21858 33966 21870 34018
rect 21922 33966 21934 34018
rect 19518 33954 19570 33966
rect 25342 33954 25394 33966
rect 27918 34018 27970 34030
rect 27918 33954 27970 33966
rect 28030 34018 28082 34030
rect 41358 34018 41410 34030
rect 29698 33966 29710 34018
rect 29762 34015 29774 34018
rect 29922 34015 29934 34018
rect 29762 33969 29934 34015
rect 29762 33966 29774 33969
rect 29922 33966 29934 33969
rect 29986 33966 29998 34018
rect 31938 33966 31950 34018
rect 32002 33966 32014 34018
rect 36082 33966 36094 34018
rect 36146 33966 36158 34018
rect 37426 33966 37438 34018
rect 37490 33966 37502 34018
rect 39666 33966 39678 34018
rect 39730 33966 39742 34018
rect 28030 33954 28082 33966
rect 41358 33954 41410 33966
rect 48750 34018 48802 34030
rect 51326 34018 51378 34030
rect 49186 33966 49198 34018
rect 49250 33966 49262 34018
rect 48750 33954 48802 33966
rect 51326 33954 51378 33966
rect 54014 34018 54066 34030
rect 54014 33954 54066 33966
rect 55358 34018 55410 34030
rect 55358 33954 55410 33966
rect 55470 34018 55522 34030
rect 63646 34018 63698 34030
rect 69358 34018 69410 34030
rect 57138 33966 57150 34018
rect 57202 33966 57214 34018
rect 61506 33966 61518 34018
rect 61570 33966 61582 34018
rect 68562 33966 68574 34018
rect 68626 33966 68638 34018
rect 73938 33966 73950 34018
rect 74002 33966 74014 34018
rect 55470 33954 55522 33966
rect 63646 33954 63698 33966
rect 69358 33954 69410 33966
rect 1934 33906 1986 33918
rect 38894 33906 38946 33918
rect 77982 33906 78034 33918
rect 32386 33854 32398 33906
rect 32450 33854 32462 33906
rect 56914 33854 56926 33906
rect 56978 33854 56990 33906
rect 1934 33842 1986 33854
rect 38894 33842 38946 33854
rect 77982 33842 78034 33854
rect 1344 33738 78624 33772
rect 1344 33686 10874 33738
rect 10926 33686 10978 33738
rect 11030 33686 11082 33738
rect 11134 33686 30194 33738
rect 30246 33686 30298 33738
rect 30350 33686 30402 33738
rect 30454 33686 49514 33738
rect 49566 33686 49618 33738
rect 49670 33686 49722 33738
rect 49774 33686 68834 33738
rect 68886 33686 68938 33738
rect 68990 33686 69042 33738
rect 69094 33686 78624 33738
rect 1344 33652 78624 33686
rect 12574 33570 12626 33582
rect 12574 33506 12626 33518
rect 15150 33570 15202 33582
rect 29262 33570 29314 33582
rect 15698 33518 15710 33570
rect 15762 33518 15774 33570
rect 15150 33506 15202 33518
rect 29262 33506 29314 33518
rect 31502 33570 31554 33582
rect 31502 33506 31554 33518
rect 35870 33570 35922 33582
rect 35870 33506 35922 33518
rect 37102 33570 37154 33582
rect 37102 33506 37154 33518
rect 48862 33570 48914 33582
rect 48862 33506 48914 33518
rect 56030 33570 56082 33582
rect 56030 33506 56082 33518
rect 57150 33570 57202 33582
rect 57150 33506 57202 33518
rect 61966 33570 62018 33582
rect 61966 33506 62018 33518
rect 66446 33570 66498 33582
rect 66446 33506 66498 33518
rect 3278 33458 3330 33470
rect 3278 33394 3330 33406
rect 13470 33458 13522 33470
rect 13470 33394 13522 33406
rect 19742 33458 19794 33470
rect 19742 33394 19794 33406
rect 21422 33458 21474 33470
rect 21422 33394 21474 33406
rect 23662 33458 23714 33470
rect 23662 33394 23714 33406
rect 24782 33458 24834 33470
rect 27246 33458 27298 33470
rect 25442 33406 25454 33458
rect 25506 33406 25518 33458
rect 24782 33394 24834 33406
rect 27246 33394 27298 33406
rect 31390 33458 31442 33470
rect 36206 33458 36258 33470
rect 43486 33458 43538 33470
rect 32386 33406 32398 33458
rect 32450 33406 32462 33458
rect 33954 33406 33966 33458
rect 34018 33406 34030 33458
rect 38322 33406 38334 33458
rect 38386 33406 38398 33458
rect 31390 33394 31442 33406
rect 36206 33394 36258 33406
rect 43486 33394 43538 33406
rect 44830 33458 44882 33470
rect 45378 33406 45390 33458
rect 45442 33406 45454 33458
rect 55346 33406 55358 33458
rect 55410 33406 55422 33458
rect 70802 33406 70814 33458
rect 70866 33406 70878 33458
rect 72930 33406 72942 33458
rect 72994 33406 73006 33458
rect 44830 33394 44882 33406
rect 14478 33346 14530 33358
rect 14478 33282 14530 33294
rect 14814 33346 14866 33358
rect 23550 33346 23602 33358
rect 26686 33346 26738 33358
rect 15138 33294 15150 33346
rect 15202 33294 15214 33346
rect 15698 33294 15710 33346
rect 15762 33294 15774 33346
rect 18946 33294 18958 33346
rect 19010 33294 19022 33346
rect 19282 33294 19294 33346
rect 19346 33294 19358 33346
rect 22082 33294 22094 33346
rect 22146 33294 22158 33346
rect 25330 33294 25342 33346
rect 25394 33294 25406 33346
rect 14814 33282 14866 33294
rect 23550 33282 23602 33294
rect 26686 33282 26738 33294
rect 28254 33346 28306 33358
rect 28254 33282 28306 33294
rect 29374 33346 29426 33358
rect 37214 33346 37266 33358
rect 45054 33346 45106 33358
rect 30370 33294 30382 33346
rect 30434 33294 30446 33346
rect 33842 33294 33854 33346
rect 33906 33294 33918 33346
rect 37762 33294 37774 33346
rect 37826 33294 37838 33346
rect 39442 33294 39454 33346
rect 39506 33294 39518 33346
rect 40786 33294 40798 33346
rect 40850 33294 40862 33346
rect 29374 33282 29426 33294
rect 37214 33282 37266 33294
rect 45054 33282 45106 33294
rect 45838 33346 45890 33358
rect 51662 33346 51714 33358
rect 49186 33294 49198 33346
rect 49250 33294 49262 33346
rect 45838 33282 45890 33294
rect 51662 33282 51714 33294
rect 51998 33346 52050 33358
rect 55806 33346 55858 33358
rect 58046 33346 58098 33358
rect 54898 33294 54910 33346
rect 54962 33294 54974 33346
rect 56354 33294 56366 33346
rect 56418 33294 56430 33346
rect 51998 33282 52050 33294
rect 55806 33282 55858 33294
rect 58046 33282 58098 33294
rect 58158 33346 58210 33358
rect 59054 33346 59106 33358
rect 66782 33346 66834 33358
rect 58370 33294 58382 33346
rect 58434 33294 58446 33346
rect 59266 33294 59278 33346
rect 59330 33294 59342 33346
rect 61058 33294 61070 33346
rect 61122 33294 61134 33346
rect 70018 33294 70030 33346
rect 70082 33294 70094 33346
rect 58158 33282 58210 33294
rect 59054 33282 59106 33294
rect 66782 33282 66834 33294
rect 12686 33234 12738 33246
rect 12686 33170 12738 33182
rect 13582 33234 13634 33246
rect 16270 33234 16322 33246
rect 16034 33182 16046 33234
rect 16098 33182 16110 33234
rect 13582 33170 13634 33182
rect 16270 33170 16322 33182
rect 18622 33234 18674 33246
rect 18622 33170 18674 33182
rect 18734 33234 18786 33246
rect 18734 33170 18786 33182
rect 20638 33234 20690 33246
rect 20638 33170 20690 33182
rect 20750 33234 20802 33246
rect 20750 33170 20802 33182
rect 21534 33234 21586 33246
rect 21534 33170 21586 33182
rect 21646 33234 21698 33246
rect 25566 33234 25618 33246
rect 25218 33182 25230 33234
rect 25282 33182 25294 33234
rect 21646 33170 21698 33182
rect 25566 33170 25618 33182
rect 29262 33234 29314 33246
rect 31166 33234 31218 33246
rect 30034 33182 30046 33234
rect 30098 33182 30110 33234
rect 29262 33170 29314 33182
rect 31166 33170 31218 33182
rect 31838 33234 31890 33246
rect 32286 33234 32338 33246
rect 32050 33182 32062 33234
rect 32114 33182 32126 33234
rect 31838 33170 31890 33182
rect 32286 33170 32338 33182
rect 32846 33234 32898 33246
rect 32846 33170 32898 33182
rect 36430 33234 36482 33246
rect 51774 33234 51826 33246
rect 37986 33182 37998 33234
rect 38050 33182 38062 33234
rect 43026 33182 43038 33234
rect 43090 33182 43102 33234
rect 36430 33170 36482 33182
rect 51774 33170 51826 33182
rect 54462 33234 54514 33246
rect 54462 33170 54514 33182
rect 57150 33234 57202 33246
rect 57150 33170 57202 33182
rect 57262 33234 57314 33246
rect 57262 33170 57314 33182
rect 59950 33234 60002 33246
rect 76302 33234 76354 33246
rect 66994 33182 67006 33234
rect 67058 33182 67070 33234
rect 67330 33182 67342 33234
rect 67394 33182 67406 33234
rect 59950 33170 60002 33182
rect 76302 33170 76354 33182
rect 14142 33122 14194 33134
rect 16718 33122 16770 33134
rect 15810 33070 15822 33122
rect 15874 33070 15886 33122
rect 14142 33058 14194 33070
rect 16718 33058 16770 33070
rect 18510 33122 18562 33134
rect 18510 33058 18562 33070
rect 20302 33122 20354 33134
rect 20302 33058 20354 33070
rect 20414 33122 20466 33134
rect 20414 33058 20466 33070
rect 21310 33122 21362 33134
rect 21310 33058 21362 33070
rect 22878 33122 22930 33134
rect 22878 33058 22930 33070
rect 23326 33122 23378 33134
rect 23326 33058 23378 33070
rect 23774 33122 23826 33134
rect 23774 33058 23826 33070
rect 24334 33122 24386 33134
rect 24334 33058 24386 33070
rect 25790 33122 25842 33134
rect 25790 33058 25842 33070
rect 26350 33122 26402 33134
rect 26350 33058 26402 33070
rect 28590 33122 28642 33134
rect 34750 33122 34802 33134
rect 29810 33070 29822 33122
rect 29874 33070 29886 33122
rect 28590 33058 28642 33070
rect 34750 33058 34802 33070
rect 37102 33122 37154 33134
rect 37102 33058 37154 33070
rect 42702 33122 42754 33134
rect 42702 33058 42754 33070
rect 43934 33122 43986 33134
rect 43934 33058 43986 33070
rect 46286 33122 46338 33134
rect 46286 33058 46338 33070
rect 48974 33122 49026 33134
rect 65998 33122 66050 33134
rect 57586 33070 57598 33122
rect 57650 33070 57662 33122
rect 48974 33058 49026 33070
rect 65998 33058 66050 33070
rect 75406 33122 75458 33134
rect 75406 33058 75458 33070
rect 1344 32954 78784 32988
rect 1344 32902 20534 32954
rect 20586 32902 20638 32954
rect 20690 32902 20742 32954
rect 20794 32902 39854 32954
rect 39906 32902 39958 32954
rect 40010 32902 40062 32954
rect 40114 32902 59174 32954
rect 59226 32902 59278 32954
rect 59330 32902 59382 32954
rect 59434 32902 78494 32954
rect 78546 32902 78598 32954
rect 78650 32902 78702 32954
rect 78754 32902 78784 32954
rect 1344 32868 78784 32902
rect 14254 32786 14306 32798
rect 14254 32722 14306 32734
rect 14366 32786 14418 32798
rect 14366 32722 14418 32734
rect 16382 32786 16434 32798
rect 16382 32722 16434 32734
rect 20974 32786 21026 32798
rect 20974 32722 21026 32734
rect 22990 32786 23042 32798
rect 22990 32722 23042 32734
rect 33294 32786 33346 32798
rect 33294 32722 33346 32734
rect 36990 32786 37042 32798
rect 36990 32722 37042 32734
rect 39006 32786 39058 32798
rect 45614 32786 45666 32798
rect 39330 32734 39342 32786
rect 39394 32734 39406 32786
rect 43026 32734 43038 32786
rect 43090 32734 43102 32786
rect 44258 32734 44270 32786
rect 44322 32734 44334 32786
rect 39006 32722 39058 32734
rect 45614 32722 45666 32734
rect 46286 32786 46338 32798
rect 46286 32722 46338 32734
rect 49870 32786 49922 32798
rect 49870 32722 49922 32734
rect 57374 32786 57426 32798
rect 57374 32722 57426 32734
rect 59838 32786 59890 32798
rect 59838 32722 59890 32734
rect 67790 32786 67842 32798
rect 67790 32722 67842 32734
rect 71598 32786 71650 32798
rect 71598 32722 71650 32734
rect 72382 32786 72434 32798
rect 72382 32722 72434 32734
rect 13918 32674 13970 32686
rect 13918 32610 13970 32622
rect 15374 32674 15426 32686
rect 15374 32610 15426 32622
rect 19518 32674 19570 32686
rect 19518 32610 19570 32622
rect 23662 32674 23714 32686
rect 23662 32610 23714 32622
rect 25230 32674 25282 32686
rect 38894 32674 38946 32686
rect 28242 32622 28254 32674
rect 28306 32622 28318 32674
rect 37202 32622 37214 32674
rect 37266 32622 37278 32674
rect 25230 32610 25282 32622
rect 38894 32610 38946 32622
rect 44830 32674 44882 32686
rect 44830 32610 44882 32622
rect 45166 32674 45218 32686
rect 50766 32674 50818 32686
rect 46610 32622 46622 32674
rect 46674 32622 46686 32674
rect 45166 32610 45218 32622
rect 50766 32610 50818 32622
rect 59950 32674 60002 32686
rect 66882 32622 66894 32674
rect 66946 32622 66958 32674
rect 70690 32622 70702 32674
rect 70754 32622 70766 32674
rect 59950 32610 60002 32622
rect 14142 32562 14194 32574
rect 15150 32562 15202 32574
rect 14578 32510 14590 32562
rect 14642 32510 14654 32562
rect 14914 32510 14926 32562
rect 14978 32510 14990 32562
rect 14142 32498 14194 32510
rect 15150 32498 15202 32510
rect 15486 32562 15538 32574
rect 15486 32498 15538 32510
rect 18958 32562 19010 32574
rect 19966 32562 20018 32574
rect 25790 32562 25842 32574
rect 19282 32510 19294 32562
rect 19346 32510 19358 32562
rect 25442 32510 25454 32562
rect 25506 32510 25518 32562
rect 18958 32498 19010 32510
rect 19966 32498 20018 32510
rect 25790 32498 25842 32510
rect 26126 32562 26178 32574
rect 26126 32498 26178 32510
rect 27358 32562 27410 32574
rect 30830 32562 30882 32574
rect 36654 32562 36706 32574
rect 28130 32510 28142 32562
rect 28194 32510 28206 32562
rect 29922 32510 29934 32562
rect 29986 32510 29998 32562
rect 31826 32510 31838 32562
rect 31890 32510 31902 32562
rect 27358 32498 27410 32510
rect 30830 32498 30882 32510
rect 36654 32498 36706 32510
rect 37438 32562 37490 32574
rect 37438 32498 37490 32510
rect 37886 32562 37938 32574
rect 37886 32498 37938 32510
rect 39678 32562 39730 32574
rect 39678 32498 39730 32510
rect 39902 32562 39954 32574
rect 39902 32498 39954 32510
rect 43374 32562 43426 32574
rect 43374 32498 43426 32510
rect 43710 32562 43762 32574
rect 43710 32498 43762 32510
rect 50654 32562 50706 32574
rect 50654 32498 50706 32510
rect 50990 32562 51042 32574
rect 67454 32562 67506 32574
rect 51538 32510 51550 32562
rect 51602 32510 51614 32562
rect 58146 32510 58158 32562
rect 58210 32510 58222 32562
rect 60722 32510 60734 32562
rect 60786 32510 60798 32562
rect 66658 32510 66670 32562
rect 66722 32510 66734 32562
rect 70466 32510 70478 32562
rect 70530 32510 70542 32562
rect 72706 32510 72718 32562
rect 72770 32510 72782 32562
rect 75618 32510 75630 32562
rect 75682 32510 75694 32562
rect 50990 32498 51042 32510
rect 67454 32498 67506 32510
rect 15934 32450 15986 32462
rect 15934 32386 15986 32398
rect 19182 32450 19234 32462
rect 19182 32386 19234 32398
rect 20414 32450 20466 32462
rect 20414 32386 20466 32398
rect 22542 32450 22594 32462
rect 26574 32450 26626 32462
rect 23650 32398 23662 32450
rect 23714 32398 23726 32450
rect 25330 32398 25342 32450
rect 25394 32398 25406 32450
rect 22542 32386 22594 32398
rect 26574 32386 26626 32398
rect 27918 32450 27970 32462
rect 27918 32386 27970 32398
rect 30718 32450 30770 32462
rect 30718 32386 30770 32398
rect 33854 32450 33906 32462
rect 33854 32386 33906 32398
rect 34302 32450 34354 32462
rect 34302 32386 34354 32398
rect 35758 32450 35810 32462
rect 35758 32386 35810 32398
rect 36318 32450 36370 32462
rect 38446 32450 38498 32462
rect 37538 32398 37550 32450
rect 37602 32398 37614 32450
rect 36318 32386 36370 32398
rect 38446 32386 38498 32398
rect 42030 32450 42082 32462
rect 42030 32386 42082 32398
rect 42702 32450 42754 32462
rect 42702 32386 42754 32398
rect 50430 32450 50482 32462
rect 63646 32450 63698 32462
rect 52322 32398 52334 32450
rect 52386 32398 52398 32450
rect 54450 32398 54462 32450
rect 54514 32398 54526 32450
rect 58482 32398 58494 32450
rect 58546 32398 58558 32450
rect 59378 32398 59390 32450
rect 59442 32398 59454 32450
rect 61506 32398 61518 32450
rect 61570 32398 61582 32450
rect 50430 32386 50482 32398
rect 63646 32386 63698 32398
rect 66222 32450 66274 32462
rect 66222 32386 66274 32398
rect 69246 32450 69298 32462
rect 69246 32386 69298 32398
rect 69806 32450 69858 32462
rect 69806 32386 69858 32398
rect 75070 32450 75122 32462
rect 75070 32386 75122 32398
rect 23886 32338 23938 32350
rect 23886 32274 23938 32286
rect 36542 32338 36594 32350
rect 36542 32274 36594 32286
rect 43934 32338 43986 32350
rect 43934 32274 43986 32286
rect 59726 32338 59778 32350
rect 59726 32274 59778 32286
rect 71262 32338 71314 32350
rect 71262 32274 71314 32286
rect 77982 32338 78034 32350
rect 77982 32274 78034 32286
rect 1344 32170 78624 32204
rect 1344 32118 10874 32170
rect 10926 32118 10978 32170
rect 11030 32118 11082 32170
rect 11134 32118 30194 32170
rect 30246 32118 30298 32170
rect 30350 32118 30402 32170
rect 30454 32118 49514 32170
rect 49566 32118 49618 32170
rect 49670 32118 49722 32170
rect 49774 32118 68834 32170
rect 68886 32118 68938 32170
rect 68990 32118 69042 32170
rect 69094 32118 78624 32170
rect 1344 32084 78624 32118
rect 29822 32002 29874 32014
rect 29822 31938 29874 31950
rect 37102 32002 37154 32014
rect 37102 31938 37154 31950
rect 44830 32002 44882 32014
rect 44830 31938 44882 31950
rect 60958 32002 61010 32014
rect 60958 31938 61010 31950
rect 1934 31890 1986 31902
rect 1934 31826 1986 31838
rect 15262 31890 15314 31902
rect 23326 31890 23378 31902
rect 18386 31838 18398 31890
rect 18450 31838 18462 31890
rect 20402 31838 20414 31890
rect 20466 31838 20478 31890
rect 15262 31826 15314 31838
rect 23326 31826 23378 31838
rect 25454 31890 25506 31902
rect 25454 31826 25506 31838
rect 29486 31890 29538 31902
rect 29486 31826 29538 31838
rect 31390 31890 31442 31902
rect 37326 31890 37378 31902
rect 33170 31838 33182 31890
rect 33234 31838 33246 31890
rect 31390 31826 31442 31838
rect 37326 31826 37378 31838
rect 39230 31890 39282 31902
rect 39230 31826 39282 31838
rect 46174 31890 46226 31902
rect 46174 31826 46226 31838
rect 53454 31890 53506 31902
rect 53454 31826 53506 31838
rect 59726 31890 59778 31902
rect 61618 31838 61630 31890
rect 61682 31838 61694 31890
rect 73378 31838 73390 31890
rect 73442 31838 73454 31890
rect 59726 31826 59778 31838
rect 22766 31778 22818 31790
rect 4274 31726 4286 31778
rect 4338 31726 4350 31778
rect 18834 31726 18846 31778
rect 18898 31726 18910 31778
rect 20290 31726 20302 31778
rect 20354 31726 20366 31778
rect 22418 31726 22430 31778
rect 22482 31726 22494 31778
rect 22766 31714 22818 31726
rect 23550 31778 23602 31790
rect 23550 31714 23602 31726
rect 24222 31778 24274 31790
rect 24222 31714 24274 31726
rect 24670 31778 24722 31790
rect 24670 31714 24722 31726
rect 26238 31778 26290 31790
rect 26238 31714 26290 31726
rect 26462 31778 26514 31790
rect 26462 31714 26514 31726
rect 26686 31778 26738 31790
rect 26686 31714 26738 31726
rect 30158 31778 30210 31790
rect 30158 31714 30210 31726
rect 31278 31778 31330 31790
rect 31278 31714 31330 31726
rect 31502 31778 31554 31790
rect 31502 31714 31554 31726
rect 31838 31778 31890 31790
rect 31838 31714 31890 31726
rect 32174 31778 32226 31790
rect 42590 31778 42642 31790
rect 32386 31726 32398 31778
rect 32450 31726 32462 31778
rect 33506 31726 33518 31778
rect 33570 31726 33582 31778
rect 37538 31726 37550 31778
rect 37602 31726 37614 31778
rect 38322 31726 38334 31778
rect 38386 31726 38398 31778
rect 38994 31726 39006 31778
rect 39058 31726 39070 31778
rect 41234 31726 41246 31778
rect 41298 31726 41310 31778
rect 32174 31714 32226 31726
rect 42590 31714 42642 31726
rect 43150 31778 43202 31790
rect 43150 31714 43202 31726
rect 51662 31778 51714 31790
rect 51662 31714 51714 31726
rect 53566 31778 53618 31790
rect 53566 31714 53618 31726
rect 53902 31778 53954 31790
rect 70466 31726 70478 31778
rect 70530 31726 70542 31778
rect 75394 31726 75406 31778
rect 75458 31726 75470 31778
rect 53902 31714 53954 31726
rect 8990 31666 9042 31678
rect 8990 31602 9042 31614
rect 16158 31666 16210 31678
rect 16158 31602 16210 31614
rect 17838 31666 17890 31678
rect 17838 31602 17890 31614
rect 22878 31666 22930 31678
rect 22878 31602 22930 31614
rect 25006 31666 25058 31678
rect 30382 31666 30434 31678
rect 27346 31614 27358 31666
rect 27410 31614 27422 31666
rect 25006 31602 25058 31614
rect 30382 31602 30434 31614
rect 30942 31666 30994 31678
rect 30942 31602 30994 31614
rect 32062 31666 32114 31678
rect 32062 31602 32114 31614
rect 41022 31666 41074 31678
rect 41022 31602 41074 31614
rect 42254 31666 42306 31678
rect 42254 31602 42306 31614
rect 42366 31666 42418 31678
rect 42366 31602 42418 31614
rect 42926 31666 42978 31678
rect 42926 31602 42978 31614
rect 43486 31666 43538 31678
rect 43486 31602 43538 31614
rect 44942 31666 44994 31678
rect 44942 31602 44994 31614
rect 49646 31666 49698 31678
rect 49646 31602 49698 31614
rect 49870 31666 49922 31678
rect 49870 31602 49922 31614
rect 50206 31666 50258 31678
rect 50206 31602 50258 31614
rect 50654 31666 50706 31678
rect 50654 31602 50706 31614
rect 50766 31666 50818 31678
rect 50766 31602 50818 31614
rect 51438 31666 51490 31678
rect 51438 31602 51490 31614
rect 51998 31666 52050 31678
rect 51998 31602 52050 31614
rect 53342 31666 53394 31678
rect 53342 31602 53394 31614
rect 60622 31666 60674 31678
rect 60622 31602 60674 31614
rect 60846 31666 60898 31678
rect 60846 31602 60898 31614
rect 61294 31666 61346 31678
rect 61294 31602 61346 31614
rect 61518 31666 61570 31678
rect 61518 31602 61570 31614
rect 64878 31666 64930 31678
rect 64878 31602 64930 31614
rect 65214 31666 65266 31678
rect 65214 31602 65266 31614
rect 65886 31666 65938 31678
rect 65886 31602 65938 31614
rect 69134 31666 69186 31678
rect 69134 31602 69186 31614
rect 69806 31666 69858 31678
rect 71250 31614 71262 31666
rect 71314 31614 71326 31666
rect 69806 31602 69858 31614
rect 8654 31554 8706 31566
rect 8654 31490 8706 31502
rect 9438 31554 9490 31566
rect 9438 31490 9490 31502
rect 15934 31554 15986 31566
rect 15934 31490 15986 31502
rect 16046 31554 16098 31566
rect 27134 31554 27186 31566
rect 23874 31502 23886 31554
rect 23938 31502 23950 31554
rect 16046 31490 16098 31502
rect 27134 31490 27186 31502
rect 27694 31554 27746 31566
rect 27694 31490 27746 31502
rect 32846 31554 32898 31566
rect 32846 31490 32898 31502
rect 37438 31554 37490 31566
rect 37438 31490 37490 31502
rect 38110 31554 38162 31566
rect 38110 31490 38162 31502
rect 43150 31554 43202 31566
rect 43150 31490 43202 31502
rect 43934 31554 43986 31566
rect 43934 31490 43986 31502
rect 45390 31554 45442 31566
rect 45390 31490 45442 31502
rect 46734 31554 46786 31566
rect 46734 31490 46786 31502
rect 48638 31554 48690 31566
rect 49982 31554 50034 31566
rect 48962 31502 48974 31554
rect 49026 31502 49038 31554
rect 48638 31490 48690 31502
rect 49982 31490 50034 31502
rect 50990 31554 51042 31566
rect 50990 31490 51042 31502
rect 51886 31554 51938 31566
rect 51886 31490 51938 31502
rect 58718 31554 58770 31566
rect 58718 31490 58770 31502
rect 65550 31554 65602 31566
rect 65550 31490 65602 31502
rect 66334 31554 66386 31566
rect 66334 31490 66386 31502
rect 69470 31554 69522 31566
rect 69470 31490 69522 31502
rect 70142 31554 70194 31566
rect 70142 31490 70194 31502
rect 75630 31554 75682 31566
rect 75630 31490 75682 31502
rect 1344 31386 78784 31420
rect 1344 31334 20534 31386
rect 20586 31334 20638 31386
rect 20690 31334 20742 31386
rect 20794 31334 39854 31386
rect 39906 31334 39958 31386
rect 40010 31334 40062 31386
rect 40114 31334 59174 31386
rect 59226 31334 59278 31386
rect 59330 31334 59382 31386
rect 59434 31334 78494 31386
rect 78546 31334 78598 31386
rect 78650 31334 78702 31386
rect 78754 31334 78784 31386
rect 1344 31300 78784 31334
rect 17950 31218 18002 31230
rect 17950 31154 18002 31166
rect 18510 31218 18562 31230
rect 18510 31154 18562 31166
rect 20414 31218 20466 31230
rect 33406 31218 33458 31230
rect 31490 31166 31502 31218
rect 31554 31166 31566 31218
rect 20414 31154 20466 31166
rect 33406 31154 33458 31166
rect 35646 31218 35698 31230
rect 35646 31154 35698 31166
rect 36990 31218 37042 31230
rect 43710 31218 43762 31230
rect 40002 31166 40014 31218
rect 40066 31166 40078 31218
rect 40226 31166 40238 31218
rect 40290 31166 40302 31218
rect 36990 31154 37042 31166
rect 43710 31154 43762 31166
rect 49422 31218 49474 31230
rect 49422 31154 49474 31166
rect 49646 31218 49698 31230
rect 49646 31154 49698 31166
rect 51102 31218 51154 31230
rect 51102 31154 51154 31166
rect 60062 31218 60114 31230
rect 60062 31154 60114 31166
rect 71038 31218 71090 31230
rect 71038 31154 71090 31166
rect 9550 31106 9602 31118
rect 19630 31106 19682 31118
rect 16370 31054 16382 31106
rect 16434 31054 16446 31106
rect 9550 31042 9602 31054
rect 19630 31042 19682 31054
rect 19854 31106 19906 31118
rect 19854 31042 19906 31054
rect 20078 31106 20130 31118
rect 20078 31042 20130 31054
rect 20190 31106 20242 31118
rect 44606 31106 44658 31118
rect 22866 31054 22878 31106
rect 22930 31054 22942 31106
rect 24098 31054 24110 31106
rect 24162 31054 24174 31106
rect 30146 31054 30158 31106
rect 30210 31054 30222 31106
rect 30818 31054 30830 31106
rect 30882 31054 30894 31106
rect 36082 31054 36094 31106
rect 36146 31054 36158 31106
rect 39330 31054 39342 31106
rect 39394 31054 39406 31106
rect 20190 31042 20242 31054
rect 44606 31042 44658 31054
rect 48974 31106 49026 31118
rect 48974 31042 49026 31054
rect 49310 31106 49362 31118
rect 49310 31042 49362 31054
rect 51774 31106 51826 31118
rect 51774 31042 51826 31054
rect 51998 31106 52050 31118
rect 69806 31106 69858 31118
rect 65426 31054 65438 31106
rect 65490 31054 65502 31106
rect 51998 31042 52050 31054
rect 69806 31042 69858 31054
rect 74174 31106 74226 31118
rect 74174 31042 74226 31054
rect 74510 31106 74562 31118
rect 74510 31042 74562 31054
rect 14814 30994 14866 31006
rect 18398 30994 18450 31006
rect 19518 30994 19570 31006
rect 26238 30994 26290 31006
rect 9762 30942 9774 30994
rect 9826 30942 9838 30994
rect 14466 30942 14478 30994
rect 14530 30942 14542 30994
rect 15474 30942 15486 30994
rect 15538 30942 15550 30994
rect 15810 30942 15822 30994
rect 15874 30942 15886 30994
rect 18610 30942 18622 30994
rect 18674 30942 18686 30994
rect 21410 30942 21422 30994
rect 21474 30942 21486 30994
rect 24658 30942 24670 30994
rect 24722 30942 24734 30994
rect 25890 30942 25902 30994
rect 25954 30942 25966 30994
rect 14814 30930 14866 30942
rect 18398 30930 18450 30942
rect 19518 30930 19570 30942
rect 26238 30930 26290 30942
rect 28254 30994 28306 31006
rect 37998 30994 38050 31006
rect 28578 30942 28590 30994
rect 28642 30942 28654 30994
rect 29922 30942 29934 30994
rect 29986 30942 29998 30994
rect 30482 30942 30494 30994
rect 30546 30942 30558 30994
rect 31602 30942 31614 30994
rect 31666 30942 31678 30994
rect 35970 30942 35982 30994
rect 36034 30942 36046 30994
rect 37202 30942 37214 30994
rect 37266 30942 37278 30994
rect 37426 30942 37438 30994
rect 37490 30942 37502 30994
rect 37762 30942 37774 30994
rect 37826 30942 37838 30994
rect 28254 30930 28306 30942
rect 37998 30930 38050 30942
rect 38110 30994 38162 31006
rect 41022 30994 41074 31006
rect 39442 30942 39454 30994
rect 39506 30942 39518 30994
rect 39778 30942 39790 30994
rect 39842 30942 39854 30994
rect 38110 30930 38162 30942
rect 41022 30930 41074 30942
rect 42142 30994 42194 31006
rect 42142 30930 42194 30942
rect 43598 30994 43650 31006
rect 43598 30930 43650 30942
rect 43822 30994 43874 31006
rect 43822 30930 43874 30942
rect 44270 30994 44322 31006
rect 44270 30930 44322 30942
rect 47518 30994 47570 31006
rect 47518 30930 47570 30942
rect 50990 30994 51042 31006
rect 50990 30930 51042 30942
rect 51326 30994 51378 31006
rect 51326 30930 51378 30942
rect 51550 30994 51602 31006
rect 51550 30930 51602 30942
rect 52222 30994 52274 31006
rect 59390 30994 59442 31006
rect 57810 30942 57822 30994
rect 57874 30942 57886 30994
rect 59042 30942 59054 30994
rect 59106 30942 59118 30994
rect 52222 30930 52274 30942
rect 59390 30930 59442 30942
rect 59950 30994 60002 31006
rect 59950 30930 60002 30942
rect 60398 30994 60450 31006
rect 70142 30994 70194 31006
rect 64754 30942 64766 30994
rect 64818 30942 64830 30994
rect 60398 30930 60450 30942
rect 70142 30930 70194 30942
rect 71374 30994 71426 31006
rect 74834 30942 74846 30994
rect 74898 30942 74910 30994
rect 71374 30930 71426 30942
rect 14926 30882 14978 30894
rect 16830 30882 16882 30894
rect 20750 30882 20802 30894
rect 34638 30882 34690 30894
rect 41806 30882 41858 30894
rect 43150 30882 43202 30894
rect 50654 30882 50706 30894
rect 58606 30882 58658 30894
rect 16258 30830 16270 30882
rect 16322 30830 16334 30882
rect 18050 30830 18062 30882
rect 18114 30830 18126 30882
rect 23426 30830 23438 30882
rect 23490 30830 23502 30882
rect 25330 30830 25342 30882
rect 25394 30830 25406 30882
rect 36642 30830 36654 30882
rect 36706 30830 36718 30882
rect 36978 30830 36990 30882
rect 37042 30830 37054 30882
rect 42578 30830 42590 30882
rect 42642 30830 42654 30882
rect 47954 30830 47966 30882
rect 48018 30830 48030 30882
rect 57586 30830 57598 30882
rect 57650 30830 57662 30882
rect 14926 30818 14978 30830
rect 16830 30818 16882 30830
rect 20750 30818 20802 30830
rect 34638 30818 34690 30830
rect 41806 30818 41858 30830
rect 43150 30818 43202 30830
rect 50654 30818 50706 30830
rect 58606 30818 58658 30830
rect 59726 30882 59778 30894
rect 68126 30882 68178 30894
rect 67554 30830 67566 30882
rect 67618 30830 67630 30882
rect 59726 30818 59778 30830
rect 68126 30818 68178 30830
rect 72494 30882 72546 30894
rect 75618 30830 75630 30882
rect 75682 30830 75694 30882
rect 77746 30830 77758 30882
rect 77810 30830 77822 30882
rect 72494 30818 72546 30830
rect 17726 30770 17778 30782
rect 59502 30770 59554 30782
rect 38546 30718 38558 30770
rect 38610 30718 38622 30770
rect 44370 30718 44382 30770
rect 44434 30767 44446 30770
rect 44706 30767 44718 30770
rect 44434 30721 44718 30767
rect 44434 30718 44446 30721
rect 44706 30718 44718 30721
rect 44770 30718 44782 30770
rect 57362 30718 57374 30770
rect 57426 30718 57438 30770
rect 58258 30718 58270 30770
rect 58322 30767 58334 30770
rect 58482 30767 58494 30770
rect 58322 30721 58494 30767
rect 58322 30718 58334 30721
rect 58482 30718 58494 30721
rect 58546 30718 58558 30770
rect 17726 30706 17778 30718
rect 59502 30706 59554 30718
rect 1344 30602 78624 30636
rect 1344 30550 10874 30602
rect 10926 30550 10978 30602
rect 11030 30550 11082 30602
rect 11134 30550 30194 30602
rect 30246 30550 30298 30602
rect 30350 30550 30402 30602
rect 30454 30550 49514 30602
rect 49566 30550 49618 30602
rect 49670 30550 49722 30602
rect 49774 30550 68834 30602
rect 68886 30550 68938 30602
rect 68990 30550 69042 30602
rect 69094 30550 78624 30602
rect 1344 30516 78624 30550
rect 17950 30434 18002 30446
rect 36094 30434 36146 30446
rect 16482 30382 16494 30434
rect 16546 30382 16558 30434
rect 20066 30382 20078 30434
rect 20130 30382 20142 30434
rect 26002 30382 26014 30434
rect 26066 30382 26078 30434
rect 17950 30370 18002 30382
rect 36094 30370 36146 30382
rect 36430 30434 36482 30446
rect 36430 30370 36482 30382
rect 53790 30434 53842 30446
rect 53790 30370 53842 30382
rect 19070 30322 19122 30334
rect 34526 30322 34578 30334
rect 9202 30270 9214 30322
rect 9266 30270 9278 30322
rect 11330 30270 11342 30322
rect 11394 30270 11406 30322
rect 23314 30270 23326 30322
rect 23378 30270 23390 30322
rect 24882 30270 24894 30322
rect 24946 30270 24958 30322
rect 25778 30270 25790 30322
rect 25842 30270 25854 30322
rect 28354 30270 28366 30322
rect 28418 30270 28430 30322
rect 19070 30258 19122 30270
rect 34526 30258 34578 30270
rect 35870 30322 35922 30334
rect 35870 30258 35922 30270
rect 39454 30322 39506 30334
rect 43710 30322 43762 30334
rect 61294 30322 61346 30334
rect 73390 30322 73442 30334
rect 41906 30270 41918 30322
rect 41970 30270 41982 30322
rect 46834 30270 46846 30322
rect 46898 30270 46910 30322
rect 69794 30270 69806 30322
rect 69858 30270 69870 30322
rect 39454 30258 39506 30270
rect 43710 30258 43762 30270
rect 61294 30258 61346 30270
rect 73390 30258 73442 30270
rect 74734 30322 74786 30334
rect 74734 30258 74786 30270
rect 76638 30322 76690 30334
rect 76638 30258 76690 30270
rect 15598 30210 15650 30222
rect 17838 30210 17890 30222
rect 8530 30158 8542 30210
rect 8594 30158 8606 30210
rect 14354 30158 14366 30210
rect 14418 30158 14430 30210
rect 14690 30158 14702 30210
rect 14754 30158 14766 30210
rect 17266 30158 17278 30210
rect 17330 30158 17342 30210
rect 15598 30146 15650 30158
rect 17838 30146 17890 30158
rect 18622 30210 18674 30222
rect 31726 30210 31778 30222
rect 19506 30158 19518 30210
rect 19570 30158 19582 30210
rect 21746 30158 21758 30210
rect 21810 30158 21822 30210
rect 22082 30158 22094 30210
rect 22146 30158 22158 30210
rect 23762 30158 23774 30210
rect 23826 30158 23838 30210
rect 23986 30158 23998 30210
rect 24050 30158 24062 30210
rect 24770 30158 24782 30210
rect 24834 30158 24846 30210
rect 25666 30158 25678 30210
rect 25730 30158 25742 30210
rect 28242 30158 28254 30210
rect 28306 30158 28318 30210
rect 29586 30158 29598 30210
rect 29650 30158 29662 30210
rect 18622 30146 18674 30158
rect 31726 30146 31778 30158
rect 34078 30210 34130 30222
rect 34078 30146 34130 30158
rect 34302 30210 34354 30222
rect 34302 30146 34354 30158
rect 34862 30210 34914 30222
rect 39118 30210 39170 30222
rect 42590 30210 42642 30222
rect 37650 30158 37662 30210
rect 37714 30158 37726 30210
rect 38098 30158 38110 30210
rect 38162 30158 38174 30210
rect 38658 30158 38670 30210
rect 38722 30158 38734 30210
rect 41458 30158 41470 30210
rect 41522 30158 41534 30210
rect 34862 30146 34914 30158
rect 39118 30146 39170 30158
rect 42590 30146 42642 30158
rect 48078 30210 48130 30222
rect 48078 30146 48130 30158
rect 53566 30210 53618 30222
rect 53566 30146 53618 30158
rect 56702 30210 56754 30222
rect 60958 30210 61010 30222
rect 58146 30158 58158 30210
rect 58210 30158 58222 30210
rect 58930 30158 58942 30210
rect 58994 30158 59006 30210
rect 59490 30158 59502 30210
rect 59554 30158 59566 30210
rect 60498 30158 60510 30210
rect 60562 30158 60574 30210
rect 56702 30146 56754 30158
rect 60958 30146 61010 30158
rect 61182 30210 61234 30222
rect 73726 30210 73778 30222
rect 77982 30210 78034 30222
rect 64642 30158 64654 30210
rect 64706 30158 64718 30210
rect 68562 30158 68574 30210
rect 68626 30158 68638 30210
rect 69122 30158 69134 30210
rect 69186 30158 69198 30210
rect 72818 30158 72830 30210
rect 72882 30158 72894 30210
rect 75506 30158 75518 30210
rect 75570 30158 75582 30210
rect 61182 30146 61234 30158
rect 73726 30146 73778 30158
rect 77982 30146 78034 30158
rect 3726 30098 3778 30110
rect 15934 30098 15986 30110
rect 20526 30098 20578 30110
rect 43598 30098 43650 30110
rect 15250 30046 15262 30098
rect 15314 30046 15326 30098
rect 16370 30046 16382 30098
rect 16434 30046 16446 30098
rect 28354 30046 28366 30098
rect 28418 30046 28430 30098
rect 29698 30046 29710 30098
rect 29762 30046 29774 30098
rect 33282 30046 33294 30098
rect 33346 30046 33358 30098
rect 37314 30046 37326 30098
rect 37378 30046 37390 30098
rect 3726 30034 3778 30046
rect 15934 30034 15986 30046
rect 20526 30034 20578 30046
rect 43598 30034 43650 30046
rect 43822 30098 43874 30110
rect 43822 30034 43874 30046
rect 47406 30098 47458 30110
rect 61406 30098 61458 30110
rect 57810 30046 57822 30098
rect 57874 30046 57886 30098
rect 58818 30046 58830 30098
rect 58882 30046 58894 30098
rect 60722 30046 60734 30098
rect 60786 30046 60798 30098
rect 47406 30034 47458 30046
rect 61406 30034 61458 30046
rect 61742 30098 61794 30110
rect 76302 30098 76354 30110
rect 65314 30046 65326 30098
rect 65378 30046 65390 30098
rect 72706 30046 72718 30098
rect 72770 30046 72782 30098
rect 75282 30046 75294 30098
rect 75346 30046 75358 30098
rect 76962 30046 76974 30098
rect 77026 30046 77038 30098
rect 77410 30046 77422 30098
rect 77474 30046 77486 30098
rect 61742 30034 61794 30046
rect 76302 30034 76354 30046
rect 3390 29986 3442 29998
rect 3390 29922 3442 29934
rect 5854 29986 5906 29998
rect 5854 29922 5906 29934
rect 15822 29986 15874 29998
rect 15822 29922 15874 29934
rect 26686 29986 26738 29998
rect 26686 29922 26738 29934
rect 29262 29986 29314 29998
rect 29262 29922 29314 29934
rect 31166 29986 31218 29998
rect 31166 29922 31218 29934
rect 33854 29986 33906 29998
rect 33854 29922 33906 29934
rect 33966 29986 34018 29998
rect 43150 29986 43202 29998
rect 35186 29934 35198 29986
rect 35250 29934 35262 29986
rect 38098 29934 38110 29986
rect 38162 29934 38174 29986
rect 33966 29922 34018 29934
rect 43150 29922 43202 29934
rect 44046 29986 44098 29998
rect 44046 29922 44098 29934
rect 44942 29986 44994 29998
rect 45726 29986 45778 29998
rect 45266 29934 45278 29986
rect 45330 29934 45342 29986
rect 44942 29922 44994 29934
rect 45726 29922 45778 29934
rect 46846 29986 46898 29998
rect 46846 29922 46898 29934
rect 46958 29986 47010 29998
rect 46958 29922 47010 29934
rect 47182 29986 47234 29998
rect 57150 29986 57202 29998
rect 47730 29934 47742 29986
rect 47794 29934 47806 29986
rect 54114 29934 54126 29986
rect 54178 29934 54190 29986
rect 47182 29922 47234 29934
rect 57150 29922 57202 29934
rect 60062 29986 60114 29998
rect 74398 29986 74450 29998
rect 62066 29934 62078 29986
rect 62130 29934 62142 29986
rect 67554 29934 67566 29986
rect 67618 29934 67630 29986
rect 68338 29934 68350 29986
rect 68402 29934 68414 29986
rect 72034 29934 72046 29986
rect 72098 29934 72110 29986
rect 60062 29922 60114 29934
rect 74398 29922 74450 29934
rect 1344 29818 78784 29852
rect 1344 29766 20534 29818
rect 20586 29766 20638 29818
rect 20690 29766 20742 29818
rect 20794 29766 39854 29818
rect 39906 29766 39958 29818
rect 40010 29766 40062 29818
rect 40114 29766 59174 29818
rect 59226 29766 59278 29818
rect 59330 29766 59382 29818
rect 59434 29766 78494 29818
rect 78546 29766 78598 29818
rect 78650 29766 78702 29818
rect 78754 29766 78784 29818
rect 1344 29732 78784 29766
rect 5742 29650 5794 29662
rect 5742 29586 5794 29598
rect 9662 29650 9714 29662
rect 9662 29586 9714 29598
rect 16270 29650 16322 29662
rect 16270 29586 16322 29598
rect 17390 29650 17442 29662
rect 17390 29586 17442 29598
rect 17502 29650 17554 29662
rect 17502 29586 17554 29598
rect 19182 29650 19234 29662
rect 19182 29586 19234 29598
rect 20750 29650 20802 29662
rect 29934 29650 29986 29662
rect 22754 29598 22766 29650
rect 22818 29598 22830 29650
rect 20750 29586 20802 29598
rect 29934 29586 29986 29598
rect 30158 29650 30210 29662
rect 30158 29586 30210 29598
rect 32286 29650 32338 29662
rect 32286 29586 32338 29598
rect 35646 29650 35698 29662
rect 35646 29586 35698 29598
rect 38222 29650 38274 29662
rect 42030 29650 42082 29662
rect 38994 29598 39006 29650
rect 39058 29598 39070 29650
rect 40002 29598 40014 29650
rect 40066 29598 40078 29650
rect 38222 29586 38274 29598
rect 42030 29586 42082 29598
rect 42478 29650 42530 29662
rect 42478 29586 42530 29598
rect 43038 29650 43090 29662
rect 49086 29650 49138 29662
rect 47730 29598 47742 29650
rect 47794 29598 47806 29650
rect 43038 29586 43090 29598
rect 49086 29586 49138 29598
rect 49198 29650 49250 29662
rect 49198 29586 49250 29598
rect 51774 29650 51826 29662
rect 51774 29586 51826 29598
rect 51886 29650 51938 29662
rect 59726 29650 59778 29662
rect 53442 29598 53454 29650
rect 53506 29598 53518 29650
rect 54674 29598 54686 29650
rect 54738 29598 54750 29650
rect 51886 29586 51938 29598
rect 59726 29586 59778 29598
rect 60398 29650 60450 29662
rect 60398 29586 60450 29598
rect 62638 29650 62690 29662
rect 62638 29586 62690 29598
rect 65102 29650 65154 29662
rect 65102 29586 65154 29598
rect 65438 29650 65490 29662
rect 65438 29586 65490 29598
rect 70142 29650 70194 29662
rect 70142 29586 70194 29598
rect 74510 29650 74562 29662
rect 74510 29586 74562 29598
rect 7982 29538 8034 29550
rect 13134 29538 13186 29550
rect 3154 29486 3166 29538
rect 3218 29486 3230 29538
rect 6738 29486 6750 29538
rect 6802 29486 6814 29538
rect 10210 29486 10222 29538
rect 10274 29486 10286 29538
rect 10546 29486 10558 29538
rect 10610 29486 10622 29538
rect 7982 29474 8034 29486
rect 13134 29474 13186 29486
rect 13246 29538 13298 29550
rect 17838 29538 17890 29550
rect 15138 29486 15150 29538
rect 15202 29486 15214 29538
rect 13246 29474 13298 29486
rect 17838 29474 17890 29486
rect 20302 29538 20354 29550
rect 20302 29474 20354 29486
rect 20414 29538 20466 29550
rect 20414 29474 20466 29486
rect 20638 29538 20690 29550
rect 20638 29474 20690 29486
rect 20974 29538 21026 29550
rect 26126 29538 26178 29550
rect 32062 29538 32114 29550
rect 35534 29538 35586 29550
rect 38446 29538 38498 29550
rect 49646 29538 49698 29550
rect 22082 29486 22094 29538
rect 22146 29486 22158 29538
rect 24210 29486 24222 29538
rect 24274 29486 24286 29538
rect 26450 29486 26462 29538
rect 26514 29486 26526 29538
rect 27122 29486 27134 29538
rect 27186 29486 27198 29538
rect 33170 29486 33182 29538
rect 33234 29486 33246 29538
rect 35410 29486 35422 29538
rect 35474 29486 35486 29538
rect 36418 29486 36430 29538
rect 36482 29486 36494 29538
rect 40226 29486 40238 29538
rect 40290 29486 40302 29538
rect 43922 29486 43934 29538
rect 43986 29486 43998 29538
rect 46162 29486 46174 29538
rect 46226 29486 46238 29538
rect 47842 29486 47854 29538
rect 47906 29486 47918 29538
rect 20974 29474 21026 29486
rect 26126 29474 26178 29486
rect 32062 29474 32114 29486
rect 35534 29474 35586 29486
rect 38446 29474 38498 29486
rect 49646 29474 49698 29486
rect 49758 29538 49810 29550
rect 64766 29538 64818 29550
rect 55346 29486 55358 29538
rect 55410 29486 55422 29538
rect 60834 29486 60846 29538
rect 60898 29486 60910 29538
rect 66882 29486 66894 29538
rect 66946 29486 66958 29538
rect 67218 29486 67230 29538
rect 67282 29486 67294 29538
rect 70690 29486 70702 29538
rect 70754 29486 70766 29538
rect 71026 29486 71038 29538
rect 71090 29486 71102 29538
rect 72258 29486 72270 29538
rect 72322 29486 72334 29538
rect 75618 29486 75630 29538
rect 75682 29486 75694 29538
rect 49758 29474 49810 29486
rect 64766 29474 64818 29486
rect 8318 29426 8370 29438
rect 2482 29374 2494 29426
rect 2546 29374 2558 29426
rect 6514 29374 6526 29426
rect 6578 29374 6590 29426
rect 8318 29362 8370 29374
rect 9998 29426 10050 29438
rect 9998 29362 10050 29374
rect 13694 29426 13746 29438
rect 13694 29362 13746 29374
rect 14254 29426 14306 29438
rect 17614 29426 17666 29438
rect 19294 29426 19346 29438
rect 14914 29374 14926 29426
rect 14978 29374 14990 29426
rect 15586 29374 15598 29426
rect 15650 29374 15662 29426
rect 16482 29374 16494 29426
rect 16546 29374 16558 29426
rect 16706 29374 16718 29426
rect 16770 29374 16782 29426
rect 19058 29374 19070 29426
rect 19122 29374 19134 29426
rect 14254 29362 14306 29374
rect 17614 29362 17666 29374
rect 19294 29362 19346 29374
rect 21086 29426 21138 29438
rect 25566 29426 25618 29438
rect 29598 29426 29650 29438
rect 35870 29426 35922 29438
rect 22418 29374 22430 29426
rect 22482 29374 22494 29426
rect 23426 29374 23438 29426
rect 23490 29374 23502 29426
rect 26562 29374 26574 29426
rect 26626 29374 26638 29426
rect 27570 29374 27582 29426
rect 27634 29374 27646 29426
rect 30818 29374 30830 29426
rect 30882 29374 30894 29426
rect 31042 29374 31054 29426
rect 31106 29374 31118 29426
rect 33058 29374 33070 29426
rect 33122 29374 33134 29426
rect 33954 29374 33966 29426
rect 34018 29374 34030 29426
rect 21086 29362 21138 29374
rect 25566 29362 25618 29374
rect 29598 29362 29650 29374
rect 35870 29362 35922 29374
rect 36206 29426 36258 29438
rect 38558 29426 38610 29438
rect 42366 29426 42418 29438
rect 36866 29374 36878 29426
rect 36930 29374 36942 29426
rect 37650 29374 37662 29426
rect 37714 29374 37726 29426
rect 38882 29374 38894 29426
rect 38946 29374 38958 29426
rect 40114 29374 40126 29426
rect 40178 29374 40190 29426
rect 36206 29362 36258 29374
rect 38558 29362 38610 29374
rect 42366 29362 42418 29374
rect 42702 29426 42754 29438
rect 42702 29362 42754 29374
rect 43374 29426 43426 29438
rect 44718 29426 44770 29438
rect 44146 29374 44158 29426
rect 44210 29374 44222 29426
rect 43374 29362 43426 29374
rect 44718 29362 44770 29374
rect 48638 29426 48690 29438
rect 48638 29362 48690 29374
rect 49310 29426 49362 29438
rect 49310 29362 49362 29374
rect 51662 29426 51714 29438
rect 51662 29362 51714 29374
rect 51998 29426 52050 29438
rect 53118 29426 53170 29438
rect 52210 29374 52222 29426
rect 52274 29374 52286 29426
rect 51998 29362 52050 29374
rect 53118 29362 53170 29374
rect 53678 29426 53730 29438
rect 53678 29362 53730 29374
rect 54126 29426 54178 29438
rect 54126 29362 54178 29374
rect 54238 29426 54290 29438
rect 62414 29426 62466 29438
rect 54898 29374 54910 29426
rect 54962 29374 54974 29426
rect 55570 29374 55582 29426
rect 55634 29374 55646 29426
rect 58034 29374 58046 29426
rect 58098 29374 58110 29426
rect 58258 29374 58270 29426
rect 58322 29374 58334 29426
rect 59378 29374 59390 29426
rect 59442 29374 59454 29426
rect 59938 29374 59950 29426
rect 60002 29374 60014 29426
rect 60946 29374 60958 29426
rect 61010 29374 61022 29426
rect 61170 29374 61182 29426
rect 61234 29374 61246 29426
rect 62178 29374 62190 29426
rect 62242 29374 62254 29426
rect 54238 29362 54290 29374
rect 62414 29362 62466 29374
rect 62750 29426 62802 29438
rect 62750 29362 62802 29374
rect 62974 29426 63026 29438
rect 62974 29362 63026 29374
rect 65774 29426 65826 29438
rect 65774 29362 65826 29374
rect 66222 29426 66274 29438
rect 72482 29374 72494 29426
rect 72546 29374 72558 29426
rect 74274 29374 74286 29426
rect 74338 29374 74350 29426
rect 74834 29374 74846 29426
rect 74898 29374 74910 29426
rect 66222 29362 66274 29374
rect 7422 29314 7474 29326
rect 5282 29262 5294 29314
rect 5346 29262 5358 29314
rect 7422 29250 7474 29262
rect 11342 29314 11394 29326
rect 11342 29250 11394 29262
rect 11790 29314 11842 29326
rect 16606 29314 16658 29326
rect 15362 29262 15374 29314
rect 15426 29262 15438 29314
rect 11790 29250 11842 29262
rect 16606 29250 16658 29262
rect 19742 29314 19794 29326
rect 19742 29250 19794 29262
rect 28030 29314 28082 29326
rect 28030 29250 28082 29262
rect 28590 29314 28642 29326
rect 35758 29314 35810 29326
rect 30034 29262 30046 29314
rect 30098 29262 30110 29314
rect 31490 29262 31502 29314
rect 31554 29262 31566 29314
rect 33170 29262 33182 29314
rect 33234 29262 33246 29314
rect 28590 29250 28642 29262
rect 35758 29250 35810 29262
rect 41246 29314 41298 29326
rect 41246 29250 41298 29262
rect 41694 29314 41746 29326
rect 52894 29314 52946 29326
rect 45938 29262 45950 29314
rect 46002 29262 46014 29314
rect 41694 29250 41746 29262
rect 52894 29250 52946 29262
rect 53902 29314 53954 29326
rect 53902 29250 53954 29262
rect 67902 29314 67954 29326
rect 67902 29250 67954 29262
rect 69694 29314 69746 29326
rect 69694 29250 69746 29262
rect 73838 29314 73890 29326
rect 77746 29262 77758 29314
rect 77810 29262 77822 29314
rect 73838 29250 73890 29262
rect 6078 29202 6130 29214
rect 6078 29138 6130 29150
rect 13246 29202 13298 29214
rect 32398 29202 32450 29214
rect 49758 29202 49810 29214
rect 59614 29202 59666 29214
rect 31602 29150 31614 29202
rect 31666 29150 31678 29202
rect 36530 29150 36542 29202
rect 36594 29150 36606 29202
rect 58258 29150 58270 29202
rect 58322 29150 58334 29202
rect 13246 29138 13298 29150
rect 32398 29138 32450 29150
rect 49758 29138 49810 29150
rect 59614 29138 59666 29150
rect 66558 29202 66610 29214
rect 66558 29138 66610 29150
rect 70478 29202 70530 29214
rect 70478 29138 70530 29150
rect 1344 29034 78624 29068
rect 1344 28982 10874 29034
rect 10926 28982 10978 29034
rect 11030 28982 11082 29034
rect 11134 28982 30194 29034
rect 30246 28982 30298 29034
rect 30350 28982 30402 29034
rect 30454 28982 49514 29034
rect 49566 28982 49618 29034
rect 49670 28982 49722 29034
rect 49774 28982 68834 29034
rect 68886 28982 68938 29034
rect 68990 28982 69042 29034
rect 69094 28982 78624 29034
rect 1344 28948 78624 28982
rect 13694 28866 13746 28878
rect 24670 28866 24722 28878
rect 21970 28814 21982 28866
rect 22034 28814 22046 28866
rect 13694 28802 13746 28814
rect 24670 28802 24722 28814
rect 25454 28866 25506 28878
rect 25454 28802 25506 28814
rect 25790 28866 25842 28878
rect 25790 28802 25842 28814
rect 35198 28866 35250 28878
rect 35198 28802 35250 28814
rect 40350 28866 40402 28878
rect 40350 28802 40402 28814
rect 40686 28866 40738 28878
rect 40686 28802 40738 28814
rect 48302 28866 48354 28878
rect 48302 28802 48354 28814
rect 54574 28866 54626 28878
rect 54574 28802 54626 28814
rect 57486 28866 57538 28878
rect 57486 28802 57538 28814
rect 59614 28866 59666 28878
rect 59614 28802 59666 28814
rect 59950 28866 60002 28878
rect 59950 28802 60002 28814
rect 66334 28866 66386 28878
rect 66334 28802 66386 28814
rect 66670 28866 66722 28878
rect 66670 28802 66722 28814
rect 13806 28754 13858 28766
rect 5058 28702 5070 28754
rect 5122 28702 5134 28754
rect 7858 28702 7870 28754
rect 7922 28702 7934 28754
rect 9986 28702 9998 28754
rect 10050 28702 10062 28754
rect 13806 28690 13858 28702
rect 14702 28754 14754 28766
rect 20750 28754 20802 28766
rect 20178 28702 20190 28754
rect 20242 28702 20254 28754
rect 14702 28690 14754 28702
rect 20750 28690 20802 28702
rect 30270 28754 30322 28766
rect 38558 28754 38610 28766
rect 31266 28702 31278 28754
rect 31330 28702 31342 28754
rect 37650 28702 37662 28754
rect 37714 28702 37726 28754
rect 30270 28690 30322 28702
rect 38558 28690 38610 28702
rect 40910 28754 40962 28766
rect 42366 28754 42418 28766
rect 41570 28702 41582 28754
rect 41634 28702 41646 28754
rect 40910 28690 40962 28702
rect 42366 28690 42418 28702
rect 42814 28754 42866 28766
rect 53006 28754 53058 28766
rect 46050 28702 46062 28754
rect 46114 28702 46126 28754
rect 49970 28702 49982 28754
rect 50034 28702 50046 28754
rect 42814 28690 42866 28702
rect 53006 28690 53058 28702
rect 54798 28754 54850 28766
rect 54798 28690 54850 28702
rect 58046 28754 58098 28766
rect 58046 28690 58098 28702
rect 58942 28754 58994 28766
rect 72718 28754 72770 28766
rect 61506 28702 61518 28754
rect 61570 28702 61582 28754
rect 58942 28690 58994 28702
rect 72718 28690 72770 28702
rect 75406 28754 75458 28766
rect 75406 28690 75458 28702
rect 18286 28642 18338 28654
rect 21310 28642 21362 28654
rect 24894 28642 24946 28654
rect 26238 28642 26290 28654
rect 34526 28642 34578 28654
rect 2258 28590 2270 28642
rect 2322 28590 2334 28642
rect 2930 28590 2942 28642
rect 2994 28590 3006 28642
rect 5842 28590 5854 28642
rect 5906 28590 5918 28642
rect 7074 28590 7086 28642
rect 7138 28590 7150 28642
rect 14242 28590 14254 28642
rect 14306 28590 14318 28642
rect 16146 28590 16158 28642
rect 16210 28590 16222 28642
rect 17042 28590 17054 28642
rect 17106 28590 17118 28642
rect 19058 28590 19070 28642
rect 19122 28590 19134 28642
rect 19618 28590 19630 28642
rect 19682 28590 19694 28642
rect 21634 28590 21646 28642
rect 21698 28590 21710 28642
rect 23874 28590 23886 28642
rect 23938 28590 23950 28642
rect 25778 28590 25790 28642
rect 25842 28590 25854 28642
rect 27906 28590 27918 28642
rect 27970 28590 27982 28642
rect 29810 28590 29822 28642
rect 29874 28590 29886 28642
rect 30034 28590 30046 28642
rect 30098 28590 30110 28642
rect 31154 28590 31166 28642
rect 31218 28590 31230 28642
rect 32386 28590 32398 28642
rect 32450 28590 32462 28642
rect 33954 28590 33966 28642
rect 34018 28590 34030 28642
rect 18286 28578 18338 28590
rect 21310 28578 21362 28590
rect 24894 28578 24946 28590
rect 26238 28578 26290 28590
rect 34526 28578 34578 28590
rect 35310 28642 35362 28654
rect 35310 28578 35362 28590
rect 35870 28642 35922 28654
rect 35870 28578 35922 28590
rect 36094 28642 36146 28654
rect 39342 28642 39394 28654
rect 36978 28590 36990 28642
rect 37042 28590 37054 28642
rect 36094 28578 36146 28590
rect 39342 28578 39394 28590
rect 39790 28642 39842 28654
rect 47294 28642 47346 28654
rect 41682 28590 41694 28642
rect 41746 28590 41758 28642
rect 46610 28590 46622 28642
rect 46674 28590 46686 28642
rect 39790 28578 39842 28590
rect 47294 28578 47346 28590
rect 47854 28642 47906 28654
rect 53230 28642 53282 28654
rect 51426 28590 51438 28642
rect 51490 28590 51502 28642
rect 52658 28590 52670 28642
rect 52722 28590 52734 28642
rect 47854 28578 47906 28590
rect 53230 28578 53282 28590
rect 54014 28642 54066 28654
rect 55918 28642 55970 28654
rect 54338 28590 54350 28642
rect 54402 28590 54414 28642
rect 54014 28578 54066 28590
rect 55918 28578 55970 28590
rect 57934 28642 57986 28654
rect 57934 28578 57986 28590
rect 58270 28642 58322 28654
rect 58270 28578 58322 28590
rect 58494 28642 58546 28654
rect 58494 28578 58546 28590
rect 58718 28642 58770 28654
rect 62078 28642 62130 28654
rect 59938 28590 59950 28642
rect 60002 28590 60014 28642
rect 61618 28590 61630 28642
rect 61682 28590 61694 28642
rect 58718 28578 58770 28590
rect 62078 28578 62130 28590
rect 62302 28642 62354 28654
rect 62302 28578 62354 28590
rect 65886 28642 65938 28654
rect 71934 28642 71986 28654
rect 67106 28590 67118 28642
rect 67170 28590 67182 28642
rect 73042 28590 73054 28642
rect 73106 28590 73118 28642
rect 65886 28578 65938 28590
rect 71934 28578 71986 28590
rect 5630 28530 5682 28542
rect 26462 28530 26514 28542
rect 15698 28478 15710 28530
rect 15762 28478 15774 28530
rect 5630 28466 5682 28478
rect 26462 28466 26514 28478
rect 26574 28530 26626 28542
rect 26574 28466 26626 28478
rect 27134 28530 27186 28542
rect 34862 28530 34914 28542
rect 28130 28478 28142 28530
rect 28194 28478 28206 28530
rect 30930 28478 30942 28530
rect 30994 28478 31006 28530
rect 27134 28466 27186 28478
rect 34862 28466 34914 28478
rect 36430 28530 36482 28542
rect 46398 28530 46450 28542
rect 38658 28478 38670 28530
rect 38722 28478 38734 28530
rect 38994 28478 39006 28530
rect 39058 28478 39070 28530
rect 41570 28478 41582 28530
rect 41634 28478 41646 28530
rect 36430 28466 36482 28478
rect 46398 28466 46450 28478
rect 48190 28530 48242 28542
rect 48190 28466 48242 28478
rect 48302 28530 48354 28542
rect 53790 28530 53842 28542
rect 50306 28478 50318 28530
rect 50370 28478 50382 28530
rect 48302 28466 48354 28478
rect 53790 28466 53842 28478
rect 54910 28530 54962 28542
rect 54910 28466 54962 28478
rect 55022 28530 55074 28542
rect 55022 28466 55074 28478
rect 55694 28530 55746 28542
rect 55694 28466 55746 28478
rect 57598 28530 57650 28542
rect 57598 28466 57650 28478
rect 59054 28530 59106 28542
rect 59054 28466 59106 28478
rect 59278 28530 59330 28542
rect 59278 28466 59330 28478
rect 62638 28530 62690 28542
rect 67218 28478 67230 28530
rect 67282 28478 67294 28530
rect 62638 28466 62690 28478
rect 11230 28418 11282 28430
rect 24334 28418 24386 28430
rect 17154 28366 17166 28418
rect 17218 28366 17230 28418
rect 11230 28354 11282 28366
rect 24334 28354 24386 28366
rect 24558 28418 24610 28430
rect 24558 28354 24610 28366
rect 26798 28418 26850 28430
rect 26798 28354 26850 28366
rect 27022 28418 27074 28430
rect 27022 28354 27074 28366
rect 34750 28418 34802 28430
rect 34750 28354 34802 28366
rect 36318 28418 36370 28430
rect 36318 28354 36370 28366
rect 39566 28418 39618 28430
rect 39566 28354 39618 28366
rect 39902 28418 39954 28430
rect 39902 28354 39954 28366
rect 40126 28418 40178 28430
rect 40126 28354 40178 28366
rect 46062 28418 46114 28430
rect 46062 28354 46114 28366
rect 46174 28418 46226 28430
rect 52894 28418 52946 28430
rect 51986 28366 51998 28418
rect 52050 28366 52062 28418
rect 46174 28354 46226 28366
rect 52894 28354 52946 28366
rect 53118 28418 53170 28430
rect 56702 28418 56754 28430
rect 57486 28418 57538 28430
rect 56242 28366 56254 28418
rect 56306 28366 56318 28418
rect 57026 28366 57038 28418
rect 57090 28366 57102 28418
rect 53118 28354 53170 28366
rect 56702 28354 56754 28366
rect 57486 28354 57538 28366
rect 60734 28418 60786 28430
rect 60734 28354 60786 28366
rect 62526 28418 62578 28430
rect 62526 28354 62578 28366
rect 76302 28418 76354 28430
rect 76302 28354 76354 28366
rect 1344 28250 78784 28284
rect 1344 28198 20534 28250
rect 20586 28198 20638 28250
rect 20690 28198 20742 28250
rect 20794 28198 39854 28250
rect 39906 28198 39958 28250
rect 40010 28198 40062 28250
rect 40114 28198 59174 28250
rect 59226 28198 59278 28250
rect 59330 28198 59382 28250
rect 59434 28198 78494 28250
rect 78546 28198 78598 28250
rect 78650 28198 78702 28250
rect 78754 28198 78784 28250
rect 1344 28164 78784 28198
rect 5854 28082 5906 28094
rect 5854 28018 5906 28030
rect 9662 28082 9714 28094
rect 19854 28082 19906 28094
rect 15026 28030 15038 28082
rect 15090 28030 15102 28082
rect 17714 28030 17726 28082
rect 17778 28030 17790 28082
rect 19282 28030 19294 28082
rect 19346 28030 19358 28082
rect 9662 28018 9714 28030
rect 19854 28018 19906 28030
rect 21758 28082 21810 28094
rect 21758 28018 21810 28030
rect 23326 28082 23378 28094
rect 23326 28018 23378 28030
rect 24558 28082 24610 28094
rect 27806 28082 27858 28094
rect 25442 28030 25454 28082
rect 25506 28030 25518 28082
rect 24558 28018 24610 28030
rect 27806 28018 27858 28030
rect 28030 28082 28082 28094
rect 28030 28018 28082 28030
rect 28702 28082 28754 28094
rect 34638 28082 34690 28094
rect 33282 28030 33294 28082
rect 33346 28030 33358 28082
rect 34402 28030 34414 28082
rect 34466 28030 34478 28082
rect 28702 28018 28754 28030
rect 34638 28018 34690 28030
rect 35422 28082 35474 28094
rect 41134 28082 41186 28094
rect 38770 28030 38782 28082
rect 38834 28030 38846 28082
rect 35422 28018 35474 28030
rect 41134 28018 41186 28030
rect 43262 28082 43314 28094
rect 43262 28018 43314 28030
rect 43934 28082 43986 28094
rect 43934 28018 43986 28030
rect 44158 28082 44210 28094
rect 44158 28018 44210 28030
rect 44382 28082 44434 28094
rect 44382 28018 44434 28030
rect 48862 28082 48914 28094
rect 48862 28018 48914 28030
rect 49758 28082 49810 28094
rect 49758 28018 49810 28030
rect 49982 28082 50034 28094
rect 51438 28082 51490 28094
rect 50306 28030 50318 28082
rect 50370 28030 50382 28082
rect 49982 28018 50034 28030
rect 51438 28018 51490 28030
rect 54574 28082 54626 28094
rect 61294 28082 61346 28094
rect 60498 28030 60510 28082
rect 60562 28030 60574 28082
rect 54574 28018 54626 28030
rect 61294 28018 61346 28030
rect 61406 28082 61458 28094
rect 74174 28082 74226 28094
rect 72370 28030 72382 28082
rect 72434 28030 72446 28082
rect 72594 28030 72606 28082
rect 72658 28030 72670 28082
rect 61406 28018 61458 28030
rect 74174 28018 74226 28030
rect 11342 27970 11394 27982
rect 20078 27970 20130 27982
rect 4946 27918 4958 27970
rect 5010 27918 5022 27970
rect 5282 27918 5294 27970
rect 5346 27918 5358 27970
rect 10210 27918 10222 27970
rect 10274 27918 10286 27970
rect 10546 27918 10558 27970
rect 10610 27918 10622 27970
rect 18722 27918 18734 27970
rect 18786 27918 18798 27970
rect 11342 27906 11394 27918
rect 20078 27906 20130 27918
rect 21870 27970 21922 27982
rect 21870 27906 21922 27918
rect 22878 27970 22930 27982
rect 22878 27906 22930 27918
rect 23102 27970 23154 27982
rect 23102 27906 23154 27918
rect 24446 27970 24498 27982
rect 34862 27970 34914 27982
rect 25890 27918 25902 27970
rect 25954 27918 25966 27970
rect 32274 27918 32286 27970
rect 32338 27918 32350 27970
rect 33618 27918 33630 27970
rect 33682 27918 33694 27970
rect 24446 27906 24498 27918
rect 34862 27906 34914 27918
rect 38446 27970 38498 27982
rect 38446 27906 38498 27918
rect 39790 27970 39842 27982
rect 39790 27906 39842 27918
rect 40238 27970 40290 27982
rect 40238 27906 40290 27918
rect 41358 27970 41410 27982
rect 41358 27906 41410 27918
rect 42702 27970 42754 27982
rect 42702 27906 42754 27918
rect 42814 27970 42866 27982
rect 70142 27970 70194 27982
rect 48066 27918 48078 27970
rect 48130 27918 48142 27970
rect 49186 27918 49198 27970
rect 49250 27918 49262 27970
rect 50642 27918 50654 27970
rect 50706 27918 50718 27970
rect 59602 27918 59614 27970
rect 59666 27918 59678 27970
rect 42814 27906 42866 27918
rect 70142 27906 70194 27918
rect 71374 27970 71426 27982
rect 75070 27970 75122 27982
rect 73266 27918 73278 27970
rect 73330 27918 73342 27970
rect 71374 27906 71426 27918
rect 75070 27906 75122 27918
rect 11678 27858 11730 27870
rect 4274 27806 4286 27858
rect 4338 27806 4350 27858
rect 11678 27794 11730 27806
rect 15374 27858 15426 27870
rect 19630 27858 19682 27870
rect 17826 27806 17838 27858
rect 17890 27806 17902 27858
rect 18162 27806 18174 27858
rect 18226 27806 18238 27858
rect 15374 27794 15426 27806
rect 19630 27794 19682 27806
rect 20190 27858 20242 27870
rect 20190 27794 20242 27806
rect 20750 27858 20802 27870
rect 20750 27794 20802 27806
rect 23438 27858 23490 27870
rect 28142 27858 28194 27870
rect 25218 27806 25230 27858
rect 25282 27806 25294 27858
rect 26338 27806 26350 27858
rect 26402 27806 26414 27858
rect 23438 27794 23490 27806
rect 28142 27794 28194 27806
rect 29038 27858 29090 27870
rect 29038 27794 29090 27806
rect 30382 27858 30434 27870
rect 30382 27794 30434 27806
rect 30494 27858 30546 27870
rect 30494 27794 30546 27806
rect 30718 27858 30770 27870
rect 34974 27858 35026 27870
rect 38334 27858 38386 27870
rect 31490 27806 31502 27858
rect 31554 27806 31566 27858
rect 32162 27806 32174 27858
rect 32226 27806 32238 27858
rect 33730 27806 33742 27858
rect 33794 27806 33806 27858
rect 34178 27806 34190 27858
rect 34242 27806 34254 27858
rect 37986 27806 37998 27858
rect 38050 27806 38062 27858
rect 30718 27794 30770 27806
rect 34974 27794 35026 27806
rect 38334 27794 38386 27806
rect 41470 27858 41522 27870
rect 41470 27794 41522 27806
rect 42478 27858 42530 27870
rect 42478 27794 42530 27806
rect 44494 27858 44546 27870
rect 44494 27794 44546 27806
rect 46958 27858 47010 27870
rect 60174 27858 60226 27870
rect 47730 27806 47742 27858
rect 47794 27806 47806 27858
rect 50866 27806 50878 27858
rect 50930 27806 50942 27858
rect 52098 27806 52110 27858
rect 52162 27806 52174 27858
rect 53666 27806 53678 27858
rect 53730 27806 53742 27858
rect 54898 27806 54910 27858
rect 54962 27806 54974 27858
rect 58706 27806 58718 27858
rect 58770 27806 58782 27858
rect 59042 27806 59054 27858
rect 59106 27806 59118 27858
rect 46958 27794 47010 27806
rect 60174 27794 60226 27806
rect 60734 27858 60786 27870
rect 60734 27794 60786 27806
rect 61182 27858 61234 27870
rect 68574 27858 68626 27870
rect 62066 27806 62078 27858
rect 62130 27806 62142 27858
rect 62514 27806 62526 27858
rect 62578 27806 62590 27858
rect 63410 27806 63422 27858
rect 63474 27806 63486 27858
rect 61182 27794 61234 27806
rect 68574 27794 68626 27806
rect 68686 27858 68738 27870
rect 68686 27794 68738 27806
rect 68910 27858 68962 27870
rect 70702 27858 70754 27870
rect 71150 27858 71202 27870
rect 69122 27806 69134 27858
rect 69186 27806 69198 27858
rect 70354 27806 70366 27858
rect 70418 27806 70430 27858
rect 70914 27806 70926 27858
rect 70978 27806 70990 27858
rect 68910 27794 68962 27806
rect 70702 27794 70754 27806
rect 71150 27794 71202 27806
rect 71262 27858 71314 27870
rect 74734 27858 74786 27870
rect 71586 27806 71598 27858
rect 71650 27806 71662 27858
rect 72818 27806 72830 27858
rect 72882 27806 72894 27858
rect 73154 27806 73166 27858
rect 73218 27806 73230 27858
rect 75618 27806 75630 27858
rect 75682 27806 75694 27858
rect 71262 27794 71314 27806
rect 74734 27794 74786 27806
rect 1934 27746 1986 27758
rect 1934 27682 1986 27694
rect 6414 27746 6466 27758
rect 6414 27682 6466 27694
rect 6862 27746 6914 27758
rect 6862 27682 6914 27694
rect 12126 27746 12178 27758
rect 12126 27682 12178 27694
rect 15598 27746 15650 27758
rect 15598 27682 15650 27694
rect 16270 27746 16322 27758
rect 16270 27682 16322 27694
rect 16830 27746 16882 27758
rect 16830 27682 16882 27694
rect 20526 27746 20578 27758
rect 20526 27682 20578 27694
rect 21086 27746 21138 27758
rect 21086 27682 21138 27694
rect 23998 27746 24050 27758
rect 23998 27682 24050 27694
rect 26798 27746 26850 27758
rect 26798 27682 26850 27694
rect 27358 27746 27410 27758
rect 37102 27746 37154 27758
rect 31714 27694 31726 27746
rect 31778 27694 31790 27746
rect 27358 27682 27410 27694
rect 37102 27682 37154 27694
rect 39342 27746 39394 27758
rect 39342 27682 39394 27694
rect 45054 27746 45106 27758
rect 45054 27682 45106 27694
rect 45390 27746 45442 27758
rect 55246 27746 55298 27758
rect 51874 27694 51886 27746
rect 51938 27694 51950 27746
rect 55010 27694 55022 27746
rect 55074 27694 55086 27746
rect 45390 27682 45442 27694
rect 55246 27682 55298 27694
rect 56702 27746 56754 27758
rect 68798 27746 68850 27758
rect 59266 27694 59278 27746
rect 59330 27694 59342 27746
rect 56702 27682 56754 27694
rect 68798 27682 68850 27694
rect 5518 27634 5570 27646
rect 5518 27570 5570 27582
rect 9998 27634 10050 27646
rect 9998 27570 10050 27582
rect 16494 27634 16546 27646
rect 16494 27570 16546 27582
rect 24670 27634 24722 27646
rect 24670 27570 24722 27582
rect 30830 27634 30882 27646
rect 30830 27570 30882 27582
rect 39118 27634 39170 27646
rect 39118 27570 39170 27582
rect 39678 27634 39730 27646
rect 39678 27570 39730 27582
rect 40126 27634 40178 27646
rect 40126 27570 40178 27582
rect 47294 27634 47346 27646
rect 70030 27634 70082 27646
rect 53554 27582 53566 27634
rect 53618 27582 53630 27634
rect 62290 27582 62302 27634
rect 62354 27582 62366 27634
rect 47294 27570 47346 27582
rect 70030 27570 70082 27582
rect 77982 27634 78034 27646
rect 77982 27570 78034 27582
rect 1344 27466 78624 27500
rect 1344 27414 10874 27466
rect 10926 27414 10978 27466
rect 11030 27414 11082 27466
rect 11134 27414 30194 27466
rect 30246 27414 30298 27466
rect 30350 27414 30402 27466
rect 30454 27414 49514 27466
rect 49566 27414 49618 27466
rect 49670 27414 49722 27466
rect 49774 27414 68834 27466
rect 68886 27414 68938 27466
rect 68990 27414 69042 27466
rect 69094 27414 78624 27466
rect 1344 27380 78624 27414
rect 18286 27298 18338 27310
rect 18286 27234 18338 27246
rect 24782 27298 24834 27310
rect 24782 27234 24834 27246
rect 30382 27298 30434 27310
rect 30382 27234 30434 27246
rect 39006 27298 39058 27310
rect 39006 27234 39058 27246
rect 42366 27298 42418 27310
rect 58830 27298 58882 27310
rect 53442 27246 53454 27298
rect 53506 27246 53518 27298
rect 42366 27234 42418 27246
rect 58830 27234 58882 27246
rect 66222 27298 66274 27310
rect 66222 27234 66274 27246
rect 73726 27298 73778 27310
rect 73726 27234 73778 27246
rect 74398 27298 74450 27310
rect 74398 27234 74450 27246
rect 4510 27186 4562 27198
rect 19070 27186 19122 27198
rect 9538 27134 9550 27186
rect 9602 27134 9614 27186
rect 10770 27134 10782 27186
rect 10834 27134 10846 27186
rect 12898 27134 12910 27186
rect 12962 27134 12974 27186
rect 18498 27134 18510 27186
rect 18562 27134 18574 27186
rect 4510 27122 4562 27134
rect 19070 27122 19122 27134
rect 25118 27186 25170 27198
rect 37550 27186 37602 27198
rect 28354 27134 28366 27186
rect 28418 27134 28430 27186
rect 25118 27122 25170 27134
rect 37550 27122 37602 27134
rect 38222 27186 38274 27198
rect 38222 27122 38274 27134
rect 44942 27186 44994 27198
rect 58942 27186 58994 27198
rect 53554 27134 53566 27186
rect 53618 27134 53630 27186
rect 44942 27122 44994 27134
rect 58942 27122 58994 27134
rect 59390 27186 59442 27198
rect 59390 27122 59442 27134
rect 60622 27186 60674 27198
rect 62066 27134 62078 27186
rect 62130 27134 62142 27186
rect 69346 27134 69358 27186
rect 69410 27134 69422 27186
rect 60622 27122 60674 27134
rect 17390 27074 17442 27086
rect 26350 27074 26402 27086
rect 6738 27022 6750 27074
rect 6802 27022 6814 27074
rect 10098 27022 10110 27074
rect 10162 27022 10174 27074
rect 18610 27022 18622 27074
rect 18674 27022 18686 27074
rect 25778 27022 25790 27074
rect 25842 27022 25854 27074
rect 17390 27010 17442 27022
rect 26350 27010 26402 27022
rect 26686 27074 26738 27086
rect 26686 27010 26738 27022
rect 27022 27074 27074 27086
rect 38558 27074 38610 27086
rect 42702 27074 42754 27086
rect 44270 27074 44322 27086
rect 59278 27074 59330 27086
rect 27570 27022 27582 27074
rect 27634 27022 27646 27074
rect 30818 27022 30830 27074
rect 30882 27022 30894 27074
rect 31714 27022 31726 27074
rect 31778 27022 31790 27074
rect 32498 27022 32510 27074
rect 32562 27022 32574 27074
rect 33954 27022 33966 27074
rect 34018 27022 34030 27074
rect 36082 27022 36094 27074
rect 36146 27022 36158 27074
rect 37874 27022 37886 27074
rect 37938 27022 37950 27074
rect 38770 27022 38782 27074
rect 38834 27022 38846 27074
rect 39330 27022 39342 27074
rect 39394 27022 39406 27074
rect 40226 27022 40238 27074
rect 40290 27022 40302 27074
rect 43474 27022 43486 27074
rect 43538 27022 43550 27074
rect 53442 27022 53454 27074
rect 53506 27022 53518 27074
rect 54338 27022 54350 27074
rect 54402 27022 54414 27074
rect 27022 27010 27074 27022
rect 38558 27010 38610 27022
rect 42702 27010 42754 27022
rect 44270 27010 44322 27022
rect 59278 27010 59330 27022
rect 59726 27074 59778 27086
rect 66334 27074 66386 27086
rect 74734 27074 74786 27086
rect 61618 27022 61630 27074
rect 61682 27022 61694 27074
rect 62738 27022 62750 27074
rect 62802 27022 62814 27074
rect 66994 27022 67006 27074
rect 67058 27022 67070 27074
rect 67554 27022 67566 27074
rect 67618 27022 67630 27074
rect 69234 27022 69246 27074
rect 69298 27022 69310 27074
rect 70354 27022 70366 27074
rect 70418 27022 70430 27074
rect 72146 27022 72158 27074
rect 72210 27022 72222 27074
rect 73714 27022 73726 27074
rect 73778 27022 73790 27074
rect 75506 27022 75518 27074
rect 75570 27022 75582 27074
rect 76402 27022 76414 27074
rect 76466 27022 76478 27074
rect 59726 27010 59778 27022
rect 66334 27010 66386 27022
rect 74734 27010 74786 27022
rect 3166 26962 3218 26974
rect 16494 26962 16546 26974
rect 7410 26910 7422 26962
rect 7474 26910 7486 26962
rect 3166 26898 3218 26910
rect 16494 26898 16546 26910
rect 16830 26962 16882 26974
rect 16830 26898 16882 26910
rect 17166 26962 17218 26974
rect 17166 26898 17218 26910
rect 21534 26962 21586 26974
rect 21534 26898 21586 26910
rect 21646 26962 21698 26974
rect 21646 26898 21698 26910
rect 21758 26962 21810 26974
rect 22206 26962 22258 26974
rect 21858 26910 21870 26962
rect 21922 26959 21934 26962
rect 22082 26959 22094 26962
rect 21922 26913 22094 26959
rect 21922 26910 21934 26913
rect 22082 26910 22094 26913
rect 22146 26910 22158 26962
rect 21758 26898 21810 26910
rect 22206 26898 22258 26910
rect 22654 26962 22706 26974
rect 22654 26898 22706 26910
rect 24558 26962 24610 26974
rect 24558 26898 24610 26910
rect 26462 26962 26514 26974
rect 26462 26898 26514 26910
rect 30382 26962 30434 26974
rect 30382 26898 30434 26910
rect 30494 26962 30546 26974
rect 39678 26962 39730 26974
rect 31266 26910 31278 26962
rect 31330 26910 31342 26962
rect 32274 26910 32286 26962
rect 32338 26910 32350 26962
rect 35522 26910 35534 26962
rect 35586 26910 35598 26962
rect 30494 26898 30546 26910
rect 39678 26898 39730 26910
rect 39902 26962 39954 26974
rect 39902 26898 39954 26910
rect 41358 26962 41410 26974
rect 41358 26898 41410 26910
rect 41694 26962 41746 26974
rect 44830 26962 44882 26974
rect 43362 26910 43374 26962
rect 43426 26910 43438 26962
rect 43922 26910 43934 26962
rect 43986 26910 43998 26962
rect 41694 26898 41746 26910
rect 44830 26898 44882 26910
rect 45502 26962 45554 26974
rect 59614 26962 59666 26974
rect 45826 26910 45838 26962
rect 45890 26910 45902 26962
rect 61282 26910 61294 26962
rect 61346 26910 61358 26962
rect 66546 26910 66558 26962
rect 66610 26910 66622 26962
rect 70018 26910 70030 26962
rect 70082 26910 70094 26962
rect 73154 26910 73166 26962
rect 73218 26910 73230 26962
rect 75282 26910 75294 26962
rect 75346 26910 75358 26962
rect 45502 26898 45554 26910
rect 59614 26898 59666 26910
rect 2830 26850 2882 26862
rect 22766 26850 22818 26862
rect 17714 26798 17726 26850
rect 17778 26798 17790 26850
rect 2830 26786 2882 26798
rect 22766 26786 22818 26798
rect 22990 26850 23042 26862
rect 22990 26786 23042 26798
rect 26910 26850 26962 26862
rect 38110 26850 38162 26862
rect 31826 26798 31838 26850
rect 31890 26798 31902 26850
rect 32722 26798 32734 26850
rect 32786 26798 32798 26850
rect 26910 26786 26962 26798
rect 38110 26786 38162 26798
rect 39342 26850 39394 26862
rect 39342 26786 39394 26798
rect 39790 26850 39842 26862
rect 39790 26786 39842 26798
rect 40798 26850 40850 26862
rect 40798 26786 40850 26798
rect 45054 26850 45106 26862
rect 45054 26786 45106 26798
rect 48414 26850 48466 26862
rect 48414 26786 48466 26798
rect 50430 26850 50482 26862
rect 50430 26786 50482 26798
rect 76190 26850 76242 26862
rect 76190 26786 76242 26798
rect 1344 26682 78784 26716
rect 1344 26630 20534 26682
rect 20586 26630 20638 26682
rect 20690 26630 20742 26682
rect 20794 26630 39854 26682
rect 39906 26630 39958 26682
rect 40010 26630 40062 26682
rect 40114 26630 59174 26682
rect 59226 26630 59278 26682
rect 59330 26630 59382 26682
rect 59434 26630 78494 26682
rect 78546 26630 78598 26682
rect 78650 26630 78702 26682
rect 78754 26630 78784 26682
rect 1344 26596 78784 26630
rect 7310 26514 7362 26526
rect 11342 26514 11394 26526
rect 10994 26462 11006 26514
rect 11058 26462 11070 26514
rect 7310 26450 7362 26462
rect 11342 26450 11394 26462
rect 11790 26514 11842 26526
rect 23662 26514 23714 26526
rect 22082 26462 22094 26514
rect 22146 26462 22158 26514
rect 11790 26450 11842 26462
rect 23662 26450 23714 26462
rect 25902 26514 25954 26526
rect 25902 26450 25954 26462
rect 32398 26514 32450 26526
rect 38782 26514 38834 26526
rect 36642 26462 36654 26514
rect 36706 26462 36718 26514
rect 32398 26450 32450 26462
rect 38782 26450 38834 26462
rect 42702 26514 42754 26526
rect 42702 26450 42754 26462
rect 44606 26514 44658 26526
rect 44606 26450 44658 26462
rect 46286 26514 46338 26526
rect 46286 26450 46338 26462
rect 50542 26514 50594 26526
rect 50542 26450 50594 26462
rect 50766 26514 50818 26526
rect 50766 26450 50818 26462
rect 52782 26514 52834 26526
rect 52782 26450 52834 26462
rect 54126 26514 54178 26526
rect 54126 26450 54178 26462
rect 57038 26514 57090 26526
rect 57038 26450 57090 26462
rect 58606 26514 58658 26526
rect 58606 26450 58658 26462
rect 59614 26514 59666 26526
rect 59614 26450 59666 26462
rect 59950 26514 60002 26526
rect 59950 26450 60002 26462
rect 61630 26514 61682 26526
rect 61630 26450 61682 26462
rect 63086 26514 63138 26526
rect 63086 26450 63138 26462
rect 65326 26514 65378 26526
rect 65326 26450 65378 26462
rect 66110 26514 66162 26526
rect 70018 26462 70030 26514
rect 70082 26462 70094 26514
rect 73154 26462 73166 26514
rect 73218 26462 73230 26514
rect 66110 26450 66162 26462
rect 16494 26402 16546 26414
rect 26126 26402 26178 26414
rect 2482 26350 2494 26402
rect 2546 26350 2558 26402
rect 8418 26350 8430 26402
rect 8482 26350 8494 26402
rect 8866 26350 8878 26402
rect 8930 26350 8942 26402
rect 20626 26350 20638 26402
rect 20690 26350 20702 26402
rect 16494 26338 16546 26350
rect 26126 26338 26178 26350
rect 26238 26402 26290 26414
rect 32174 26402 32226 26414
rect 31154 26350 31166 26402
rect 31218 26350 31230 26402
rect 26238 26338 26290 26350
rect 32174 26338 32226 26350
rect 33742 26402 33794 26414
rect 37886 26402 37938 26414
rect 36754 26350 36766 26402
rect 36818 26350 36830 26402
rect 33742 26338 33794 26350
rect 37886 26338 37938 26350
rect 45166 26402 45218 26414
rect 51102 26402 51154 26414
rect 48962 26350 48974 26402
rect 49026 26350 49038 26402
rect 45166 26338 45218 26350
rect 51102 26338 51154 26350
rect 57262 26402 57314 26414
rect 57262 26338 57314 26350
rect 58942 26402 58994 26414
rect 58942 26338 58994 26350
rect 59166 26402 59218 26414
rect 59166 26338 59218 26350
rect 59502 26402 59554 26414
rect 63310 26402 63362 26414
rect 61954 26350 61966 26402
rect 62018 26350 62030 26402
rect 59502 26338 59554 26350
rect 63310 26338 63362 26350
rect 63422 26402 63474 26414
rect 63422 26338 63474 26350
rect 65438 26402 65490 26414
rect 72494 26402 72546 26414
rect 71026 26350 71038 26402
rect 71090 26350 71102 26402
rect 73602 26350 73614 26402
rect 73666 26350 73678 26402
rect 74946 26350 74958 26402
rect 75010 26350 75022 26402
rect 65438 26338 65490 26350
rect 72494 26338 72546 26350
rect 7758 26290 7810 26302
rect 1810 26238 1822 26290
rect 1874 26238 1886 26290
rect 7074 26238 7086 26290
rect 7138 26238 7150 26290
rect 7758 26226 7810 26238
rect 8094 26290 8146 26302
rect 19854 26290 19906 26302
rect 27134 26290 27186 26302
rect 14914 26238 14926 26290
rect 14978 26238 14990 26290
rect 16818 26238 16830 26290
rect 16882 26238 16894 26290
rect 18050 26238 18062 26290
rect 18114 26238 18126 26290
rect 19394 26238 19406 26290
rect 19458 26238 19470 26290
rect 21186 26238 21198 26290
rect 21250 26238 21262 26290
rect 21746 26238 21758 26290
rect 21810 26238 21822 26290
rect 24322 26238 24334 26290
rect 24386 26238 24398 26290
rect 8094 26226 8146 26238
rect 19854 26226 19906 26238
rect 27134 26226 27186 26238
rect 27470 26290 27522 26302
rect 29374 26290 29426 26302
rect 37998 26290 38050 26302
rect 28914 26238 28926 26290
rect 28978 26238 28990 26290
rect 31042 26238 31054 26290
rect 31106 26238 31118 26290
rect 33058 26238 33070 26290
rect 33122 26238 33134 26290
rect 35298 26238 35310 26290
rect 35362 26238 35374 26290
rect 27470 26226 27522 26238
rect 29374 26226 29426 26238
rect 37998 26226 38050 26238
rect 38446 26290 38498 26302
rect 38446 26226 38498 26238
rect 38670 26290 38722 26302
rect 42478 26290 42530 26302
rect 40114 26238 40126 26290
rect 40178 26238 40190 26290
rect 38670 26226 38722 26238
rect 42478 26226 42530 26238
rect 42702 26290 42754 26302
rect 42702 26226 42754 26238
rect 43038 26290 43090 26302
rect 43038 26226 43090 26238
rect 45054 26290 45106 26302
rect 45054 26226 45106 26238
rect 45278 26290 45330 26302
rect 50654 26290 50706 26302
rect 46050 26238 46062 26290
rect 46114 26238 46126 26290
rect 49074 26238 49086 26290
rect 49138 26238 49150 26290
rect 50194 26238 50206 26290
rect 50258 26238 50270 26290
rect 45278 26226 45330 26238
rect 50654 26226 50706 26238
rect 50878 26290 50930 26302
rect 50878 26226 50930 26238
rect 52558 26290 52610 26302
rect 52558 26226 52610 26238
rect 52670 26290 52722 26302
rect 52670 26226 52722 26238
rect 52894 26290 52946 26302
rect 57374 26290 57426 26302
rect 53106 26238 53118 26290
rect 53170 26238 53182 26290
rect 52894 26226 52946 26238
rect 57374 26226 57426 26238
rect 59726 26290 59778 26302
rect 59726 26226 59778 26238
rect 64878 26290 64930 26302
rect 64878 26226 64930 26238
rect 65214 26290 65266 26302
rect 65214 26226 65266 26238
rect 65886 26290 65938 26302
rect 65886 26226 65938 26238
rect 65998 26290 66050 26302
rect 65998 26226 66050 26238
rect 66222 26290 66274 26302
rect 66434 26238 66446 26290
rect 66498 26238 66510 26290
rect 66770 26238 66782 26290
rect 66834 26238 66846 26290
rect 68114 26238 68126 26290
rect 68178 26238 68190 26290
rect 68562 26238 68574 26290
rect 68626 26238 68638 26290
rect 69570 26238 69582 26290
rect 69634 26238 69646 26290
rect 71474 26238 71486 26290
rect 71538 26238 71550 26290
rect 72818 26238 72830 26290
rect 72882 26238 72894 26290
rect 73154 26238 73166 26290
rect 73218 26238 73230 26290
rect 74274 26238 74286 26290
rect 74338 26238 74350 26290
rect 66222 26226 66274 26238
rect 9662 26178 9714 26190
rect 16606 26178 16658 26190
rect 18734 26178 18786 26190
rect 4610 26126 4622 26178
rect 4674 26126 4686 26178
rect 16034 26126 16046 26178
rect 16098 26126 16110 26178
rect 18386 26126 18398 26178
rect 18450 26126 18462 26178
rect 9662 26114 9714 26126
rect 16606 26114 16658 26126
rect 18734 26114 18786 26126
rect 19182 26178 19234 26190
rect 22654 26178 22706 26190
rect 20962 26126 20974 26178
rect 21026 26126 21038 26178
rect 19182 26114 19234 26126
rect 22654 26114 22706 26126
rect 25678 26178 25730 26190
rect 28030 26178 28082 26190
rect 30718 26178 30770 26190
rect 37438 26178 37490 26190
rect 26674 26126 26686 26178
rect 26738 26126 26750 26178
rect 28578 26126 28590 26178
rect 28642 26126 28654 26178
rect 29810 26126 29822 26178
rect 29874 26126 29886 26178
rect 31266 26126 31278 26178
rect 31330 26126 31342 26178
rect 32498 26126 32510 26178
rect 32562 26126 32574 26178
rect 25678 26114 25730 26126
rect 28030 26114 28082 26126
rect 30718 26114 30770 26126
rect 37438 26114 37490 26126
rect 37550 26178 37602 26190
rect 43486 26178 43538 26190
rect 39666 26126 39678 26178
rect 39730 26126 39742 26178
rect 37550 26114 37602 26126
rect 43486 26114 43538 26126
rect 48190 26178 48242 26190
rect 64542 26178 64594 26190
rect 49522 26126 49534 26178
rect 49586 26126 49598 26178
rect 77074 26126 77086 26178
rect 77138 26126 77150 26178
rect 48190 26114 48242 26126
rect 64542 26114 64594 26126
rect 19070 26066 19122 26078
rect 19070 26002 19122 26014
rect 22430 26066 22482 26078
rect 46398 26066 46450 26078
rect 45714 26014 45726 26066
rect 45778 26014 45790 26066
rect 22430 26002 22482 26014
rect 46398 26002 46450 26014
rect 58830 26066 58882 26078
rect 58830 26002 58882 26014
rect 1344 25898 78624 25932
rect 1344 25846 10874 25898
rect 10926 25846 10978 25898
rect 11030 25846 11082 25898
rect 11134 25846 30194 25898
rect 30246 25846 30298 25898
rect 30350 25846 30402 25898
rect 30454 25846 49514 25898
rect 49566 25846 49618 25898
rect 49670 25846 49722 25898
rect 49774 25846 68834 25898
rect 68886 25846 68938 25898
rect 68990 25846 69042 25898
rect 69094 25846 78624 25898
rect 1344 25812 78624 25846
rect 1934 25730 1986 25742
rect 1934 25666 1986 25678
rect 11678 25730 11730 25742
rect 11678 25666 11730 25678
rect 12014 25730 12066 25742
rect 12014 25666 12066 25678
rect 27806 25730 27858 25742
rect 50094 25730 50146 25742
rect 33954 25678 33966 25730
rect 34018 25678 34030 25730
rect 27806 25666 27858 25678
rect 50094 25666 50146 25678
rect 76302 25730 76354 25742
rect 76302 25666 76354 25678
rect 76638 25730 76690 25742
rect 76638 25666 76690 25678
rect 24110 25618 24162 25630
rect 15474 25566 15486 25618
rect 15538 25566 15550 25618
rect 18498 25566 18510 25618
rect 18562 25566 18574 25618
rect 19842 25566 19854 25618
rect 19906 25566 19918 25618
rect 24110 25554 24162 25566
rect 27918 25618 27970 25630
rect 27918 25554 27970 25566
rect 30270 25618 30322 25630
rect 35758 25618 35810 25630
rect 35186 25566 35198 25618
rect 35250 25566 35262 25618
rect 30270 25554 30322 25566
rect 35758 25554 35810 25566
rect 39006 25618 39058 25630
rect 43822 25618 43874 25630
rect 40226 25566 40238 25618
rect 40290 25566 40302 25618
rect 39006 25554 39058 25566
rect 43822 25554 43874 25566
rect 44270 25618 44322 25630
rect 44270 25554 44322 25566
rect 46398 25618 46450 25630
rect 46398 25554 46450 25566
rect 47294 25618 47346 25630
rect 55582 25618 55634 25630
rect 48738 25566 48750 25618
rect 48802 25566 48814 25618
rect 49746 25566 49758 25618
rect 49810 25566 49822 25618
rect 47294 25554 47346 25566
rect 55582 25554 55634 25566
rect 58942 25618 58994 25630
rect 67454 25618 67506 25630
rect 73726 25618 73778 25630
rect 66210 25566 66222 25618
rect 66274 25566 66286 25618
rect 69682 25566 69694 25618
rect 69746 25566 69758 25618
rect 58942 25554 58994 25566
rect 67454 25554 67506 25566
rect 73726 25554 73778 25566
rect 77982 25618 78034 25630
rect 77982 25554 78034 25566
rect 11118 25506 11170 25518
rect 20750 25506 20802 25518
rect 24222 25506 24274 25518
rect 26350 25506 26402 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 12786 25454 12798 25506
rect 12850 25454 12862 25506
rect 14914 25454 14926 25506
rect 14978 25454 14990 25506
rect 16034 25454 16046 25506
rect 16098 25454 16110 25506
rect 16706 25454 16718 25506
rect 16770 25454 16782 25506
rect 17938 25454 17950 25506
rect 18002 25454 18014 25506
rect 20066 25454 20078 25506
rect 20130 25454 20142 25506
rect 21634 25454 21646 25506
rect 21698 25454 21710 25506
rect 23538 25454 23550 25506
rect 23602 25454 23614 25506
rect 24994 25454 25006 25506
rect 25058 25454 25070 25506
rect 11118 25442 11170 25454
rect 20750 25442 20802 25454
rect 24222 25442 24274 25454
rect 26350 25442 26402 25454
rect 27470 25506 27522 25518
rect 33406 25506 33458 25518
rect 28130 25454 28142 25506
rect 28194 25454 28206 25506
rect 27470 25442 27522 25454
rect 33406 25442 33458 25454
rect 33630 25506 33682 25518
rect 38446 25506 38498 25518
rect 34850 25454 34862 25506
rect 34914 25454 34926 25506
rect 33630 25442 33682 25454
rect 38446 25442 38498 25454
rect 40126 25506 40178 25518
rect 44830 25506 44882 25518
rect 40338 25454 40350 25506
rect 40402 25454 40414 25506
rect 40126 25442 40178 25454
rect 44830 25442 44882 25454
rect 45166 25506 45218 25518
rect 45166 25442 45218 25454
rect 45390 25506 45442 25518
rect 48078 25506 48130 25518
rect 50430 25506 50482 25518
rect 46834 25454 46846 25506
rect 46898 25454 46910 25506
rect 48290 25454 48302 25506
rect 48354 25454 48366 25506
rect 49410 25454 49422 25506
rect 49474 25454 49486 25506
rect 45390 25442 45442 25454
rect 48078 25442 48130 25454
rect 50430 25442 50482 25454
rect 53230 25506 53282 25518
rect 59838 25506 59890 25518
rect 67342 25506 67394 25518
rect 53666 25454 53678 25506
rect 53730 25454 53742 25506
rect 54562 25454 54574 25506
rect 54626 25454 54638 25506
rect 56242 25454 56254 25506
rect 56306 25454 56318 25506
rect 56914 25454 56926 25506
rect 56978 25454 56990 25506
rect 59602 25454 59614 25506
rect 59666 25454 59678 25506
rect 63410 25454 63422 25506
rect 63474 25454 63486 25506
rect 67106 25454 67118 25506
rect 67170 25454 67182 25506
rect 68338 25454 68350 25506
rect 68402 25454 68414 25506
rect 69234 25454 69246 25506
rect 69298 25454 69310 25506
rect 71586 25454 71598 25506
rect 71650 25454 71662 25506
rect 71922 25454 71934 25506
rect 71986 25454 71998 25506
rect 72258 25454 72270 25506
rect 72322 25454 72334 25506
rect 73490 25454 73502 25506
rect 73554 25454 73566 25506
rect 75170 25454 75182 25506
rect 75234 25454 75246 25506
rect 53230 25442 53282 25454
rect 59838 25442 59890 25454
rect 67342 25442 67394 25454
rect 13694 25394 13746 25406
rect 26014 25394 26066 25406
rect 12562 25342 12574 25394
rect 12626 25342 12638 25394
rect 22306 25342 22318 25394
rect 22370 25342 22382 25394
rect 13694 25330 13746 25342
rect 26014 25330 26066 25342
rect 26910 25394 26962 25406
rect 29262 25394 29314 25406
rect 27122 25342 27134 25394
rect 27186 25342 27198 25394
rect 26910 25330 26962 25342
rect 29262 25330 29314 25342
rect 29374 25394 29426 25406
rect 29374 25330 29426 25342
rect 38894 25394 38946 25406
rect 38894 25330 38946 25342
rect 39118 25394 39170 25406
rect 39118 25330 39170 25342
rect 39678 25394 39730 25406
rect 39678 25330 39730 25342
rect 47742 25394 47794 25406
rect 47742 25330 47794 25342
rect 47854 25394 47906 25406
rect 54126 25394 54178 25406
rect 67790 25394 67842 25406
rect 48626 25342 48638 25394
rect 48690 25342 48702 25394
rect 50754 25342 50766 25394
rect 50818 25342 50830 25394
rect 54786 25342 54798 25394
rect 54850 25342 54862 25394
rect 57138 25342 57150 25394
rect 57202 25342 57214 25394
rect 64082 25342 64094 25394
rect 64146 25342 64158 25394
rect 69346 25342 69358 25394
rect 69410 25342 69422 25394
rect 73938 25342 73950 25394
rect 74002 25342 74014 25394
rect 76850 25342 76862 25394
rect 76914 25342 76926 25394
rect 77410 25342 77422 25394
rect 77474 25342 77486 25394
rect 47854 25330 47906 25342
rect 54126 25330 54178 25342
rect 67790 25330 67842 25342
rect 4846 25282 4898 25294
rect 4846 25218 4898 25230
rect 10222 25282 10274 25294
rect 10222 25218 10274 25230
rect 10782 25282 10834 25294
rect 10782 25218 10834 25230
rect 28590 25282 28642 25294
rect 28590 25218 28642 25230
rect 29038 25282 29090 25294
rect 29038 25218 29090 25230
rect 29934 25282 29986 25294
rect 29934 25218 29986 25230
rect 33070 25282 33122 25294
rect 33070 25218 33122 25230
rect 37214 25282 37266 25294
rect 37214 25218 37266 25230
rect 37550 25282 37602 25294
rect 37550 25218 37602 25230
rect 38222 25282 38274 25294
rect 38222 25218 38274 25230
rect 39902 25282 39954 25294
rect 39902 25218 39954 25230
rect 40910 25282 40962 25294
rect 40910 25218 40962 25230
rect 41806 25282 41858 25294
rect 41806 25218 41858 25230
rect 45054 25282 45106 25294
rect 45054 25218 45106 25230
rect 49870 25282 49922 25294
rect 49870 25218 49922 25230
rect 58382 25282 58434 25294
rect 58382 25218 58434 25230
rect 67566 25282 67618 25294
rect 67566 25218 67618 25230
rect 68574 25282 68626 25294
rect 68574 25218 68626 25230
rect 1344 25114 78784 25148
rect 1344 25062 20534 25114
rect 20586 25062 20638 25114
rect 20690 25062 20742 25114
rect 20794 25062 39854 25114
rect 39906 25062 39958 25114
rect 40010 25062 40062 25114
rect 40114 25062 59174 25114
rect 59226 25062 59278 25114
rect 59330 25062 59382 25114
rect 59434 25062 78494 25114
rect 78546 25062 78598 25114
rect 78650 25062 78702 25114
rect 78754 25062 78784 25114
rect 1344 25028 78784 25062
rect 3726 24946 3778 24958
rect 26014 24946 26066 24958
rect 9874 24894 9886 24946
rect 9938 24894 9950 24946
rect 3726 24882 3778 24894
rect 26014 24882 26066 24894
rect 27246 24946 27298 24958
rect 27246 24882 27298 24894
rect 28926 24946 28978 24958
rect 28926 24882 28978 24894
rect 29710 24946 29762 24958
rect 38782 24946 38834 24958
rect 47518 24946 47570 24958
rect 37090 24894 37102 24946
rect 37154 24894 37166 24946
rect 46610 24894 46622 24946
rect 46674 24894 46686 24946
rect 29710 24882 29762 24894
rect 38782 24882 38834 24894
rect 47518 24882 47570 24894
rect 49534 24946 49586 24958
rect 49534 24882 49586 24894
rect 52670 24946 52722 24958
rect 52670 24882 52722 24894
rect 53006 24946 53058 24958
rect 53006 24882 53058 24894
rect 55134 24946 55186 24958
rect 55134 24882 55186 24894
rect 59278 24946 59330 24958
rect 59278 24882 59330 24894
rect 63870 24946 63922 24958
rect 69806 24946 69858 24958
rect 69122 24894 69134 24946
rect 69186 24894 69198 24946
rect 63870 24882 63922 24894
rect 69806 24882 69858 24894
rect 72158 24946 72210 24958
rect 72158 24882 72210 24894
rect 74622 24946 74674 24958
rect 74622 24882 74674 24894
rect 19630 24834 19682 24846
rect 4722 24782 4734 24834
rect 4786 24782 4798 24834
rect 5506 24782 5518 24834
rect 5570 24782 5582 24834
rect 14578 24782 14590 24834
rect 14642 24782 14654 24834
rect 14802 24782 14814 24834
rect 14866 24782 14878 24834
rect 15474 24782 15486 24834
rect 15538 24782 15550 24834
rect 17490 24782 17502 24834
rect 17554 24782 17566 24834
rect 19630 24770 19682 24782
rect 19742 24834 19794 24846
rect 19742 24770 19794 24782
rect 28142 24834 28194 24846
rect 37550 24834 37602 24846
rect 41358 24834 41410 24846
rect 31826 24782 31838 24834
rect 31890 24782 31902 24834
rect 40002 24782 40014 24834
rect 40066 24782 40078 24834
rect 28142 24770 28194 24782
rect 37550 24770 37602 24782
rect 41358 24770 41410 24782
rect 45390 24834 45442 24846
rect 57934 24834 57986 24846
rect 45826 24782 45838 24834
rect 45890 24782 45902 24834
rect 45390 24770 45442 24782
rect 57934 24770 57986 24782
rect 58382 24834 58434 24846
rect 60050 24782 60062 24834
rect 60114 24782 60126 24834
rect 65426 24782 65438 24834
rect 65490 24782 65502 24834
rect 65986 24782 65998 24834
rect 66050 24782 66062 24834
rect 68674 24782 68686 24834
rect 68738 24782 68750 24834
rect 72258 24782 72270 24834
rect 72322 24782 72334 24834
rect 74274 24782 74286 24834
rect 74338 24782 74350 24834
rect 76066 24782 76078 24834
rect 76130 24782 76142 24834
rect 58382 24770 58434 24782
rect 4062 24722 4114 24734
rect 5854 24722 5906 24734
rect 4834 24670 4846 24722
rect 4898 24670 4910 24722
rect 4062 24658 4114 24670
rect 5854 24658 5906 24670
rect 9550 24722 9602 24734
rect 18734 24722 18786 24734
rect 19406 24722 19458 24734
rect 27918 24722 27970 24734
rect 10546 24670 10558 24722
rect 10610 24670 10622 24722
rect 15810 24670 15822 24722
rect 15874 24670 15886 24722
rect 16706 24670 16718 24722
rect 16770 24670 16782 24722
rect 19170 24670 19182 24722
rect 19234 24670 19246 24722
rect 20290 24670 20302 24722
rect 20354 24670 20366 24722
rect 20514 24670 20526 24722
rect 20578 24670 20590 24722
rect 22306 24670 22318 24722
rect 22370 24670 22382 24722
rect 23538 24670 23550 24722
rect 23602 24670 23614 24722
rect 9550 24658 9602 24670
rect 18734 24658 18786 24670
rect 19406 24658 19458 24670
rect 27918 24658 27970 24670
rect 28478 24722 28530 24734
rect 28478 24658 28530 24670
rect 29038 24722 29090 24734
rect 29038 24658 29090 24670
rect 33182 24722 33234 24734
rect 37662 24722 37714 24734
rect 41470 24722 41522 24734
rect 45278 24722 45330 24734
rect 51102 24722 51154 24734
rect 34066 24670 34078 24722
rect 34130 24670 34142 24722
rect 36306 24670 36318 24722
rect 36370 24670 36382 24722
rect 37874 24670 37886 24722
rect 37938 24670 37950 24722
rect 39218 24670 39230 24722
rect 39282 24670 39294 24722
rect 39666 24670 39678 24722
rect 39730 24670 39742 24722
rect 42466 24670 42478 24722
rect 42530 24670 42542 24722
rect 44706 24670 44718 24722
rect 44770 24670 44782 24722
rect 46162 24670 46174 24722
rect 46226 24670 46238 24722
rect 46610 24670 46622 24722
rect 46674 24670 46686 24722
rect 33182 24658 33234 24670
rect 37662 24658 37714 24670
rect 41470 24658 41522 24670
rect 45278 24658 45330 24670
rect 51102 24658 51154 24670
rect 51662 24722 51714 24734
rect 51662 24658 51714 24670
rect 53902 24722 53954 24734
rect 53902 24658 53954 24670
rect 55470 24722 55522 24734
rect 55470 24658 55522 24670
rect 56590 24722 56642 24734
rect 56590 24658 56642 24670
rect 57822 24722 57874 24734
rect 57822 24658 57874 24670
rect 58158 24722 58210 24734
rect 62190 24722 62242 24734
rect 64878 24722 64930 24734
rect 59714 24670 59726 24722
rect 59778 24670 59790 24722
rect 63634 24670 63646 24722
rect 63698 24670 63710 24722
rect 58158 24658 58210 24670
rect 62190 24658 62242 24670
rect 64878 24658 64930 24670
rect 65214 24722 65266 24734
rect 69010 24670 69022 24722
rect 69074 24670 69086 24722
rect 69458 24670 69470 24722
rect 69522 24670 69534 24722
rect 72594 24670 72606 24722
rect 72658 24670 72670 24722
rect 73378 24670 73390 24722
rect 73442 24670 73454 24722
rect 73714 24670 73726 24722
rect 73778 24670 73790 24722
rect 75282 24670 75294 24722
rect 75346 24670 75358 24722
rect 65214 24658 65266 24670
rect 6302 24610 6354 24622
rect 26798 24610 26850 24622
rect 30718 24610 30770 24622
rect 11330 24558 11342 24610
rect 11394 24558 11406 24610
rect 13458 24558 13470 24610
rect 13522 24558 13534 24610
rect 16146 24558 16158 24610
rect 16210 24558 16222 24610
rect 17714 24558 17726 24610
rect 17778 24558 17790 24610
rect 20178 24558 20190 24610
rect 20242 24558 20254 24610
rect 23874 24558 23886 24610
rect 23938 24558 23950 24610
rect 30146 24558 30158 24610
rect 30210 24558 30222 24610
rect 6302 24546 6354 24558
rect 26798 24546 26850 24558
rect 30718 24546 30770 24558
rect 32174 24610 32226 24622
rect 38334 24610 38386 24622
rect 41806 24610 41858 24622
rect 43262 24610 43314 24622
rect 33618 24558 33630 24610
rect 33682 24558 33694 24610
rect 36754 24558 36766 24610
rect 36818 24558 36830 24610
rect 39778 24558 39790 24610
rect 39842 24558 39854 24610
rect 42690 24558 42702 24610
rect 42754 24558 42766 24610
rect 32174 24546 32226 24558
rect 38334 24546 38386 24558
rect 41806 24546 41858 24558
rect 43262 24546 43314 24558
rect 44046 24610 44098 24622
rect 44046 24546 44098 24558
rect 50766 24610 50818 24622
rect 50766 24546 50818 24558
rect 53566 24610 53618 24622
rect 53566 24546 53618 24558
rect 56030 24610 56082 24622
rect 56030 24546 56082 24558
rect 57150 24610 57202 24622
rect 57150 24546 57202 24558
rect 58830 24610 58882 24622
rect 60958 24610 61010 24622
rect 60386 24558 60398 24610
rect 60450 24558 60462 24610
rect 58830 24546 58882 24558
rect 60958 24546 61010 24558
rect 62750 24610 62802 24622
rect 62750 24546 62802 24558
rect 71710 24610 71762 24622
rect 78194 24558 78206 24610
rect 78258 24558 78270 24610
rect 71710 24546 71762 24558
rect 13918 24498 13970 24510
rect 13918 24434 13970 24446
rect 14254 24498 14306 24510
rect 14254 24434 14306 24446
rect 19070 24498 19122 24510
rect 19070 24434 19122 24446
rect 28926 24498 28978 24510
rect 41358 24498 41410 24510
rect 36082 24446 36094 24498
rect 36146 24446 36158 24498
rect 28926 24434 28978 24446
rect 41358 24434 41410 24446
rect 54686 24498 54738 24510
rect 54686 24434 54738 24446
rect 1344 24330 78624 24364
rect 1344 24278 10874 24330
rect 10926 24278 10978 24330
rect 11030 24278 11082 24330
rect 11134 24278 30194 24330
rect 30246 24278 30298 24330
rect 30350 24278 30402 24330
rect 30454 24278 49514 24330
rect 49566 24278 49618 24330
rect 49670 24278 49722 24330
rect 49774 24278 68834 24330
rect 68886 24278 68938 24330
rect 68990 24278 69042 24330
rect 69094 24278 78624 24330
rect 1344 24244 78624 24278
rect 21422 24162 21474 24174
rect 21422 24098 21474 24110
rect 22094 24162 22146 24174
rect 22094 24098 22146 24110
rect 28366 24162 28418 24174
rect 28366 24098 28418 24110
rect 31502 24162 31554 24174
rect 31502 24098 31554 24110
rect 31838 24162 31890 24174
rect 31838 24098 31890 24110
rect 34302 24162 34354 24174
rect 34302 24098 34354 24110
rect 36318 24162 36370 24174
rect 61394 24110 61406 24162
rect 61458 24110 61470 24162
rect 36318 24098 36370 24110
rect 1934 24050 1986 24062
rect 1934 23986 1986 23998
rect 4846 24050 4898 24062
rect 21870 24050 21922 24062
rect 8642 23998 8654 24050
rect 8706 23998 8718 24050
rect 16258 23998 16270 24050
rect 16322 23998 16334 24050
rect 19842 23998 19854 24050
rect 19906 23998 19918 24050
rect 4846 23986 4898 23998
rect 21870 23986 21922 23998
rect 25230 24050 25282 24062
rect 25230 23986 25282 23998
rect 26014 24050 26066 24062
rect 26014 23986 26066 23998
rect 27470 24050 27522 24062
rect 44158 24050 44210 24062
rect 29810 23998 29822 24050
rect 29874 23998 29886 24050
rect 33842 23998 33854 24050
rect 33906 23998 33918 24050
rect 39778 23998 39790 24050
rect 39842 23998 39854 24050
rect 27470 23986 27522 23998
rect 44158 23986 44210 23998
rect 45390 24050 45442 24062
rect 45390 23986 45442 23998
rect 45950 24050 46002 24062
rect 45950 23986 46002 23998
rect 49422 24050 49474 24062
rect 49422 23986 49474 23998
rect 52222 24050 52274 24062
rect 52222 23986 52274 23998
rect 52894 24050 52946 24062
rect 52894 23986 52946 23998
rect 54126 24050 54178 24062
rect 54126 23986 54178 23998
rect 56254 24050 56306 24062
rect 56254 23986 56306 23998
rect 58718 24050 58770 24062
rect 64766 24050 64818 24062
rect 75406 24050 75458 24062
rect 61842 23998 61854 24050
rect 61906 23998 61918 24050
rect 72258 23998 72270 24050
rect 72322 23998 72334 24050
rect 58718 23986 58770 23998
rect 64766 23986 64818 23998
rect 75406 23986 75458 23998
rect 9438 23938 9490 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 5730 23886 5742 23938
rect 5794 23886 5806 23938
rect 9438 23874 9490 23886
rect 11678 23938 11730 23950
rect 11678 23874 11730 23886
rect 15262 23938 15314 23950
rect 21310 23938 21362 23950
rect 16706 23886 16718 23938
rect 16770 23886 16782 23938
rect 17490 23886 17502 23938
rect 17554 23886 17566 23938
rect 18498 23886 18510 23938
rect 18562 23886 18574 23938
rect 19058 23886 19070 23938
rect 19122 23886 19134 23938
rect 15262 23874 15314 23886
rect 21310 23874 21362 23886
rect 23438 23938 23490 23950
rect 35982 23938 36034 23950
rect 38110 23938 38162 23950
rect 29698 23886 29710 23938
rect 29762 23886 29774 23938
rect 32610 23886 32622 23938
rect 32674 23886 32686 23938
rect 33394 23886 33406 23938
rect 33458 23886 33470 23938
rect 34066 23886 34078 23938
rect 34130 23886 34142 23938
rect 35522 23886 35534 23938
rect 35586 23886 35598 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 23438 23874 23490 23886
rect 35982 23874 36034 23886
rect 38110 23874 38162 23886
rect 38222 23938 38274 23950
rect 42702 23938 42754 23950
rect 38434 23886 38446 23938
rect 38498 23886 38510 23938
rect 38770 23886 38782 23938
rect 38834 23886 38846 23938
rect 39442 23886 39454 23938
rect 39506 23886 39518 23938
rect 41682 23886 41694 23938
rect 41746 23886 41758 23938
rect 38222 23874 38274 23886
rect 42702 23874 42754 23886
rect 42926 23938 42978 23950
rect 42926 23874 42978 23886
rect 43710 23938 43762 23950
rect 57598 23938 57650 23950
rect 47842 23886 47854 23938
rect 47906 23886 47918 23938
rect 48738 23886 48750 23938
rect 48802 23886 48814 23938
rect 53218 23886 53230 23938
rect 53282 23886 53294 23938
rect 54450 23886 54462 23938
rect 54514 23886 54526 23938
rect 43710 23874 43762 23886
rect 57598 23874 57650 23886
rect 58830 23938 58882 23950
rect 70030 23938 70082 23950
rect 72158 23938 72210 23950
rect 61618 23886 61630 23938
rect 61682 23886 61694 23938
rect 62514 23886 62526 23938
rect 62578 23886 62590 23938
rect 70802 23886 70814 23938
rect 70866 23886 70878 23938
rect 71026 23886 71038 23938
rect 71090 23886 71102 23938
rect 72706 23886 72718 23938
rect 72770 23886 72782 23938
rect 73042 23886 73054 23938
rect 73106 23886 73118 23938
rect 58830 23874 58882 23886
rect 70030 23874 70082 23886
rect 72158 23874 72210 23886
rect 11342 23826 11394 23838
rect 6514 23774 6526 23826
rect 6578 23774 6590 23826
rect 9650 23774 9662 23826
rect 9714 23774 9726 23826
rect 9986 23774 9998 23826
rect 10050 23774 10062 23826
rect 11342 23762 11394 23774
rect 22766 23826 22818 23838
rect 22766 23762 22818 23774
rect 22990 23826 23042 23838
rect 28254 23826 28306 23838
rect 30606 23826 30658 23838
rect 26338 23774 26350 23826
rect 26402 23774 26414 23826
rect 29474 23774 29486 23826
rect 29538 23774 29550 23826
rect 22990 23762 23042 23774
rect 28254 23762 28306 23774
rect 30606 23762 30658 23774
rect 31054 23826 31106 23838
rect 41470 23826 41522 23838
rect 32386 23774 32398 23826
rect 32450 23774 32462 23826
rect 35298 23774 35310 23826
rect 35362 23774 35374 23826
rect 31054 23762 31106 23774
rect 41470 23762 41522 23774
rect 43262 23826 43314 23838
rect 43262 23762 43314 23774
rect 43598 23826 43650 23838
rect 55022 23826 55074 23838
rect 47506 23774 47518 23826
rect 47570 23774 47582 23826
rect 43598 23762 43650 23774
rect 55022 23762 55074 23774
rect 57374 23826 57426 23838
rect 57374 23762 57426 23774
rect 59054 23826 59106 23838
rect 59054 23762 59106 23774
rect 59390 23826 59442 23838
rect 59390 23762 59442 23774
rect 59502 23826 59554 23838
rect 59502 23762 59554 23774
rect 66446 23826 66498 23838
rect 72270 23826 72322 23838
rect 69570 23774 69582 23826
rect 69634 23774 69646 23826
rect 71586 23774 71598 23826
rect 71650 23774 71662 23826
rect 66446 23762 66498 23774
rect 72270 23762 72322 23774
rect 9102 23714 9154 23726
rect 9102 23650 9154 23662
rect 13582 23714 13634 23726
rect 13582 23650 13634 23662
rect 21422 23714 21474 23726
rect 23102 23714 23154 23726
rect 22418 23662 22430 23714
rect 22482 23662 22494 23714
rect 21422 23650 21474 23662
rect 23102 23650 23154 23662
rect 23774 23714 23826 23726
rect 23774 23650 23826 23662
rect 25790 23714 25842 23726
rect 27022 23714 27074 23726
rect 26674 23662 26686 23714
rect 26738 23662 26750 23714
rect 25790 23650 25842 23662
rect 27022 23650 27074 23662
rect 28030 23714 28082 23726
rect 28030 23650 28082 23662
rect 28366 23714 28418 23726
rect 28366 23650 28418 23662
rect 37102 23714 37154 23726
rect 37102 23650 37154 23662
rect 43038 23714 43090 23726
rect 43038 23650 43090 23662
rect 50766 23714 50818 23726
rect 50766 23650 50818 23662
rect 53566 23714 53618 23726
rect 53566 23650 53618 23662
rect 54574 23714 54626 23726
rect 54574 23650 54626 23662
rect 57710 23714 57762 23726
rect 57710 23650 57762 23662
rect 57822 23714 57874 23726
rect 57822 23650 57874 23662
rect 57934 23714 57986 23726
rect 57934 23650 57986 23662
rect 58494 23714 58546 23726
rect 58494 23650 58546 23662
rect 58606 23714 58658 23726
rect 58606 23650 58658 23662
rect 59726 23714 59778 23726
rect 59726 23650 59778 23662
rect 60622 23714 60674 23726
rect 60622 23650 60674 23662
rect 64206 23714 64258 23726
rect 64206 23650 64258 23662
rect 66782 23714 66834 23726
rect 66782 23650 66834 23662
rect 69246 23714 69298 23726
rect 72494 23714 72546 23726
rect 69906 23662 69918 23714
rect 69970 23662 69982 23714
rect 69246 23650 69298 23662
rect 72494 23650 72546 23662
rect 76526 23714 76578 23726
rect 76526 23650 76578 23662
rect 1344 23546 78784 23580
rect 1344 23494 20534 23546
rect 20586 23494 20638 23546
rect 20690 23494 20742 23546
rect 20794 23494 39854 23546
rect 39906 23494 39958 23546
rect 40010 23494 40062 23546
rect 40114 23494 59174 23546
rect 59226 23494 59278 23546
rect 59330 23494 59382 23546
rect 59434 23494 78494 23546
rect 78546 23494 78598 23546
rect 78650 23494 78702 23546
rect 78754 23494 78784 23546
rect 1344 23460 78784 23494
rect 6862 23378 6914 23390
rect 6862 23314 6914 23326
rect 8654 23378 8706 23390
rect 8654 23314 8706 23326
rect 15710 23378 15762 23390
rect 15710 23314 15762 23326
rect 16270 23378 16322 23390
rect 19630 23378 19682 23390
rect 18162 23326 18174 23378
rect 18226 23326 18238 23378
rect 16270 23314 16322 23326
rect 19630 23314 19682 23326
rect 22206 23378 22258 23390
rect 22206 23314 22258 23326
rect 22430 23378 22482 23390
rect 22430 23314 22482 23326
rect 22878 23378 22930 23390
rect 22878 23314 22930 23326
rect 23438 23378 23490 23390
rect 23438 23314 23490 23326
rect 24558 23378 24610 23390
rect 27246 23378 27298 23390
rect 25330 23326 25342 23378
rect 25394 23326 25406 23378
rect 24558 23314 24610 23326
rect 27246 23314 27298 23326
rect 30494 23378 30546 23390
rect 33518 23378 33570 23390
rect 31602 23326 31614 23378
rect 31666 23326 31678 23378
rect 30494 23314 30546 23326
rect 33518 23314 33570 23326
rect 33742 23378 33794 23390
rect 33742 23314 33794 23326
rect 36094 23378 36146 23390
rect 41470 23378 41522 23390
rect 40226 23326 40238 23378
rect 40290 23326 40302 23378
rect 36094 23314 36146 23326
rect 41470 23314 41522 23326
rect 42814 23378 42866 23390
rect 42814 23314 42866 23326
rect 46174 23378 46226 23390
rect 47518 23378 47570 23390
rect 47170 23326 47182 23378
rect 47234 23326 47246 23378
rect 46174 23314 46226 23326
rect 47518 23314 47570 23326
rect 50094 23378 50146 23390
rect 51662 23378 51714 23390
rect 52782 23378 52834 23390
rect 51314 23326 51326 23378
rect 51378 23326 51390 23378
rect 51986 23326 51998 23378
rect 52050 23326 52062 23378
rect 50094 23314 50146 23326
rect 51662 23314 51714 23326
rect 52782 23314 52834 23326
rect 53118 23378 53170 23390
rect 53118 23314 53170 23326
rect 60398 23378 60450 23390
rect 60398 23314 60450 23326
rect 60622 23378 60674 23390
rect 60622 23314 60674 23326
rect 61742 23378 61794 23390
rect 61742 23314 61794 23326
rect 62974 23378 63026 23390
rect 62974 23314 63026 23326
rect 65102 23378 65154 23390
rect 65102 23314 65154 23326
rect 65662 23378 65714 23390
rect 70354 23326 70366 23378
rect 70418 23326 70430 23378
rect 65662 23314 65714 23326
rect 7198 23266 7250 23278
rect 7198 23202 7250 23214
rect 15486 23266 15538 23278
rect 15486 23202 15538 23214
rect 16046 23266 16098 23278
rect 21982 23266 22034 23278
rect 19058 23214 19070 23266
rect 19122 23214 19134 23266
rect 16046 23202 16098 23214
rect 21982 23202 22034 23214
rect 22766 23266 22818 23278
rect 30382 23266 30434 23278
rect 26226 23214 26238 23266
rect 26290 23214 26302 23266
rect 28354 23214 28366 23266
rect 28418 23214 28430 23266
rect 22766 23202 22818 23214
rect 30382 23202 30434 23214
rect 36654 23266 36706 23278
rect 42366 23266 42418 23278
rect 39666 23214 39678 23266
rect 39730 23214 39742 23266
rect 36654 23202 36706 23214
rect 42366 23202 42418 23214
rect 53006 23266 53058 23278
rect 53006 23202 53058 23214
rect 55470 23266 55522 23278
rect 55470 23202 55522 23214
rect 57150 23266 57202 23278
rect 61182 23266 61234 23278
rect 59714 23214 59726 23266
rect 59778 23214 59790 23266
rect 57150 23202 57202 23214
rect 61182 23202 61234 23214
rect 63198 23266 63250 23278
rect 66770 23214 66782 23266
rect 66834 23214 66846 23266
rect 71362 23214 71374 23266
rect 71426 23214 71438 23266
rect 73154 23214 73166 23266
rect 73218 23214 73230 23266
rect 76962 23214 76974 23266
rect 77026 23214 77038 23266
rect 63198 23202 63250 23214
rect 15374 23154 15426 23166
rect 1810 23102 1822 23154
rect 1874 23102 1886 23154
rect 15374 23090 15426 23102
rect 15934 23154 15986 23166
rect 31054 23154 31106 23166
rect 18050 23102 18062 23154
rect 18114 23102 18126 23154
rect 18722 23102 18734 23154
rect 18786 23102 18798 23154
rect 25666 23102 25678 23154
rect 25730 23102 25742 23154
rect 26674 23102 26686 23154
rect 26738 23102 26750 23154
rect 27458 23102 27470 23154
rect 27522 23102 27534 23154
rect 29586 23102 29598 23154
rect 29650 23102 29662 23154
rect 30706 23102 30718 23154
rect 30770 23102 30782 23154
rect 15934 23090 15986 23102
rect 31054 23090 31106 23102
rect 31278 23154 31330 23166
rect 32510 23154 32562 23166
rect 32050 23102 32062 23154
rect 32114 23102 32126 23154
rect 31278 23090 31330 23102
rect 32510 23090 32562 23102
rect 34190 23154 34242 23166
rect 34190 23090 34242 23102
rect 34638 23154 34690 23166
rect 34638 23090 34690 23102
rect 35534 23154 35586 23166
rect 35534 23090 35586 23102
rect 36542 23154 36594 23166
rect 41246 23154 41298 23166
rect 37202 23102 37214 23154
rect 37266 23102 37278 23154
rect 39778 23102 39790 23154
rect 39842 23102 39854 23154
rect 40114 23102 40126 23154
rect 40178 23102 40190 23154
rect 40898 23102 40910 23154
rect 40962 23102 40974 23154
rect 36542 23090 36594 23102
rect 41246 23090 41298 23102
rect 42702 23154 42754 23166
rect 42702 23090 42754 23102
rect 43038 23154 43090 23166
rect 50654 23154 50706 23166
rect 45938 23102 45950 23154
rect 46002 23102 46014 23154
rect 43038 23090 43090 23102
rect 50654 23090 50706 23102
rect 50990 23154 51042 23166
rect 50990 23090 51042 23102
rect 54238 23154 54290 23166
rect 58382 23154 58434 23166
rect 60734 23154 60786 23166
rect 56018 23102 56030 23154
rect 56082 23102 56094 23154
rect 58146 23102 58158 23154
rect 58210 23102 58222 23154
rect 59490 23102 59502 23154
rect 59554 23102 59566 23154
rect 54238 23090 54290 23102
rect 58382 23090 58434 23102
rect 60734 23090 60786 23102
rect 60958 23154 61010 23166
rect 60958 23090 61010 23102
rect 61294 23154 61346 23166
rect 61294 23090 61346 23102
rect 62638 23154 62690 23166
rect 62638 23090 62690 23102
rect 63310 23154 63362 23166
rect 72830 23154 72882 23166
rect 65986 23102 65998 23154
rect 66050 23102 66062 23154
rect 70578 23102 70590 23154
rect 70642 23102 70654 23154
rect 71138 23102 71150 23154
rect 71202 23102 71214 23154
rect 73602 23102 73614 23154
rect 73666 23102 73678 23154
rect 76850 23102 76862 23154
rect 76914 23102 76926 23154
rect 63310 23090 63362 23102
rect 72830 23090 72882 23102
rect 15038 23042 15090 23054
rect 2482 22990 2494 23042
rect 2546 22990 2558 23042
rect 4610 22990 4622 23042
rect 4674 22990 4686 23042
rect 15038 22978 15090 22990
rect 16606 23042 16658 23054
rect 16606 22978 16658 22990
rect 22094 23042 22146 23054
rect 35310 23042 35362 23054
rect 39006 23042 39058 23054
rect 24098 22990 24110 23042
rect 24162 22990 24174 23042
rect 26002 22990 26014 23042
rect 26066 22990 26078 23042
rect 29138 22990 29150 23042
rect 29202 22990 29214 23042
rect 38210 22990 38222 23042
rect 38274 22990 38286 23042
rect 22094 22978 22146 22990
rect 35310 22978 35362 22990
rect 39006 22978 39058 22990
rect 41358 23042 41410 23054
rect 41358 22978 41410 22990
rect 41918 23042 41970 23054
rect 41918 22978 41970 22990
rect 43374 23042 43426 23054
rect 43374 22978 43426 22990
rect 43822 23042 43874 23054
rect 43822 22978 43874 22990
rect 44606 23042 44658 23054
rect 44606 22978 44658 22990
rect 45054 23042 45106 23054
rect 45054 22978 45106 22990
rect 45502 23042 45554 23054
rect 45502 22978 45554 22990
rect 46734 23042 46786 23054
rect 46734 22978 46786 22990
rect 49422 23042 49474 23054
rect 49422 22978 49474 22990
rect 54126 23042 54178 23054
rect 54126 22978 54178 22990
rect 58494 23042 58546 23054
rect 62190 23042 62242 23054
rect 72494 23042 72546 23054
rect 60162 22990 60174 23042
rect 60226 22990 60238 23042
rect 68898 22990 68910 23042
rect 68962 22990 68974 23042
rect 71474 22990 71486 23042
rect 71538 22990 71550 23042
rect 74274 22990 74286 23042
rect 74338 22990 74350 23042
rect 76402 22990 76414 23042
rect 76466 22990 76478 23042
rect 58494 22978 58546 22990
rect 62190 22978 62242 22990
rect 72494 22978 72546 22990
rect 34414 22930 34466 22942
rect 77646 22930 77698 22942
rect 64866 22878 64878 22930
rect 64930 22927 64942 22930
rect 65090 22927 65102 22930
rect 64930 22881 65102 22927
rect 64930 22878 64942 22881
rect 65090 22878 65102 22881
rect 65154 22878 65166 22930
rect 34414 22866 34466 22878
rect 77646 22866 77698 22878
rect 77982 22930 78034 22942
rect 77982 22866 78034 22878
rect 1344 22762 78624 22796
rect 1344 22710 10874 22762
rect 10926 22710 10978 22762
rect 11030 22710 11082 22762
rect 11134 22710 30194 22762
rect 30246 22710 30298 22762
rect 30350 22710 30402 22762
rect 30454 22710 49514 22762
rect 49566 22710 49618 22762
rect 49670 22710 49722 22762
rect 49774 22710 68834 22762
rect 68886 22710 68938 22762
rect 68990 22710 69042 22762
rect 69094 22710 78624 22762
rect 1344 22676 78624 22710
rect 22206 22594 22258 22606
rect 40462 22594 40514 22606
rect 26338 22542 26350 22594
rect 26402 22542 26414 22594
rect 22206 22530 22258 22542
rect 40462 22530 40514 22542
rect 51326 22594 51378 22606
rect 66446 22594 66498 22606
rect 62290 22542 62302 22594
rect 62354 22542 62366 22594
rect 51326 22530 51378 22542
rect 66446 22530 66498 22542
rect 66782 22594 66834 22606
rect 66782 22530 66834 22542
rect 68350 22594 68402 22606
rect 68350 22530 68402 22542
rect 76638 22594 76690 22606
rect 76638 22530 76690 22542
rect 2046 22482 2098 22494
rect 2046 22418 2098 22430
rect 5742 22482 5794 22494
rect 5742 22418 5794 22430
rect 19406 22482 19458 22494
rect 19406 22418 19458 22430
rect 19854 22482 19906 22494
rect 19854 22418 19906 22430
rect 20302 22482 20354 22494
rect 20302 22418 20354 22430
rect 30830 22482 30882 22494
rect 51102 22482 51154 22494
rect 35746 22430 35758 22482
rect 35810 22430 35822 22482
rect 37202 22430 37214 22482
rect 37266 22430 37278 22482
rect 39778 22430 39790 22482
rect 39842 22430 39854 22482
rect 44930 22430 44942 22482
rect 44994 22430 45006 22482
rect 46610 22430 46622 22482
rect 46674 22430 46686 22482
rect 50194 22430 50206 22482
rect 50258 22430 50270 22482
rect 30830 22418 30882 22430
rect 51102 22418 51154 22430
rect 56142 22482 56194 22494
rect 56142 22418 56194 22430
rect 58046 22482 58098 22494
rect 58046 22418 58098 22430
rect 65774 22482 65826 22494
rect 75630 22482 75682 22494
rect 69346 22430 69358 22482
rect 69410 22430 69422 22482
rect 65774 22418 65826 22430
rect 75630 22418 75682 22430
rect 4174 22370 4226 22382
rect 18174 22370 18226 22382
rect 4946 22318 4958 22370
rect 5010 22318 5022 22370
rect 17266 22318 17278 22370
rect 17330 22318 17342 22370
rect 4174 22306 4226 22318
rect 18174 22306 18226 22318
rect 18286 22370 18338 22382
rect 18286 22306 18338 22318
rect 18510 22370 18562 22382
rect 22094 22370 22146 22382
rect 26462 22370 26514 22382
rect 18722 22318 18734 22370
rect 18786 22318 18798 22370
rect 23986 22318 23998 22370
rect 24050 22318 24062 22370
rect 24434 22318 24446 22370
rect 24498 22318 24510 22370
rect 24994 22318 25006 22370
rect 25058 22318 25070 22370
rect 18510 22306 18562 22318
rect 22094 22306 22146 22318
rect 26462 22306 26514 22318
rect 26574 22370 26626 22382
rect 28702 22370 28754 22382
rect 27458 22318 27470 22370
rect 27522 22318 27534 22370
rect 27906 22318 27918 22370
rect 27970 22318 27982 22370
rect 28242 22318 28254 22370
rect 28306 22318 28318 22370
rect 26574 22306 26626 22318
rect 28702 22306 28754 22318
rect 29150 22370 29202 22382
rect 29150 22306 29202 22318
rect 29598 22370 29650 22382
rect 42478 22370 42530 22382
rect 31378 22318 31390 22370
rect 31442 22318 31454 22370
rect 32162 22318 32174 22370
rect 32226 22318 32238 22370
rect 32722 22318 32734 22370
rect 32786 22318 32798 22370
rect 33618 22318 33630 22370
rect 33682 22318 33694 22370
rect 35410 22318 35422 22370
rect 35474 22318 35486 22370
rect 36194 22318 36206 22370
rect 36258 22318 36270 22370
rect 37090 22318 37102 22370
rect 37154 22318 37166 22370
rect 39330 22318 39342 22370
rect 39394 22318 39406 22370
rect 39890 22318 39902 22370
rect 39954 22318 39966 22370
rect 41010 22318 41022 22370
rect 41074 22318 41086 22370
rect 42130 22318 42142 22370
rect 42194 22318 42206 22370
rect 29598 22306 29650 22318
rect 42478 22306 42530 22318
rect 43262 22370 43314 22382
rect 43262 22306 43314 22318
rect 44270 22370 44322 22382
rect 44270 22306 44322 22318
rect 45054 22370 45106 22382
rect 45054 22306 45106 22318
rect 45278 22370 45330 22382
rect 46174 22370 46226 22382
rect 65326 22370 65378 22382
rect 45490 22318 45502 22370
rect 45554 22318 45566 22370
rect 47058 22318 47070 22370
rect 47122 22318 47134 22370
rect 48178 22318 48190 22370
rect 48242 22318 48254 22370
rect 48962 22318 48974 22370
rect 49026 22318 49038 22370
rect 54338 22318 54350 22370
rect 54402 22318 54414 22370
rect 58258 22318 58270 22370
rect 58322 22318 58334 22370
rect 60498 22318 60510 22370
rect 60562 22318 60574 22370
rect 61842 22318 61854 22370
rect 61906 22318 61918 22370
rect 63074 22318 63086 22370
rect 63138 22318 63150 22370
rect 65090 22318 65102 22370
rect 65154 22318 65166 22370
rect 45278 22306 45330 22318
rect 46174 22306 46226 22318
rect 65326 22306 65378 22318
rect 69022 22370 69074 22382
rect 69022 22306 69074 22318
rect 69694 22370 69746 22382
rect 70354 22318 70366 22370
rect 70418 22318 70430 22370
rect 72258 22318 72270 22370
rect 72322 22318 72334 22370
rect 74834 22318 74846 22370
rect 74898 22318 74910 22370
rect 78082 22318 78094 22370
rect 78146 22318 78158 22370
rect 69694 22306 69746 22318
rect 2830 22258 2882 22270
rect 2830 22194 2882 22206
rect 3166 22258 3218 22270
rect 3166 22194 3218 22206
rect 3838 22258 3890 22270
rect 16270 22258 16322 22270
rect 4722 22206 4734 22258
rect 4786 22206 4798 22258
rect 3838 22194 3890 22206
rect 16270 22194 16322 22206
rect 16606 22258 16658 22270
rect 25678 22258 25730 22270
rect 24546 22206 24558 22258
rect 24610 22206 24622 22258
rect 16606 22194 16658 22206
rect 25678 22194 25730 22206
rect 29934 22258 29986 22270
rect 29934 22194 29986 22206
rect 30606 22258 30658 22270
rect 30606 22194 30658 22206
rect 31166 22258 31218 22270
rect 40350 22258 40402 22270
rect 54910 22258 54962 22270
rect 32274 22206 32286 22258
rect 32338 22206 32350 22258
rect 34626 22206 34638 22258
rect 34690 22206 34702 22258
rect 36418 22206 36430 22258
rect 36482 22206 36494 22258
rect 36978 22206 36990 22258
rect 37042 22206 37054 22258
rect 41682 22206 41694 22258
rect 41746 22206 41758 22258
rect 42802 22206 42814 22258
rect 42866 22206 42878 22258
rect 31166 22194 31218 22206
rect 40350 22194 40402 22206
rect 54910 22194 54962 22206
rect 59278 22258 59330 22270
rect 68462 22258 68514 22270
rect 60834 22206 60846 22258
rect 60898 22206 60910 22258
rect 66994 22206 67006 22258
rect 67058 22206 67070 22258
rect 67442 22206 67454 22258
rect 67506 22206 67518 22258
rect 59278 22194 59330 22206
rect 68462 22194 68514 22206
rect 69358 22258 69410 22270
rect 69358 22194 69410 22206
rect 69918 22258 69970 22270
rect 71586 22262 71598 22314
rect 71650 22262 71662 22314
rect 74174 22258 74226 22270
rect 73378 22206 73390 22258
rect 73442 22206 73454 22258
rect 76850 22206 76862 22258
rect 76914 22206 76926 22258
rect 77186 22206 77198 22258
rect 77250 22206 77262 22258
rect 69918 22194 69970 22206
rect 74174 22194 74226 22206
rect 12238 22146 12290 22158
rect 11890 22094 11902 22146
rect 11954 22094 11966 22146
rect 12238 22082 12290 22094
rect 12686 22146 12738 22158
rect 13806 22146 13858 22158
rect 13458 22094 13470 22146
rect 13522 22094 13534 22146
rect 12686 22082 12738 22094
rect 13806 22082 13858 22094
rect 14254 22146 14306 22158
rect 14254 22082 14306 22094
rect 16830 22146 16882 22158
rect 16830 22082 16882 22094
rect 16942 22146 16994 22158
rect 16942 22082 16994 22094
rect 17054 22146 17106 22158
rect 17054 22082 17106 22094
rect 18398 22146 18450 22158
rect 18398 22082 18450 22094
rect 22206 22146 22258 22158
rect 22206 22082 22258 22094
rect 22878 22146 22930 22158
rect 22878 22082 22930 22094
rect 23550 22146 23602 22158
rect 23550 22082 23602 22094
rect 25790 22146 25842 22158
rect 25790 22082 25842 22094
rect 26014 22146 26066 22158
rect 26014 22082 26066 22094
rect 30718 22146 30770 22158
rect 30718 22082 30770 22094
rect 30942 22146 30994 22158
rect 43710 22146 43762 22158
rect 41122 22094 41134 22146
rect 41186 22094 41198 22146
rect 30942 22082 30994 22094
rect 43710 22082 43762 22094
rect 44942 22146 44994 22158
rect 44942 22082 44994 22094
rect 47182 22146 47234 22158
rect 47182 22082 47234 22094
rect 49758 22146 49810 22158
rect 49758 22082 49810 22094
rect 50878 22146 50930 22158
rect 52222 22146 52274 22158
rect 51650 22094 51662 22146
rect 51714 22094 51726 22146
rect 50878 22082 50930 22094
rect 52222 22082 52274 22094
rect 54462 22146 54514 22158
rect 54462 22082 54514 22094
rect 57486 22146 57538 22158
rect 68686 22146 68738 22158
rect 61058 22094 61070 22146
rect 61122 22094 61134 22146
rect 57486 22082 57538 22094
rect 68686 22082 68738 22094
rect 69470 22146 69522 22158
rect 76302 22146 76354 22158
rect 75058 22094 75070 22146
rect 75122 22094 75134 22146
rect 69470 22082 69522 22094
rect 76302 22082 76354 22094
rect 77870 22146 77922 22158
rect 77870 22082 77922 22094
rect 1344 21978 78784 22012
rect 1344 21926 20534 21978
rect 20586 21926 20638 21978
rect 20690 21926 20742 21978
rect 20794 21926 39854 21978
rect 39906 21926 39958 21978
rect 40010 21926 40062 21978
rect 40114 21926 59174 21978
rect 59226 21926 59278 21978
rect 59330 21926 59382 21978
rect 59434 21926 78494 21978
rect 78546 21926 78598 21978
rect 78650 21926 78702 21978
rect 78754 21926 78784 21978
rect 1344 21892 78784 21926
rect 2158 21810 2210 21822
rect 2158 21746 2210 21758
rect 12686 21810 12738 21822
rect 14142 21810 14194 21822
rect 16606 21810 16658 21822
rect 13458 21758 13470 21810
rect 13522 21758 13534 21810
rect 14466 21758 14478 21810
rect 14530 21758 14542 21810
rect 15138 21758 15150 21810
rect 15202 21758 15214 21810
rect 12686 21746 12738 21758
rect 14142 21746 14194 21758
rect 16606 21746 16658 21758
rect 18510 21810 18562 21822
rect 22990 21810 23042 21822
rect 19954 21758 19966 21810
rect 20018 21758 20030 21810
rect 18510 21746 18562 21758
rect 22990 21746 23042 21758
rect 23998 21810 24050 21822
rect 23998 21746 24050 21758
rect 24110 21810 24162 21822
rect 24110 21746 24162 21758
rect 27806 21810 27858 21822
rect 27806 21746 27858 21758
rect 29598 21810 29650 21822
rect 29598 21746 29650 21758
rect 29934 21810 29986 21822
rect 31950 21810 32002 21822
rect 31042 21758 31054 21810
rect 31106 21758 31118 21810
rect 29934 21746 29986 21758
rect 31950 21746 32002 21758
rect 38782 21810 38834 21822
rect 38782 21746 38834 21758
rect 41022 21810 41074 21822
rect 41022 21746 41074 21758
rect 41918 21810 41970 21822
rect 41918 21746 41970 21758
rect 42366 21810 42418 21822
rect 42366 21746 42418 21758
rect 46622 21810 46674 21822
rect 46622 21746 46674 21758
rect 47966 21810 48018 21822
rect 47966 21746 48018 21758
rect 50318 21810 50370 21822
rect 50318 21746 50370 21758
rect 50878 21810 50930 21822
rect 50878 21746 50930 21758
rect 51214 21810 51266 21822
rect 51214 21746 51266 21758
rect 51998 21810 52050 21822
rect 51998 21746 52050 21758
rect 52334 21810 52386 21822
rect 52334 21746 52386 21758
rect 59726 21810 59778 21822
rect 59726 21746 59778 21758
rect 59838 21810 59890 21822
rect 59838 21746 59890 21758
rect 60062 21810 60114 21822
rect 60062 21746 60114 21758
rect 64542 21810 64594 21822
rect 66894 21810 66946 21822
rect 65314 21758 65326 21810
rect 65378 21758 65390 21810
rect 64542 21746 64594 21758
rect 66894 21746 66946 21758
rect 72606 21810 72658 21822
rect 72606 21746 72658 21758
rect 72718 21810 72770 21822
rect 72718 21746 72770 21758
rect 73502 21810 73554 21822
rect 73502 21746 73554 21758
rect 74062 21810 74114 21822
rect 74062 21746 74114 21758
rect 74398 21810 74450 21822
rect 74398 21746 74450 21758
rect 1710 21698 1762 21710
rect 1710 21634 1762 21646
rect 15598 21698 15650 21710
rect 15598 21634 15650 21646
rect 18734 21698 18786 21710
rect 18734 21634 18786 21646
rect 19518 21698 19570 21710
rect 24334 21698 24386 21710
rect 20290 21646 20302 21698
rect 20354 21646 20366 21698
rect 19518 21634 19570 21646
rect 24334 21634 24386 21646
rect 26686 21698 26738 21710
rect 26686 21634 26738 21646
rect 29822 21698 29874 21710
rect 38446 21698 38498 21710
rect 36978 21646 36990 21698
rect 37042 21646 37054 21698
rect 29822 21634 29874 21646
rect 38446 21634 38498 21646
rect 39230 21698 39282 21710
rect 39230 21634 39282 21646
rect 51774 21698 51826 21710
rect 51774 21634 51826 21646
rect 57598 21698 57650 21710
rect 57598 21634 57650 21646
rect 59502 21698 59554 21710
rect 59502 21634 59554 21646
rect 64878 21698 64930 21710
rect 67118 21698 67170 21710
rect 65538 21646 65550 21698
rect 65602 21646 65614 21698
rect 66210 21646 66222 21698
rect 66274 21646 66286 21698
rect 64878 21634 64930 21646
rect 67118 21634 67170 21646
rect 67678 21698 67730 21710
rect 67678 21634 67730 21646
rect 70478 21698 70530 21710
rect 73726 21698 73778 21710
rect 71698 21646 71710 21698
rect 71762 21646 71774 21698
rect 70478 21634 70530 21646
rect 73726 21634 73778 21646
rect 74734 21698 74786 21710
rect 75842 21646 75854 21698
rect 75906 21646 75918 21698
rect 74734 21634 74786 21646
rect 10558 21586 10610 21598
rect 2370 21534 2382 21586
rect 2434 21534 2446 21586
rect 2818 21534 2830 21586
rect 2882 21534 2894 21586
rect 6178 21534 6190 21586
rect 6242 21534 6254 21586
rect 10322 21534 10334 21586
rect 10386 21534 10398 21586
rect 10558 21522 10610 21534
rect 10670 21586 10722 21598
rect 11566 21586 11618 21598
rect 15710 21586 15762 21598
rect 18286 21586 18338 21598
rect 11106 21534 11118 21586
rect 11170 21534 11182 21586
rect 13682 21534 13694 21586
rect 13746 21534 13758 21586
rect 15922 21534 15934 21586
rect 15986 21534 15998 21586
rect 10670 21522 10722 21534
rect 11566 21522 11618 21534
rect 15710 21522 15762 21534
rect 18286 21522 18338 21534
rect 18398 21586 18450 21598
rect 18398 21522 18450 21534
rect 18622 21586 18674 21598
rect 18622 21522 18674 21534
rect 19294 21586 19346 21598
rect 19294 21522 19346 21534
rect 19406 21586 19458 21598
rect 19406 21522 19458 21534
rect 20638 21586 20690 21598
rect 20638 21522 20690 21534
rect 23438 21586 23490 21598
rect 23438 21522 23490 21534
rect 23774 21586 23826 21598
rect 23774 21522 23826 21534
rect 23886 21586 23938 21598
rect 23886 21522 23938 21534
rect 26126 21586 26178 21598
rect 26126 21522 26178 21534
rect 26462 21586 26514 21598
rect 26462 21522 26514 21534
rect 27470 21586 27522 21598
rect 27470 21522 27522 21534
rect 27918 21586 27970 21598
rect 27918 21522 27970 21534
rect 29038 21586 29090 21598
rect 29038 21522 29090 21534
rect 29262 21586 29314 21598
rect 31390 21586 31442 21598
rect 38670 21586 38722 21598
rect 30370 21534 30382 21586
rect 30434 21534 30446 21586
rect 34738 21534 34750 21586
rect 34802 21534 34814 21586
rect 35970 21534 35982 21586
rect 36034 21534 36046 21586
rect 36418 21534 36430 21586
rect 36482 21534 36494 21586
rect 29262 21522 29314 21534
rect 31390 21522 31442 21534
rect 38670 21522 38722 21534
rect 38894 21586 38946 21598
rect 42814 21586 42866 21598
rect 47742 21586 47794 21598
rect 40114 21534 40126 21586
rect 40178 21534 40190 21586
rect 43362 21534 43374 21586
rect 43426 21534 43438 21586
rect 43586 21534 43598 21586
rect 43650 21534 43662 21586
rect 44706 21534 44718 21586
rect 44770 21534 44782 21586
rect 45154 21534 45166 21586
rect 45218 21534 45230 21586
rect 45602 21534 45614 21586
rect 45666 21534 45678 21586
rect 47506 21534 47518 21586
rect 47570 21534 47582 21586
rect 38894 21522 38946 21534
rect 42814 21522 42866 21534
rect 47742 21522 47794 21534
rect 48078 21586 48130 21598
rect 48078 21522 48130 21534
rect 48862 21586 48914 21598
rect 48862 21522 48914 21534
rect 49310 21586 49362 21598
rect 49310 21522 49362 21534
rect 49870 21586 49922 21598
rect 49870 21522 49922 21534
rect 50990 21586 51042 21598
rect 50990 21522 51042 21534
rect 51326 21586 51378 21598
rect 51326 21522 51378 21534
rect 52222 21586 52274 21598
rect 58382 21586 58434 21598
rect 58146 21534 58158 21586
rect 58210 21534 58222 21586
rect 52222 21522 52274 21534
rect 58382 21522 58434 21534
rect 59950 21586 60002 21598
rect 65326 21586 65378 21598
rect 63858 21534 63870 21586
rect 63922 21534 63934 21586
rect 59950 21522 60002 21534
rect 65326 21522 65378 21534
rect 67230 21586 67282 21598
rect 72494 21586 72546 21598
rect 70802 21534 70814 21586
rect 70866 21534 70878 21586
rect 71250 21534 71262 21586
rect 71314 21534 71326 21586
rect 72258 21534 72270 21586
rect 72322 21534 72334 21586
rect 72930 21534 72942 21586
rect 72994 21534 73006 21586
rect 75170 21534 75182 21586
rect 75234 21534 75246 21586
rect 67230 21522 67282 21534
rect 72494 21522 72546 21534
rect 11342 21474 11394 21486
rect 3602 21422 3614 21474
rect 3666 21422 3678 21474
rect 5730 21422 5742 21474
rect 5794 21422 5806 21474
rect 6850 21422 6862 21474
rect 6914 21422 6926 21474
rect 8978 21422 8990 21474
rect 9042 21422 9054 21474
rect 11342 21410 11394 21422
rect 11454 21474 11506 21486
rect 11454 21410 11506 21422
rect 12350 21474 12402 21486
rect 12350 21410 12402 21422
rect 13246 21474 13298 21486
rect 13246 21410 13298 21422
rect 17838 21474 17890 21486
rect 17838 21410 17890 21422
rect 21086 21474 21138 21486
rect 21086 21410 21138 21422
rect 22094 21474 22146 21486
rect 22094 21410 22146 21422
rect 22430 21474 22482 21486
rect 22430 21410 22482 21422
rect 25566 21474 25618 21486
rect 32286 21474 32338 21486
rect 28578 21422 28590 21474
rect 28642 21422 28654 21474
rect 30258 21422 30270 21474
rect 30322 21422 30334 21474
rect 25566 21410 25618 21422
rect 32286 21410 32338 21422
rect 33182 21474 33234 21486
rect 41470 21474 41522 21486
rect 47182 21474 47234 21486
rect 34290 21422 34302 21474
rect 34354 21422 34366 21474
rect 36866 21422 36878 21474
rect 36930 21422 36942 21474
rect 39666 21422 39678 21474
rect 39730 21422 39742 21474
rect 45490 21422 45502 21474
rect 45554 21422 45566 21474
rect 33182 21410 33234 21422
rect 41470 21410 41522 21422
rect 47182 21410 47234 21422
rect 47854 21474 47906 21486
rect 58494 21474 58546 21486
rect 50866 21422 50878 21474
rect 50930 21422 50942 21474
rect 52322 21422 52334 21474
rect 52386 21422 52398 21474
rect 47854 21410 47906 21422
rect 58494 21410 58546 21422
rect 60622 21474 60674 21486
rect 77982 21474 78034 21486
rect 60946 21422 60958 21474
rect 61010 21422 61022 21474
rect 63074 21422 63086 21474
rect 63138 21422 63150 21474
rect 71362 21422 71374 21474
rect 71426 21422 71438 21474
rect 60622 21410 60674 21422
rect 77982 21410 78034 21422
rect 1822 21362 1874 21374
rect 44158 21362 44210 21374
rect 21858 21310 21870 21362
rect 21922 21359 21934 21362
rect 22530 21359 22542 21362
rect 21922 21313 22542 21359
rect 21922 21310 21934 21313
rect 22530 21310 22542 21313
rect 22594 21359 22606 21362
rect 22978 21359 22990 21362
rect 22594 21313 22990 21359
rect 22594 21310 22606 21313
rect 22978 21310 22990 21313
rect 23042 21310 23054 21362
rect 41458 21310 41470 21362
rect 41522 21359 41534 21362
rect 41682 21359 41694 21362
rect 41522 21313 41694 21359
rect 41522 21310 41534 21313
rect 41682 21310 41694 21313
rect 41746 21310 41758 21362
rect 45938 21310 45950 21362
rect 46002 21310 46014 21362
rect 1822 21298 1874 21310
rect 44158 21298 44210 21310
rect 1344 21194 78624 21228
rect 1344 21142 10874 21194
rect 10926 21142 10978 21194
rect 11030 21142 11082 21194
rect 11134 21142 30194 21194
rect 30246 21142 30298 21194
rect 30350 21142 30402 21194
rect 30454 21142 49514 21194
rect 49566 21142 49618 21194
rect 49670 21142 49722 21194
rect 49774 21142 68834 21194
rect 68886 21142 68938 21194
rect 68990 21142 69042 21194
rect 69094 21142 78624 21194
rect 1344 21108 78624 21142
rect 2718 21026 2770 21038
rect 2718 20962 2770 20974
rect 6190 21026 6242 21038
rect 73614 21026 73666 21038
rect 24434 20974 24446 21026
rect 24498 21023 24510 21026
rect 25106 21023 25118 21026
rect 24498 20977 25118 21023
rect 24498 20974 24510 20977
rect 25106 20974 25118 20977
rect 25170 20974 25182 21026
rect 25330 20974 25342 21026
rect 25394 21023 25406 21026
rect 25554 21023 25566 21026
rect 25394 20977 25566 21023
rect 25394 20974 25406 20977
rect 25554 20974 25566 20977
rect 25618 20974 25630 21026
rect 46610 20974 46622 21026
rect 46674 21023 46686 21026
rect 47170 21023 47182 21026
rect 46674 20977 47182 21023
rect 46674 20974 46686 20977
rect 47170 20974 47182 20977
rect 47234 20974 47246 21026
rect 6190 20962 6242 20974
rect 73614 20962 73666 20974
rect 11678 20914 11730 20926
rect 17838 20914 17890 20926
rect 16370 20862 16382 20914
rect 16434 20862 16446 20914
rect 17266 20862 17278 20914
rect 17330 20862 17342 20914
rect 11678 20850 11730 20862
rect 17838 20850 17890 20862
rect 20750 20914 20802 20926
rect 22990 20914 23042 20926
rect 21410 20862 21422 20914
rect 21474 20862 21486 20914
rect 20750 20850 20802 20862
rect 22990 20850 23042 20862
rect 24222 20914 24274 20926
rect 24222 20850 24274 20862
rect 24670 20914 24722 20926
rect 24670 20850 24722 20862
rect 25118 20914 25170 20926
rect 25118 20850 25170 20862
rect 25678 20914 25730 20926
rect 25678 20850 25730 20862
rect 27134 20914 27186 20926
rect 31166 20914 31218 20926
rect 28242 20862 28254 20914
rect 28306 20862 28318 20914
rect 27134 20850 27186 20862
rect 31166 20850 31218 20862
rect 31614 20914 31666 20926
rect 39006 20914 39058 20926
rect 43598 20914 43650 20926
rect 34738 20862 34750 20914
rect 34802 20862 34814 20914
rect 41010 20862 41022 20914
rect 41074 20862 41086 20914
rect 42690 20862 42702 20914
rect 42754 20862 42766 20914
rect 31614 20850 31666 20862
rect 39006 20850 39058 20862
rect 43598 20850 43650 20862
rect 45166 20914 45218 20926
rect 45166 20850 45218 20862
rect 46846 20914 46898 20926
rect 46846 20850 46898 20862
rect 47182 20914 47234 20926
rect 47182 20850 47234 20862
rect 56814 20914 56866 20926
rect 56814 20850 56866 20862
rect 59054 20914 59106 20926
rect 59054 20850 59106 20862
rect 59390 20914 59442 20926
rect 70030 20914 70082 20926
rect 67218 20862 67230 20914
rect 67282 20862 67294 20914
rect 59390 20850 59442 20862
rect 70030 20850 70082 20862
rect 9998 20802 10050 20814
rect 10782 20802 10834 20814
rect 11454 20802 11506 20814
rect 16942 20802 16994 20814
rect 21534 20802 21586 20814
rect 1810 20750 1822 20802
rect 1874 20750 1886 20802
rect 6962 20750 6974 20802
rect 7026 20750 7038 20802
rect 7970 20750 7982 20802
rect 8034 20750 8046 20802
rect 10434 20750 10446 20802
rect 10498 20750 10510 20802
rect 11218 20750 11230 20802
rect 11282 20750 11294 20802
rect 13570 20750 13582 20802
rect 13634 20750 13646 20802
rect 21298 20750 21310 20802
rect 21362 20750 21374 20802
rect 9998 20738 10050 20750
rect 10782 20738 10834 20750
rect 11454 20738 11506 20750
rect 16942 20738 16994 20750
rect 21534 20738 21586 20750
rect 21870 20802 21922 20814
rect 21870 20738 21922 20750
rect 25902 20802 25954 20814
rect 29486 20802 29538 20814
rect 27458 20750 27470 20802
rect 27522 20750 27534 20802
rect 28354 20750 28366 20802
rect 28418 20750 28430 20802
rect 25902 20738 25954 20750
rect 29486 20738 29538 20750
rect 30830 20802 30882 20814
rect 36094 20802 36146 20814
rect 32386 20750 32398 20802
rect 32450 20750 32462 20802
rect 33730 20750 33742 20802
rect 33794 20750 33806 20802
rect 30830 20738 30882 20750
rect 36094 20738 36146 20750
rect 37326 20802 37378 20814
rect 37326 20738 37378 20750
rect 41806 20802 41858 20814
rect 41806 20738 41858 20750
rect 42366 20802 42418 20814
rect 42366 20738 42418 20750
rect 44942 20802 44994 20814
rect 44942 20738 44994 20750
rect 45278 20802 45330 20814
rect 45278 20738 45330 20750
rect 45390 20802 45442 20814
rect 49870 20802 49922 20814
rect 52670 20802 52722 20814
rect 62078 20802 62130 20814
rect 48738 20750 48750 20802
rect 48802 20750 48814 20802
rect 50754 20750 50766 20802
rect 50818 20750 50830 20802
rect 53666 20750 53678 20802
rect 53730 20750 53742 20802
rect 56578 20750 56590 20802
rect 56642 20750 56654 20802
rect 58034 20750 58046 20802
rect 58098 20750 58110 20802
rect 61394 20750 61406 20802
rect 61458 20750 61470 20802
rect 45390 20738 45442 20750
rect 49870 20738 49922 20750
rect 52670 20738 52722 20750
rect 62078 20738 62130 20750
rect 62414 20802 62466 20814
rect 71374 20802 71426 20814
rect 62850 20750 62862 20802
rect 62914 20750 62926 20802
rect 63746 20750 63758 20802
rect 63810 20750 63822 20802
rect 64418 20750 64430 20802
rect 64482 20750 64494 20802
rect 73714 20750 73726 20802
rect 73778 20750 73790 20802
rect 62414 20738 62466 20750
rect 71374 20738 71426 20750
rect 4622 20690 4674 20702
rect 4622 20626 4674 20638
rect 4958 20690 5010 20702
rect 4958 20626 5010 20638
rect 5854 20690 5906 20702
rect 7758 20690 7810 20702
rect 16718 20690 16770 20702
rect 6850 20638 6862 20690
rect 6914 20638 6926 20690
rect 14242 20638 14254 20690
rect 14306 20638 14318 20690
rect 5854 20626 5906 20638
rect 7758 20626 7810 20638
rect 16718 20626 16770 20638
rect 21758 20690 21810 20702
rect 21758 20626 21810 20638
rect 22430 20690 22482 20702
rect 22430 20626 22482 20638
rect 22542 20690 22594 20702
rect 38222 20690 38274 20702
rect 26226 20638 26238 20690
rect 26290 20638 26302 20690
rect 28130 20638 28142 20690
rect 28194 20638 28206 20690
rect 29810 20638 29822 20690
rect 29874 20638 29886 20690
rect 33282 20638 33294 20690
rect 33346 20638 33358 20690
rect 34626 20638 34638 20690
rect 34690 20638 34702 20690
rect 22542 20626 22594 20638
rect 38222 20626 38274 20638
rect 40126 20690 40178 20702
rect 40126 20626 40178 20638
rect 40238 20690 40290 20702
rect 40238 20626 40290 20638
rect 43038 20690 43090 20702
rect 50206 20690 50258 20702
rect 49074 20638 49086 20690
rect 49138 20638 49150 20690
rect 43038 20626 43090 20638
rect 50206 20626 50258 20638
rect 50318 20690 50370 20702
rect 51774 20690 51826 20702
rect 50866 20638 50878 20690
rect 50930 20638 50942 20690
rect 50318 20626 50370 20638
rect 51774 20626 51826 20638
rect 51886 20690 51938 20702
rect 51886 20626 51938 20638
rect 55582 20690 55634 20702
rect 63982 20690 64034 20702
rect 63186 20638 63198 20690
rect 63250 20638 63262 20690
rect 65090 20638 65102 20690
rect 65154 20638 65166 20690
rect 72818 20638 72830 20690
rect 72882 20638 72894 20690
rect 55582 20626 55634 20638
rect 63982 20626 64034 20638
rect 10110 20578 10162 20590
rect 10110 20514 10162 20526
rect 10670 20578 10722 20590
rect 12574 20578 12626 20590
rect 11666 20526 11678 20578
rect 11730 20526 11742 20578
rect 12226 20526 12238 20578
rect 12290 20526 12302 20578
rect 10670 20514 10722 20526
rect 12574 20514 12626 20526
rect 17166 20578 17218 20590
rect 17166 20514 17218 20526
rect 17278 20578 17330 20590
rect 17278 20514 17330 20526
rect 18286 20578 18338 20590
rect 19294 20578 19346 20590
rect 18946 20526 18958 20578
rect 19010 20526 19022 20578
rect 18286 20514 18338 20526
rect 19294 20514 19346 20526
rect 19742 20578 19794 20590
rect 19742 20514 19794 20526
rect 22206 20578 22258 20590
rect 22206 20514 22258 20526
rect 23550 20578 23602 20590
rect 23550 20514 23602 20526
rect 26574 20578 26626 20590
rect 26574 20514 26626 20526
rect 30270 20578 30322 20590
rect 30270 20514 30322 20526
rect 38670 20578 38722 20590
rect 38670 20514 38722 20526
rect 40462 20578 40514 20590
rect 40462 20514 40514 20526
rect 41470 20578 41522 20590
rect 41470 20514 41522 20526
rect 43934 20578 43986 20590
rect 43934 20514 43986 20526
rect 45054 20578 45106 20590
rect 45054 20514 45106 20526
rect 45950 20578 46002 20590
rect 45950 20514 46002 20526
rect 47630 20578 47682 20590
rect 50542 20578 50594 20590
rect 52110 20578 52162 20590
rect 49298 20526 49310 20578
rect 49362 20526 49374 20578
rect 51090 20526 51102 20578
rect 51154 20526 51166 20578
rect 47630 20514 47682 20526
rect 50542 20514 50594 20526
rect 52110 20514 52162 20526
rect 52782 20578 52834 20590
rect 52782 20514 52834 20526
rect 53006 20578 53058 20590
rect 53006 20514 53058 20526
rect 53454 20578 53506 20590
rect 53454 20514 53506 20526
rect 55134 20578 55186 20590
rect 55134 20514 55186 20526
rect 58270 20578 58322 20590
rect 58270 20514 58322 20526
rect 60958 20578 61010 20590
rect 60958 20514 61010 20526
rect 61630 20578 61682 20590
rect 61630 20514 61682 20526
rect 74174 20578 74226 20590
rect 74174 20514 74226 20526
rect 75294 20578 75346 20590
rect 75294 20514 75346 20526
rect 76302 20578 76354 20590
rect 76302 20514 76354 20526
rect 1344 20410 78784 20444
rect 1344 20358 20534 20410
rect 20586 20358 20638 20410
rect 20690 20358 20742 20410
rect 20794 20358 39854 20410
rect 39906 20358 39958 20410
rect 40010 20358 40062 20410
rect 40114 20358 59174 20410
rect 59226 20358 59278 20410
rect 59330 20358 59382 20410
rect 59434 20358 78494 20410
rect 78546 20358 78598 20410
rect 78650 20358 78702 20410
rect 78754 20358 78784 20410
rect 1344 20324 78784 20358
rect 7758 20242 7810 20254
rect 7758 20178 7810 20190
rect 25790 20242 25842 20254
rect 25790 20178 25842 20190
rect 26350 20242 26402 20254
rect 26350 20178 26402 20190
rect 30158 20242 30210 20254
rect 30158 20178 30210 20190
rect 44494 20242 44546 20254
rect 44494 20178 44546 20190
rect 49086 20242 49138 20254
rect 49086 20178 49138 20190
rect 49870 20242 49922 20254
rect 56702 20242 56754 20254
rect 51874 20190 51886 20242
rect 51938 20190 51950 20242
rect 49870 20178 49922 20190
rect 56702 20178 56754 20190
rect 69022 20242 69074 20254
rect 69022 20178 69074 20190
rect 69470 20242 69522 20254
rect 69470 20178 69522 20190
rect 3166 20130 3218 20142
rect 3166 20066 3218 20078
rect 3502 20130 3554 20142
rect 3502 20066 3554 20078
rect 7310 20130 7362 20142
rect 9998 20130 10050 20142
rect 8754 20078 8766 20130
rect 8818 20078 8830 20130
rect 7310 20066 7362 20078
rect 9998 20066 10050 20078
rect 10446 20130 10498 20142
rect 10446 20066 10498 20078
rect 16270 20130 16322 20142
rect 16270 20066 16322 20078
rect 16718 20130 16770 20142
rect 16718 20066 16770 20078
rect 28366 20130 28418 20142
rect 28366 20066 28418 20078
rect 32174 20130 32226 20142
rect 32174 20066 32226 20078
rect 32510 20130 32562 20142
rect 32510 20066 32562 20078
rect 33518 20130 33570 20142
rect 33518 20066 33570 20078
rect 33742 20130 33794 20142
rect 33742 20066 33794 20078
rect 33966 20130 34018 20142
rect 42478 20130 42530 20142
rect 36306 20078 36318 20130
rect 36370 20078 36382 20130
rect 33966 20066 34018 20078
rect 42478 20066 42530 20078
rect 42702 20130 42754 20142
rect 42702 20066 42754 20078
rect 43262 20130 43314 20142
rect 43262 20066 43314 20078
rect 44830 20130 44882 20142
rect 44830 20066 44882 20078
rect 45278 20130 45330 20142
rect 45278 20066 45330 20078
rect 45838 20130 45890 20142
rect 45838 20066 45890 20078
rect 48750 20130 48802 20142
rect 48750 20066 48802 20078
rect 48862 20130 48914 20142
rect 48862 20066 48914 20078
rect 49422 20130 49474 20142
rect 64542 20130 64594 20142
rect 69694 20130 69746 20142
rect 50978 20078 50990 20130
rect 51042 20078 51054 20130
rect 55010 20078 55022 20130
rect 55074 20078 55086 20130
rect 59154 20078 59166 20130
rect 59218 20078 59230 20130
rect 61170 20078 61182 20130
rect 61234 20078 61246 20130
rect 65090 20078 65102 20130
rect 65154 20078 65166 20130
rect 65538 20078 65550 20130
rect 65602 20078 65614 20130
rect 70578 20078 70590 20130
rect 70642 20078 70654 20130
rect 49422 20066 49474 20078
rect 64542 20066 64594 20078
rect 69694 20066 69746 20078
rect 8094 20018 8146 20030
rect 9662 20018 9714 20030
rect 8866 19966 8878 20018
rect 8930 19966 8942 20018
rect 8094 19954 8146 19966
rect 9662 19954 9714 19966
rect 10110 20018 10162 20030
rect 10110 19954 10162 19966
rect 10894 20018 10946 20030
rect 16046 20018 16098 20030
rect 11666 19966 11678 20018
rect 11730 19966 11742 20018
rect 13010 19966 13022 20018
rect 13074 19966 13086 20018
rect 13458 19966 13470 20018
rect 13522 19966 13534 20018
rect 14466 19966 14478 20018
rect 14530 19966 14542 20018
rect 10894 19954 10946 19966
rect 16046 19954 16098 19966
rect 16382 20018 16434 20030
rect 27134 20018 27186 20030
rect 29598 20018 29650 20030
rect 23090 19966 23102 20018
rect 23154 19966 23166 20018
rect 27794 19966 27806 20018
rect 27858 19966 27870 20018
rect 16382 19954 16434 19966
rect 27134 19954 27186 19966
rect 29598 19954 29650 19966
rect 31054 20018 31106 20030
rect 31054 19954 31106 19966
rect 34526 20018 34578 20030
rect 37550 20018 37602 20030
rect 60846 20018 60898 20030
rect 35410 19966 35422 20018
rect 35474 19966 35486 20018
rect 37762 19966 37774 20018
rect 37826 19966 37838 20018
rect 40226 19966 40238 20018
rect 40290 19966 40302 20018
rect 41906 19966 41918 20018
rect 41970 19966 41982 20018
rect 50866 19966 50878 20018
rect 50930 19966 50942 20018
rect 52882 19966 52894 20018
rect 52946 19966 52958 20018
rect 54338 19966 54350 20018
rect 54402 19966 54414 20018
rect 59938 19966 59950 20018
rect 60002 19966 60014 20018
rect 34526 19954 34578 19966
rect 37550 19954 37602 19966
rect 60846 19954 60898 19966
rect 64878 20018 64930 20030
rect 64878 19954 64930 19966
rect 66110 20018 66162 20030
rect 66110 19954 66162 19966
rect 66670 20018 66722 20030
rect 66670 19954 66722 19966
rect 69582 20018 69634 20030
rect 69582 19954 69634 19966
rect 69806 20018 69858 20030
rect 71262 20018 71314 20030
rect 70018 19966 70030 20018
rect 70082 19966 70094 20018
rect 70802 19966 70814 20018
rect 70866 19966 70878 20018
rect 72706 19966 72718 20018
rect 72770 19966 72782 20018
rect 75730 19966 75742 20018
rect 75794 19966 75806 20018
rect 69806 19954 69858 19966
rect 71262 19954 71314 19966
rect 3950 19906 4002 19918
rect 3950 19842 4002 19854
rect 4398 19906 4450 19918
rect 17502 19906 17554 19918
rect 14802 19854 14814 19906
rect 14866 19854 14878 19906
rect 4398 19842 4450 19854
rect 17502 19842 17554 19854
rect 17950 19906 18002 19918
rect 23550 19906 23602 19918
rect 20178 19854 20190 19906
rect 20242 19854 20254 19906
rect 22306 19854 22318 19906
rect 22370 19854 22382 19906
rect 17950 19842 18002 19854
rect 23550 19842 23602 19854
rect 23998 19906 24050 19918
rect 43710 19906 43762 19918
rect 26674 19854 26686 19906
rect 26738 19854 26750 19906
rect 31490 19854 31502 19906
rect 31554 19854 31566 19906
rect 35522 19854 35534 19906
rect 35586 19854 35598 19906
rect 41346 19854 41358 19906
rect 41410 19854 41422 19906
rect 23998 19842 24050 19854
rect 43710 19842 43762 19854
rect 50318 19906 50370 19918
rect 50318 19842 50370 19854
rect 55470 19906 55522 19918
rect 55470 19842 55522 19854
rect 56030 19906 56082 19918
rect 63870 19906 63922 19918
rect 57026 19854 57038 19906
rect 57090 19854 57102 19906
rect 56030 19842 56082 19854
rect 63870 19842 63922 19854
rect 72494 19906 72546 19918
rect 72494 19842 72546 19854
rect 77982 19906 78034 19918
rect 77982 19842 78034 19854
rect 3838 19794 3890 19806
rect 3838 19730 3890 19742
rect 10558 19794 10610 19806
rect 10558 19730 10610 19742
rect 11006 19794 11058 19806
rect 16830 19794 16882 19806
rect 23438 19794 23490 19806
rect 42814 19794 42866 19806
rect 15026 19742 15038 19794
rect 15090 19742 15102 19794
rect 17378 19742 17390 19794
rect 17442 19791 17454 19794
rect 17826 19791 17838 19794
rect 17442 19745 17838 19791
rect 17442 19742 17454 19745
rect 17826 19742 17838 19745
rect 17890 19742 17902 19794
rect 33170 19742 33182 19794
rect 33234 19742 33246 19794
rect 38770 19742 38782 19794
rect 38834 19742 38846 19794
rect 11006 19730 11058 19742
rect 16830 19730 16882 19742
rect 23438 19730 23490 19742
rect 42814 19730 42866 19742
rect 71598 19794 71650 19806
rect 71598 19730 71650 19742
rect 75070 19794 75122 19806
rect 75070 19730 75122 19742
rect 1344 19626 78624 19660
rect 1344 19574 10874 19626
rect 10926 19574 10978 19626
rect 11030 19574 11082 19626
rect 11134 19574 30194 19626
rect 30246 19574 30298 19626
rect 30350 19574 30402 19626
rect 30454 19574 49514 19626
rect 49566 19574 49618 19626
rect 49670 19574 49722 19626
rect 49774 19574 68834 19626
rect 68886 19574 68938 19626
rect 68990 19574 69042 19626
rect 69094 19574 78624 19626
rect 1344 19540 78624 19574
rect 23102 19458 23154 19470
rect 18162 19406 18174 19458
rect 18226 19406 18238 19458
rect 23102 19394 23154 19406
rect 27470 19458 27522 19470
rect 27470 19394 27522 19406
rect 29934 19458 29986 19470
rect 29934 19394 29986 19406
rect 58270 19458 58322 19470
rect 69234 19406 69246 19458
rect 69298 19406 69310 19458
rect 58270 19394 58322 19406
rect 13806 19346 13858 19358
rect 2706 19294 2718 19346
rect 2770 19294 2782 19346
rect 4834 19294 4846 19346
rect 4898 19294 4910 19346
rect 13806 19282 13858 19294
rect 14702 19346 14754 19358
rect 14702 19282 14754 19294
rect 21758 19346 21810 19358
rect 27022 19346 27074 19358
rect 22306 19294 22318 19346
rect 22370 19343 22382 19346
rect 22642 19343 22654 19346
rect 22370 19297 22654 19343
rect 22370 19294 22382 19297
rect 22642 19294 22654 19297
rect 22706 19294 22718 19346
rect 21758 19282 21810 19294
rect 27022 19282 27074 19294
rect 28590 19346 28642 19358
rect 28590 19282 28642 19294
rect 33742 19346 33794 19358
rect 51438 19346 51490 19358
rect 61070 19346 61122 19358
rect 38882 19294 38894 19346
rect 38946 19294 38958 19346
rect 40562 19294 40574 19346
rect 40626 19294 40638 19346
rect 53442 19294 53454 19346
rect 53506 19294 53518 19346
rect 55570 19294 55582 19346
rect 55634 19294 55646 19346
rect 33742 19282 33794 19294
rect 51438 19282 51490 19294
rect 61070 19282 61122 19294
rect 12126 19234 12178 19246
rect 2034 19182 2046 19234
rect 2098 19182 2110 19234
rect 12126 19170 12178 19182
rect 15262 19234 15314 19246
rect 15262 19170 15314 19182
rect 15710 19234 15762 19246
rect 15710 19170 15762 19182
rect 16494 19234 16546 19246
rect 16494 19170 16546 19182
rect 16942 19234 16994 19246
rect 16942 19170 16994 19182
rect 17278 19234 17330 19246
rect 17278 19170 17330 19182
rect 18622 19234 18674 19246
rect 22878 19234 22930 19246
rect 22194 19182 22206 19234
rect 22258 19182 22270 19234
rect 18622 19170 18674 19182
rect 22878 19170 22930 19182
rect 23326 19234 23378 19246
rect 23326 19170 23378 19182
rect 26126 19234 26178 19246
rect 26126 19170 26178 19182
rect 26574 19234 26626 19246
rect 26574 19170 26626 19182
rect 27358 19234 27410 19246
rect 27358 19170 27410 19182
rect 27806 19234 27858 19246
rect 27806 19170 27858 19182
rect 28142 19234 28194 19246
rect 28142 19170 28194 19182
rect 29038 19234 29090 19246
rect 29710 19234 29762 19246
rect 33182 19234 33234 19246
rect 42590 19234 42642 19246
rect 29362 19182 29374 19234
rect 29426 19182 29438 19234
rect 30258 19182 30270 19234
rect 30322 19182 30334 19234
rect 34066 19182 34078 19234
rect 34130 19182 34142 19234
rect 35410 19182 35422 19234
rect 35474 19182 35486 19234
rect 36418 19182 36430 19234
rect 36482 19182 36494 19234
rect 39106 19182 39118 19234
rect 39170 19182 39182 19234
rect 40674 19182 40686 19234
rect 40738 19182 40750 19234
rect 42130 19182 42142 19234
rect 42194 19182 42206 19234
rect 29038 19170 29090 19182
rect 29710 19170 29762 19182
rect 33182 19170 33234 19182
rect 42590 19170 42642 19182
rect 43486 19234 43538 19246
rect 56702 19234 56754 19246
rect 43922 19182 43934 19234
rect 43986 19182 43998 19234
rect 47058 19182 47070 19234
rect 47122 19182 47134 19234
rect 52770 19182 52782 19234
rect 52834 19182 52846 19234
rect 43486 19170 43538 19182
rect 56702 19170 56754 19182
rect 57262 19234 57314 19246
rect 57262 19170 57314 19182
rect 57822 19234 57874 19246
rect 57822 19170 57874 19182
rect 58606 19234 58658 19246
rect 68910 19234 68962 19246
rect 59266 19182 59278 19234
rect 59330 19182 59342 19234
rect 61842 19182 61854 19234
rect 61906 19182 61918 19234
rect 58606 19170 58658 19182
rect 68910 19170 68962 19182
rect 10894 19122 10946 19134
rect 12350 19122 12402 19134
rect 11330 19070 11342 19122
rect 11394 19070 11406 19122
rect 11778 19070 11790 19122
rect 11842 19070 11854 19122
rect 10894 19058 10946 19070
rect 12350 19058 12402 19070
rect 14814 19122 14866 19134
rect 14814 19058 14866 19070
rect 16270 19122 16322 19134
rect 18958 19122 19010 19134
rect 18274 19070 18286 19122
rect 18338 19070 18350 19122
rect 16270 19058 16322 19070
rect 18958 19058 19010 19070
rect 21646 19122 21698 19134
rect 27918 19122 27970 19134
rect 44942 19122 44994 19134
rect 24882 19070 24894 19122
rect 24946 19070 24958 19122
rect 35634 19070 35646 19122
rect 35698 19070 35710 19122
rect 41458 19070 41470 19122
rect 41522 19070 41534 19122
rect 43026 19070 43038 19122
rect 43090 19070 43102 19122
rect 21646 19058 21698 19070
rect 27918 19058 27970 19070
rect 44942 19058 44994 19070
rect 47518 19122 47570 19134
rect 47518 19058 47570 19070
rect 56814 19122 56866 19134
rect 61406 19122 61458 19134
rect 59378 19070 59390 19122
rect 59442 19070 59454 19122
rect 56814 19058 56866 19070
rect 61406 19058 61458 19070
rect 9214 19010 9266 19022
rect 9214 18946 9266 18958
rect 12686 19010 12738 19022
rect 12686 18946 12738 18958
rect 14366 19010 14418 19022
rect 14366 18946 14418 18958
rect 14590 19010 14642 19022
rect 14590 18946 14642 18958
rect 16046 19010 16098 19022
rect 16046 18946 16098 18958
rect 16382 19010 16434 19022
rect 16382 18946 16434 18958
rect 18846 19010 18898 19022
rect 18846 18946 18898 18958
rect 20750 19010 20802 19022
rect 20750 18946 20802 18958
rect 21870 19010 21922 19022
rect 21870 18946 21922 18958
rect 23774 19010 23826 19022
rect 23774 18946 23826 18958
rect 24222 19010 24274 19022
rect 24222 18946 24274 18958
rect 25230 19010 25282 19022
rect 25230 18946 25282 18958
rect 25678 19010 25730 19022
rect 25678 18946 25730 18958
rect 29598 19010 29650 19022
rect 29598 18946 29650 18958
rect 30046 19010 30098 19022
rect 30046 18946 30098 18958
rect 37326 19010 37378 19022
rect 37326 18946 37378 18958
rect 38110 19010 38162 19022
rect 56142 19010 56194 19022
rect 41570 18958 41582 19010
rect 41634 18958 41646 19010
rect 38110 18946 38162 18958
rect 56142 18946 56194 18958
rect 56926 19010 56978 19022
rect 56926 18946 56978 18958
rect 67902 19010 67954 19022
rect 67902 18946 67954 18958
rect 68350 19010 68402 19022
rect 69249 19007 69295 19406
rect 74958 19346 75010 19358
rect 78094 19346 78146 19358
rect 70242 19294 70254 19346
rect 70306 19294 70318 19346
rect 71138 19294 71150 19346
rect 71202 19294 71214 19346
rect 76626 19294 76638 19346
rect 76690 19294 76702 19346
rect 74958 19282 75010 19294
rect 78094 19282 78146 19294
rect 70366 19234 70418 19246
rect 70366 19170 70418 19182
rect 70590 19234 70642 19246
rect 76190 19234 76242 19246
rect 73938 19182 73950 19234
rect 74002 19182 74014 19234
rect 70590 19170 70642 19182
rect 76190 19170 76242 19182
rect 69582 19122 69634 19134
rect 69582 19058 69634 19070
rect 69694 19122 69746 19134
rect 69694 19058 69746 19070
rect 70814 19122 70866 19134
rect 75630 19122 75682 19134
rect 73266 19070 73278 19122
rect 73330 19070 73342 19122
rect 70814 19058 70866 19070
rect 75630 19058 75682 19070
rect 77646 19122 77698 19134
rect 77646 19058 77698 19070
rect 77982 19122 78034 19134
rect 77982 19058 78034 19070
rect 69918 19010 69970 19022
rect 69346 19007 69358 19010
rect 69249 18961 69358 19007
rect 69346 18958 69358 18961
rect 69410 18958 69422 19010
rect 68350 18946 68402 18958
rect 69918 18946 69970 18958
rect 70254 19010 70306 19022
rect 70254 18946 70306 18958
rect 74398 19010 74450 19022
rect 74398 18946 74450 18958
rect 75294 19010 75346 19022
rect 75294 18946 75346 18958
rect 75518 19010 75570 19022
rect 75518 18946 75570 18958
rect 77198 19010 77250 19022
rect 77198 18946 77250 18958
rect 77422 19010 77474 19022
rect 77422 18946 77474 18958
rect 77534 19010 77586 19022
rect 77534 18946 77586 18958
rect 1344 18842 78784 18876
rect 1344 18790 20534 18842
rect 20586 18790 20638 18842
rect 20690 18790 20742 18842
rect 20794 18790 39854 18842
rect 39906 18790 39958 18842
rect 40010 18790 40062 18842
rect 40114 18790 59174 18842
rect 59226 18790 59278 18842
rect 59330 18790 59382 18842
rect 59434 18790 78494 18842
rect 78546 18790 78598 18842
rect 78650 18790 78702 18842
rect 78754 18790 78784 18842
rect 1344 18756 78784 18790
rect 4734 18674 4786 18686
rect 4734 18610 4786 18622
rect 19966 18674 20018 18686
rect 19966 18610 20018 18622
rect 21870 18674 21922 18686
rect 21870 18610 21922 18622
rect 28702 18674 28754 18686
rect 42478 18674 42530 18686
rect 36418 18622 36430 18674
rect 36482 18622 36494 18674
rect 28702 18610 28754 18622
rect 42478 18610 42530 18622
rect 69582 18674 69634 18686
rect 69582 18610 69634 18622
rect 69694 18674 69746 18686
rect 70578 18622 70590 18674
rect 70642 18622 70654 18674
rect 69694 18610 69746 18622
rect 17726 18562 17778 18574
rect 20750 18562 20802 18574
rect 5842 18510 5854 18562
rect 5906 18510 5918 18562
rect 19058 18510 19070 18562
rect 19122 18510 19134 18562
rect 17726 18498 17778 18510
rect 20750 18498 20802 18510
rect 20862 18562 20914 18574
rect 34974 18562 35026 18574
rect 55582 18562 55634 18574
rect 60734 18562 60786 18574
rect 63086 18562 63138 18574
rect 22530 18510 22542 18562
rect 22594 18510 22606 18562
rect 26002 18510 26014 18562
rect 26066 18510 26078 18562
rect 35522 18510 35534 18562
rect 35586 18510 35598 18562
rect 37426 18510 37438 18562
rect 37490 18510 37502 18562
rect 43474 18510 43486 18562
rect 43538 18510 43550 18562
rect 48962 18510 48974 18562
rect 49026 18510 49038 18562
rect 54898 18510 54910 18562
rect 54962 18510 54974 18562
rect 56802 18510 56814 18562
rect 56866 18510 56878 18562
rect 62178 18510 62190 18562
rect 62242 18510 62254 18562
rect 20862 18498 20914 18510
rect 34974 18498 35026 18510
rect 55582 18498 55634 18510
rect 60734 18498 60786 18510
rect 63086 18498 63138 18510
rect 70478 18562 70530 18574
rect 71362 18510 71374 18562
rect 71426 18510 71438 18562
rect 72818 18510 72830 18562
rect 72882 18510 72894 18562
rect 77410 18510 77422 18562
rect 77474 18510 77486 18562
rect 70478 18498 70530 18510
rect 6414 18450 6466 18462
rect 18062 18450 18114 18462
rect 3826 18398 3838 18450
rect 3890 18398 3902 18450
rect 5730 18398 5742 18450
rect 5794 18398 5806 18450
rect 11890 18398 11902 18450
rect 11954 18398 11966 18450
rect 12898 18398 12910 18450
rect 12962 18398 12974 18450
rect 13122 18398 13134 18450
rect 13186 18398 13198 18450
rect 14578 18398 14590 18450
rect 14642 18398 14654 18450
rect 17378 18398 17390 18450
rect 17442 18398 17454 18450
rect 6414 18386 6466 18398
rect 18062 18386 18114 18398
rect 19630 18450 19682 18462
rect 21086 18450 21138 18462
rect 23886 18450 23938 18462
rect 20178 18398 20190 18450
rect 20242 18398 20254 18450
rect 20402 18398 20414 18450
rect 20466 18398 20478 18450
rect 21410 18398 21422 18450
rect 21474 18398 21486 18450
rect 21634 18398 21646 18450
rect 21698 18398 21710 18450
rect 23426 18398 23438 18450
rect 23490 18398 23502 18450
rect 19630 18386 19682 18398
rect 21086 18386 21138 18398
rect 23886 18386 23938 18398
rect 23998 18450 24050 18462
rect 23998 18386 24050 18398
rect 26350 18450 26402 18462
rect 29038 18450 29090 18462
rect 27682 18398 27694 18450
rect 27746 18398 27758 18450
rect 26350 18386 26402 18398
rect 29038 18386 29090 18398
rect 29934 18450 29986 18462
rect 29934 18386 29986 18398
rect 30494 18450 30546 18462
rect 30494 18386 30546 18398
rect 34302 18450 34354 18462
rect 39230 18450 39282 18462
rect 34626 18398 34638 18450
rect 34690 18398 34702 18450
rect 36530 18398 36542 18450
rect 36594 18398 36606 18450
rect 37986 18398 37998 18450
rect 38050 18398 38062 18450
rect 34302 18386 34354 18398
rect 39230 18386 39282 18398
rect 40014 18450 40066 18462
rect 53790 18450 53842 18462
rect 42018 18398 42030 18450
rect 42082 18398 42094 18450
rect 43586 18398 43598 18450
rect 43650 18398 43662 18450
rect 44258 18398 44270 18450
rect 44322 18398 44334 18450
rect 44706 18398 44718 18450
rect 44770 18398 44782 18450
rect 45378 18398 45390 18450
rect 45442 18398 45454 18450
rect 48738 18398 48750 18450
rect 48802 18398 48814 18450
rect 40014 18386 40066 18398
rect 53790 18386 53842 18398
rect 54126 18450 54178 18462
rect 55694 18450 55746 18462
rect 54674 18398 54686 18450
rect 54738 18398 54750 18450
rect 55346 18398 55358 18450
rect 55410 18398 55422 18450
rect 54126 18386 54178 18398
rect 55694 18386 55746 18398
rect 55806 18450 55858 18462
rect 56478 18450 56530 18462
rect 66670 18450 66722 18462
rect 56018 18398 56030 18450
rect 56082 18398 56094 18450
rect 56690 18398 56702 18450
rect 56754 18398 56766 18450
rect 57250 18398 57262 18450
rect 57314 18398 57326 18450
rect 58034 18398 58046 18450
rect 58098 18398 58110 18450
rect 60498 18398 60510 18450
rect 60562 18398 60574 18450
rect 61954 18398 61966 18450
rect 62018 18398 62030 18450
rect 62850 18398 62862 18450
rect 62914 18398 62926 18450
rect 65314 18398 65326 18450
rect 65378 18398 65390 18450
rect 55806 18386 55858 18398
rect 56478 18386 56530 18398
rect 66670 18386 66722 18398
rect 67566 18450 67618 18462
rect 67566 18386 67618 18398
rect 68126 18450 68178 18462
rect 68126 18386 68178 18398
rect 69358 18450 69410 18462
rect 69358 18386 69410 18398
rect 69470 18450 69522 18462
rect 69906 18398 69918 18450
rect 69970 18398 69982 18450
rect 70802 18398 70814 18450
rect 70866 18398 70878 18450
rect 71138 18398 71150 18450
rect 71202 18398 71214 18450
rect 73042 18398 73054 18450
rect 73106 18398 73118 18450
rect 73938 18398 73950 18450
rect 74002 18398 74014 18450
rect 78082 18398 78094 18450
rect 78146 18398 78158 18450
rect 69470 18386 69522 18398
rect 1934 18338 1986 18350
rect 16158 18338 16210 18350
rect 14690 18286 14702 18338
rect 14754 18286 14766 18338
rect 1934 18274 1986 18286
rect 16158 18274 16210 18286
rect 16830 18338 16882 18350
rect 16830 18274 16882 18286
rect 20302 18338 20354 18350
rect 20302 18274 20354 18286
rect 24670 18338 24722 18350
rect 24670 18274 24722 18286
rect 26910 18338 26962 18350
rect 26910 18274 26962 18286
rect 27358 18338 27410 18350
rect 40350 18338 40402 18350
rect 53454 18338 53506 18350
rect 28018 18286 28030 18338
rect 28082 18286 28094 18338
rect 29474 18286 29486 18338
rect 29538 18286 29550 18338
rect 41010 18286 41022 18338
rect 41074 18286 41086 18338
rect 42914 18286 42926 18338
rect 42978 18286 42990 18338
rect 46050 18286 46062 18338
rect 46114 18286 46126 18338
rect 48178 18286 48190 18338
rect 48242 18286 48254 18338
rect 49410 18286 49422 18338
rect 49474 18286 49486 18338
rect 27358 18274 27410 18286
rect 40350 18274 40402 18286
rect 53454 18274 53506 18286
rect 60062 18338 60114 18350
rect 60062 18274 60114 18286
rect 61182 18338 61234 18350
rect 61182 18274 61234 18286
rect 63534 18338 63586 18350
rect 63534 18274 63586 18286
rect 64990 18338 65042 18350
rect 68574 18338 68626 18350
rect 65650 18286 65662 18338
rect 65714 18286 65726 18338
rect 67106 18286 67118 18338
rect 67170 18286 67182 18338
rect 72706 18286 72718 18338
rect 72770 18286 72782 18338
rect 75282 18286 75294 18338
rect 75346 18286 75358 18338
rect 64990 18274 65042 18286
rect 68574 18274 68626 18286
rect 5070 18226 5122 18238
rect 21982 18226 22034 18238
rect 45054 18226 45106 18238
rect 15026 18174 15038 18226
rect 15090 18174 15102 18226
rect 18610 18174 18622 18226
rect 18674 18174 18686 18226
rect 22642 18174 22654 18226
rect 22706 18174 22718 18226
rect 26562 18174 26574 18226
rect 26626 18223 26638 18226
rect 26898 18223 26910 18226
rect 26626 18177 26910 18223
rect 26626 18174 26638 18177
rect 26898 18174 26910 18177
rect 26962 18223 26974 18226
rect 27346 18223 27358 18226
rect 26962 18177 27358 18223
rect 26962 18174 26974 18177
rect 27346 18174 27358 18177
rect 27410 18174 27422 18226
rect 5070 18162 5122 18174
rect 21982 18162 22034 18174
rect 45054 18162 45106 18174
rect 61518 18226 61570 18238
rect 61518 18162 61570 18174
rect 1344 18058 78624 18092
rect 1344 18006 10874 18058
rect 10926 18006 10978 18058
rect 11030 18006 11082 18058
rect 11134 18006 30194 18058
rect 30246 18006 30298 18058
rect 30350 18006 30402 18058
rect 30454 18006 49514 18058
rect 49566 18006 49618 18058
rect 49670 18006 49722 18058
rect 49774 18006 68834 18058
rect 68886 18006 68938 18058
rect 68990 18006 69042 18058
rect 69094 18006 78624 18058
rect 1344 17972 78624 18006
rect 17390 17890 17442 17902
rect 17390 17826 17442 17838
rect 17502 17890 17554 17902
rect 17502 17826 17554 17838
rect 17726 17890 17778 17902
rect 17726 17826 17778 17838
rect 20078 17890 20130 17902
rect 20078 17826 20130 17838
rect 22542 17890 22594 17902
rect 22542 17826 22594 17838
rect 23326 17890 23378 17902
rect 53118 17890 53170 17902
rect 40674 17838 40686 17890
rect 40738 17838 40750 17890
rect 23326 17826 23378 17838
rect 53118 17826 53170 17838
rect 63870 17890 63922 17902
rect 63870 17826 63922 17838
rect 6078 17778 6130 17790
rect 5058 17726 5070 17778
rect 5122 17726 5134 17778
rect 6078 17714 6130 17726
rect 12574 17778 12626 17790
rect 14702 17778 14754 17790
rect 13570 17726 13582 17778
rect 13634 17726 13646 17778
rect 12574 17714 12626 17726
rect 14702 17714 14754 17726
rect 15374 17778 15426 17790
rect 21534 17778 21586 17790
rect 23102 17778 23154 17790
rect 49310 17778 49362 17790
rect 16706 17726 16718 17778
rect 16770 17726 16782 17778
rect 18834 17726 18846 17778
rect 18898 17726 18910 17778
rect 22866 17726 22878 17778
rect 22930 17726 22942 17778
rect 24994 17726 25006 17778
rect 25058 17726 25070 17778
rect 29698 17726 29710 17778
rect 29762 17726 29774 17778
rect 33394 17726 33406 17778
rect 33458 17726 33470 17778
rect 37538 17726 37550 17778
rect 37602 17726 37614 17778
rect 40562 17726 40574 17778
rect 40626 17726 40638 17778
rect 45490 17726 45502 17778
rect 45554 17726 45566 17778
rect 15374 17714 15426 17726
rect 21534 17714 21586 17726
rect 23102 17714 23154 17726
rect 49310 17714 49362 17726
rect 54462 17778 54514 17790
rect 65998 17778 66050 17790
rect 69582 17778 69634 17790
rect 57138 17726 57150 17778
rect 57202 17726 57214 17778
rect 57810 17726 57822 17778
rect 57874 17726 57886 17778
rect 58818 17726 58830 17778
rect 58882 17726 58894 17778
rect 61282 17726 61294 17778
rect 61346 17726 61358 17778
rect 63410 17726 63422 17778
rect 63474 17726 63486 17778
rect 66994 17726 67006 17778
rect 67058 17726 67070 17778
rect 68786 17726 68798 17778
rect 68850 17726 68862 17778
rect 54462 17714 54514 17726
rect 65998 17714 66050 17726
rect 69582 17714 69634 17726
rect 73054 17778 73106 17790
rect 73054 17714 73106 17726
rect 75518 17778 75570 17790
rect 75518 17714 75570 17726
rect 12462 17666 12514 17678
rect 2146 17614 2158 17666
rect 2210 17614 2222 17666
rect 6738 17614 6750 17666
rect 6802 17614 6814 17666
rect 12462 17602 12514 17614
rect 14254 17666 14306 17678
rect 20302 17666 20354 17678
rect 15698 17614 15710 17666
rect 15762 17614 15774 17666
rect 14254 17602 14306 17614
rect 20302 17602 20354 17614
rect 20750 17666 20802 17678
rect 20750 17602 20802 17614
rect 29262 17666 29314 17678
rect 29262 17602 29314 17614
rect 31614 17666 31666 17678
rect 43710 17666 43762 17678
rect 47966 17666 48018 17678
rect 57934 17666 57986 17678
rect 58942 17666 58994 17678
rect 64206 17666 64258 17678
rect 76414 17666 76466 17678
rect 76974 17666 77026 17678
rect 33282 17614 33294 17666
rect 33346 17614 33358 17666
rect 34290 17614 34302 17666
rect 34354 17614 34366 17666
rect 34626 17614 34638 17666
rect 34690 17614 34702 17666
rect 35186 17614 35198 17666
rect 35250 17614 35262 17666
rect 36194 17614 36206 17666
rect 36258 17614 36270 17666
rect 36978 17614 36990 17666
rect 37042 17614 37054 17666
rect 40226 17614 40238 17666
rect 40290 17614 40302 17666
rect 41010 17614 41022 17666
rect 41074 17614 41086 17666
rect 43250 17614 43262 17666
rect 43314 17614 43326 17666
rect 46386 17614 46398 17666
rect 46450 17614 46462 17666
rect 48738 17614 48750 17666
rect 48802 17614 48814 17666
rect 53666 17614 53678 17666
rect 53730 17614 53742 17666
rect 55906 17614 55918 17666
rect 55970 17614 55982 17666
rect 56914 17614 56926 17666
rect 56978 17614 56990 17666
rect 58706 17614 58718 17666
rect 58770 17614 58782 17666
rect 59378 17614 59390 17666
rect 59442 17614 59454 17666
rect 60610 17614 60622 17666
rect 60674 17614 60686 17666
rect 64642 17614 64654 17666
rect 64706 17614 64718 17666
rect 65538 17614 65550 17666
rect 65602 17614 65614 17666
rect 69794 17614 69806 17666
rect 69858 17614 69870 17666
rect 71138 17614 71150 17666
rect 71202 17614 71214 17666
rect 71474 17614 71486 17666
rect 71538 17614 71550 17666
rect 72258 17614 72270 17666
rect 72322 17614 72334 17666
rect 74610 17614 74622 17666
rect 74674 17614 74686 17666
rect 76738 17614 76750 17666
rect 76802 17614 76814 17666
rect 31614 17602 31666 17614
rect 43710 17602 43762 17614
rect 47966 17602 48018 17614
rect 57934 17602 57986 17614
rect 58942 17602 58994 17614
rect 64206 17602 64258 17614
rect 76414 17602 76466 17614
rect 76974 17602 77026 17614
rect 7646 17554 7698 17566
rect 15934 17554 15986 17566
rect 2930 17502 2942 17554
rect 2994 17502 3006 17554
rect 6626 17502 6638 17554
rect 6690 17502 6702 17554
rect 11666 17502 11678 17554
rect 11730 17502 11742 17554
rect 12002 17502 12014 17554
rect 12066 17502 12078 17554
rect 7646 17490 7698 17502
rect 15934 17490 15986 17502
rect 16158 17554 16210 17566
rect 16158 17490 16210 17502
rect 16494 17554 16546 17566
rect 16494 17490 16546 17502
rect 16718 17554 16770 17566
rect 16718 17490 16770 17502
rect 16942 17554 16994 17566
rect 18622 17554 18674 17566
rect 18274 17502 18286 17554
rect 18338 17502 18350 17554
rect 16942 17490 16994 17502
rect 18622 17490 18674 17502
rect 19070 17554 19122 17566
rect 19070 17490 19122 17502
rect 19742 17554 19794 17566
rect 19742 17490 19794 17502
rect 22766 17554 22818 17566
rect 30718 17554 30770 17566
rect 26786 17502 26798 17554
rect 26850 17502 26862 17554
rect 27906 17502 27918 17554
rect 27970 17502 27982 17554
rect 22766 17490 22818 17502
rect 30718 17490 30770 17502
rect 31278 17554 31330 17566
rect 44270 17554 44322 17566
rect 33618 17502 33630 17554
rect 33682 17502 33694 17554
rect 34178 17502 34190 17554
rect 34242 17502 34254 17554
rect 35410 17502 35422 17554
rect 35474 17502 35486 17554
rect 36082 17502 36094 17554
rect 36146 17502 36158 17554
rect 38658 17502 38670 17554
rect 38722 17502 38734 17554
rect 39330 17502 39342 17554
rect 39394 17502 39406 17554
rect 31278 17490 31330 17502
rect 44270 17490 44322 17502
rect 47182 17554 47234 17566
rect 47182 17490 47234 17502
rect 47630 17554 47682 17566
rect 51326 17554 51378 17566
rect 48626 17502 48638 17554
rect 48690 17502 48702 17554
rect 47630 17490 47682 17502
rect 51326 17490 51378 17502
rect 52782 17554 52834 17566
rect 58382 17554 58434 17566
rect 73726 17554 73778 17566
rect 53890 17502 53902 17554
rect 53954 17502 53966 17554
rect 55458 17502 55470 17554
rect 55522 17502 55534 17554
rect 64978 17502 64990 17554
rect 65042 17502 65054 17554
rect 52782 17490 52834 17502
rect 58382 17490 58434 17502
rect 73726 17490 73778 17502
rect 77198 17554 77250 17566
rect 77198 17490 77250 17502
rect 77310 17554 77362 17566
rect 77310 17490 77362 17502
rect 5742 17442 5794 17454
rect 5742 17378 5794 17390
rect 7310 17442 7362 17454
rect 7310 17378 7362 17390
rect 8094 17442 8146 17454
rect 8094 17378 8146 17390
rect 12910 17442 12962 17454
rect 12910 17378 12962 17390
rect 16270 17442 16322 17454
rect 16270 17378 16322 17390
rect 18846 17442 18898 17454
rect 18846 17378 18898 17390
rect 19966 17442 20018 17454
rect 19966 17378 20018 17390
rect 22094 17442 22146 17454
rect 24110 17442 24162 17454
rect 23762 17390 23774 17442
rect 23826 17390 23838 17442
rect 22094 17378 22146 17390
rect 24110 17378 24162 17390
rect 24558 17442 24610 17454
rect 24558 17378 24610 17390
rect 25566 17442 25618 17454
rect 25566 17378 25618 17390
rect 27134 17442 27186 17454
rect 27134 17378 27186 17390
rect 27694 17442 27746 17454
rect 27694 17378 27746 17390
rect 28254 17442 28306 17454
rect 28254 17378 28306 17390
rect 32174 17442 32226 17454
rect 32174 17378 32226 17390
rect 44046 17442 44098 17454
rect 44046 17378 44098 17390
rect 44382 17442 44434 17454
rect 44382 17378 44434 17390
rect 46846 17442 46898 17454
rect 46846 17378 46898 17390
rect 50990 17442 51042 17454
rect 50990 17378 51042 17390
rect 57822 17442 57874 17454
rect 57822 17378 57874 17390
rect 58158 17442 58210 17454
rect 58158 17378 58210 17390
rect 59166 17442 59218 17454
rect 59166 17378 59218 17390
rect 66558 17442 66610 17454
rect 66558 17378 66610 17390
rect 67902 17442 67954 17454
rect 67902 17378 67954 17390
rect 68350 17442 68402 17454
rect 68350 17378 68402 17390
rect 75182 17442 75234 17454
rect 75182 17378 75234 17390
rect 75630 17442 75682 17454
rect 75630 17378 75682 17390
rect 76190 17442 76242 17454
rect 76190 17378 76242 17390
rect 76302 17442 76354 17454
rect 76302 17378 76354 17390
rect 1344 17274 78784 17308
rect 1344 17222 20534 17274
rect 20586 17222 20638 17274
rect 20690 17222 20742 17274
rect 20794 17222 39854 17274
rect 39906 17222 39958 17274
rect 40010 17222 40062 17274
rect 40114 17222 59174 17274
rect 59226 17222 59278 17274
rect 59330 17222 59382 17274
rect 59434 17222 78494 17274
rect 78546 17222 78598 17274
rect 78650 17222 78702 17274
rect 78754 17222 78784 17274
rect 1344 17188 78784 17222
rect 11678 17106 11730 17118
rect 23102 17106 23154 17118
rect 16818 17054 16830 17106
rect 16882 17054 16894 17106
rect 11678 17042 11730 17054
rect 23102 17042 23154 17054
rect 24334 17106 24386 17118
rect 24334 17042 24386 17054
rect 25342 17106 25394 17118
rect 25342 17042 25394 17054
rect 27246 17106 27298 17118
rect 27246 17042 27298 17054
rect 27582 17106 27634 17118
rect 27582 17042 27634 17054
rect 28814 17106 28866 17118
rect 28814 17042 28866 17054
rect 30382 17106 30434 17118
rect 30382 17042 30434 17054
rect 34526 17106 34578 17118
rect 34526 17042 34578 17054
rect 39342 17106 39394 17118
rect 39342 17042 39394 17054
rect 40238 17106 40290 17118
rect 53342 17106 53394 17118
rect 59950 17106 60002 17118
rect 72606 17106 72658 17118
rect 41458 17054 41470 17106
rect 41522 17054 41534 17106
rect 54674 17054 54686 17106
rect 54738 17054 54750 17106
rect 55458 17054 55470 17106
rect 55522 17054 55534 17106
rect 56914 17054 56926 17106
rect 56978 17054 56990 17106
rect 71362 17054 71374 17106
rect 71426 17054 71438 17106
rect 40238 17042 40290 17054
rect 53342 17042 53394 17054
rect 59950 17042 60002 17054
rect 72606 17042 72658 17054
rect 4846 16994 4898 17006
rect 16270 16994 16322 17006
rect 24446 16994 24498 17006
rect 6850 16942 6862 16994
rect 6914 16942 6926 16994
rect 23314 16942 23326 16994
rect 23378 16942 23390 16994
rect 4846 16930 4898 16942
rect 16270 16930 16322 16942
rect 24446 16930 24498 16942
rect 25790 16994 25842 17006
rect 34750 16994 34802 17006
rect 28466 16942 28478 16994
rect 28530 16942 28542 16994
rect 25790 16930 25842 16942
rect 34750 16930 34802 16942
rect 39678 16994 39730 17006
rect 39678 16930 39730 16942
rect 41022 16994 41074 17006
rect 41022 16930 41074 16942
rect 42030 16994 42082 17006
rect 42030 16930 42082 16942
rect 42478 16994 42530 17006
rect 42478 16930 42530 16942
rect 43038 16994 43090 17006
rect 47966 16994 48018 17006
rect 56814 16994 56866 17006
rect 68910 16994 68962 17006
rect 46050 16942 46062 16994
rect 46114 16942 46126 16994
rect 50754 16942 50766 16994
rect 50818 16942 50830 16994
rect 55794 16942 55806 16994
rect 55858 16942 55870 16994
rect 57586 16942 57598 16994
rect 57650 16942 57662 16994
rect 63074 16942 63086 16994
rect 63138 16942 63150 16994
rect 67554 16942 67566 16994
rect 67618 16942 67630 16994
rect 43038 16930 43090 16942
rect 47966 16930 48018 16942
rect 56814 16930 56866 16942
rect 68910 16930 68962 16942
rect 69806 16994 69858 17006
rect 71486 16994 71538 17006
rect 70466 16942 70478 16994
rect 70530 16942 70542 16994
rect 69806 16930 69858 16942
rect 71486 16930 71538 16942
rect 72270 16994 72322 17006
rect 77074 16942 77086 16994
rect 77138 16942 77150 16994
rect 72270 16930 72322 16942
rect 10558 16882 10610 16894
rect 3938 16830 3950 16882
rect 4002 16830 4014 16882
rect 6178 16830 6190 16882
rect 6242 16830 6254 16882
rect 10322 16830 10334 16882
rect 10386 16830 10398 16882
rect 10558 16818 10610 16830
rect 10894 16882 10946 16894
rect 11342 16882 11394 16894
rect 11106 16830 11118 16882
rect 11170 16830 11182 16882
rect 10894 16818 10946 16830
rect 11342 16818 11394 16830
rect 11566 16882 11618 16894
rect 11566 16818 11618 16830
rect 11902 16882 11954 16894
rect 15598 16882 15650 16894
rect 15250 16830 15262 16882
rect 15314 16830 15326 16882
rect 11902 16818 11954 16830
rect 15598 16818 15650 16830
rect 16158 16882 16210 16894
rect 16158 16818 16210 16830
rect 16382 16882 16434 16894
rect 16382 16818 16434 16830
rect 17614 16882 17666 16894
rect 17614 16818 17666 16830
rect 19182 16882 19234 16894
rect 19182 16818 19234 16830
rect 19854 16882 19906 16894
rect 19854 16818 19906 16830
rect 20414 16882 20466 16894
rect 20414 16818 20466 16830
rect 23662 16882 23714 16894
rect 23662 16818 23714 16830
rect 24110 16882 24162 16894
rect 24110 16818 24162 16830
rect 26686 16882 26738 16894
rect 26686 16818 26738 16830
rect 30606 16882 30658 16894
rect 30606 16818 30658 16830
rect 32510 16882 32562 16894
rect 32510 16818 32562 16830
rect 33070 16882 33122 16894
rect 42366 16882 42418 16894
rect 47406 16882 47458 16894
rect 33506 16830 33518 16882
rect 33570 16830 33582 16882
rect 35634 16830 35646 16882
rect 35698 16830 35710 16882
rect 37202 16830 37214 16882
rect 37266 16830 37278 16882
rect 38546 16830 38558 16882
rect 38610 16830 38622 16882
rect 41794 16830 41806 16882
rect 41858 16830 41870 16882
rect 42914 16830 42926 16882
rect 42978 16830 42990 16882
rect 43586 16830 43598 16882
rect 43650 16830 43662 16882
rect 44146 16830 44158 16882
rect 44210 16830 44222 16882
rect 44930 16830 44942 16882
rect 44994 16830 45006 16882
rect 46946 16830 46958 16882
rect 47010 16830 47022 16882
rect 33070 16818 33122 16830
rect 42366 16818 42418 16830
rect 47406 16818 47458 16830
rect 48974 16882 49026 16894
rect 54350 16882 54402 16894
rect 58494 16882 58546 16894
rect 50082 16830 50094 16882
rect 50146 16830 50158 16882
rect 55122 16830 55134 16882
rect 55186 16830 55198 16882
rect 55458 16830 55470 16882
rect 55522 16830 55534 16882
rect 56578 16830 56590 16882
rect 56642 16830 56654 16882
rect 57474 16830 57486 16882
rect 57538 16830 57550 16882
rect 48974 16818 49026 16830
rect 54350 16818 54402 16830
rect 58494 16818 58546 16830
rect 59726 16882 59778 16894
rect 65550 16882 65602 16894
rect 60162 16830 60174 16882
rect 60226 16830 60238 16882
rect 63858 16830 63870 16882
rect 63922 16830 63934 16882
rect 59726 16818 59778 16830
rect 65550 16818 65602 16830
rect 65886 16882 65938 16894
rect 65886 16818 65938 16830
rect 66446 16882 66498 16894
rect 68350 16882 68402 16894
rect 66770 16830 66782 16882
rect 66834 16830 66846 16882
rect 66446 16818 66498 16830
rect 68350 16818 68402 16830
rect 69246 16882 69298 16894
rect 70690 16830 70702 16882
rect 70754 16830 70766 16882
rect 71698 16830 71710 16882
rect 71762 16830 71774 16882
rect 77858 16830 77870 16882
rect 77922 16830 77934 16882
rect 69246 16818 69298 16830
rect 15710 16770 15762 16782
rect 18846 16770 18898 16782
rect 44382 16770 44434 16782
rect 8978 16718 8990 16770
rect 9042 16718 9054 16770
rect 12338 16718 12350 16770
rect 12402 16718 12414 16770
rect 14466 16718 14478 16770
rect 14530 16718 14542 16770
rect 18050 16718 18062 16770
rect 18114 16718 18126 16770
rect 28018 16718 28030 16770
rect 28082 16718 28094 16770
rect 29922 16718 29934 16770
rect 29986 16718 29998 16770
rect 32050 16718 32062 16770
rect 32114 16718 32126 16770
rect 34402 16718 34414 16770
rect 34466 16718 34478 16770
rect 35522 16718 35534 16770
rect 35586 16718 35598 16770
rect 15710 16706 15762 16718
rect 18846 16706 18898 16718
rect 44382 16706 44434 16718
rect 46510 16770 46562 16782
rect 52882 16718 52894 16770
rect 52946 16718 52958 16770
rect 60946 16718 60958 16770
rect 61010 16718 61022 16770
rect 74946 16718 74958 16770
rect 75010 16718 75022 16770
rect 46510 16706 46562 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 12014 16658 12066 16670
rect 12014 16594 12066 16606
rect 19294 16658 19346 16670
rect 30830 16658 30882 16670
rect 25554 16606 25566 16658
rect 25618 16655 25630 16658
rect 25778 16655 25790 16658
rect 25618 16609 25790 16655
rect 25618 16606 25630 16609
rect 25778 16606 25790 16609
rect 25842 16606 25854 16658
rect 32274 16606 32286 16658
rect 32338 16606 32350 16658
rect 35410 16606 35422 16658
rect 35474 16606 35486 16658
rect 39218 16606 39230 16658
rect 39282 16655 39294 16658
rect 39666 16655 39678 16658
rect 39282 16609 39678 16655
rect 39282 16606 39294 16609
rect 39666 16606 39678 16609
rect 39730 16606 39742 16658
rect 19294 16594 19346 16606
rect 30830 16594 30882 16606
rect 1344 16490 78624 16524
rect 1344 16438 10874 16490
rect 10926 16438 10978 16490
rect 11030 16438 11082 16490
rect 11134 16438 30194 16490
rect 30246 16438 30298 16490
rect 30350 16438 30402 16490
rect 30454 16438 49514 16490
rect 49566 16438 49618 16490
rect 49670 16438 49722 16490
rect 49774 16438 68834 16490
rect 68886 16438 68938 16490
rect 68990 16438 69042 16490
rect 69094 16438 78624 16490
rect 1344 16404 78624 16438
rect 7758 16322 7810 16334
rect 32734 16322 32786 16334
rect 18722 16270 18734 16322
rect 18786 16270 18798 16322
rect 7758 16258 7810 16270
rect 32734 16258 32786 16270
rect 32958 16322 33010 16334
rect 32958 16258 33010 16270
rect 33406 16322 33458 16334
rect 67566 16322 67618 16334
rect 40226 16270 40238 16322
rect 40290 16270 40302 16322
rect 33406 16258 33458 16270
rect 67566 16258 67618 16270
rect 69134 16322 69186 16334
rect 69134 16258 69186 16270
rect 9438 16210 9490 16222
rect 9438 16146 9490 16158
rect 10334 16210 10386 16222
rect 10334 16146 10386 16158
rect 12686 16210 12738 16222
rect 12686 16146 12738 16158
rect 13582 16210 13634 16222
rect 13582 16146 13634 16158
rect 14590 16210 14642 16222
rect 16830 16210 16882 16222
rect 16146 16158 16158 16210
rect 16210 16158 16222 16210
rect 14590 16146 14642 16158
rect 16830 16146 16882 16158
rect 17502 16210 17554 16222
rect 34302 16210 34354 16222
rect 41806 16210 41858 16222
rect 48190 16210 48242 16222
rect 22082 16158 22094 16210
rect 22146 16158 22158 16210
rect 29362 16158 29374 16210
rect 29426 16158 29438 16210
rect 41122 16158 41134 16210
rect 41186 16158 41198 16210
rect 45826 16158 45838 16210
rect 45890 16158 45902 16210
rect 46834 16158 46846 16210
rect 46898 16158 46910 16210
rect 17502 16146 17554 16158
rect 34302 16146 34354 16158
rect 41806 16146 41858 16158
rect 48190 16146 48242 16158
rect 51550 16210 51602 16222
rect 51550 16146 51602 16158
rect 55918 16210 55970 16222
rect 58942 16210 58994 16222
rect 58370 16158 58382 16210
rect 58434 16158 58446 16210
rect 55918 16146 55970 16158
rect 58942 16146 58994 16158
rect 59390 16210 59442 16222
rect 59390 16146 59442 16158
rect 66222 16210 66274 16222
rect 66222 16146 66274 16158
rect 69582 16210 69634 16222
rect 69582 16146 69634 16158
rect 76414 16210 76466 16222
rect 76414 16146 76466 16158
rect 3726 16098 3778 16110
rect 3726 16034 3778 16046
rect 8094 16098 8146 16110
rect 15934 16098 15986 16110
rect 8530 16046 8542 16098
rect 8594 16046 8606 16098
rect 11106 16046 11118 16098
rect 11170 16046 11182 16098
rect 15698 16046 15710 16098
rect 15762 16046 15774 16098
rect 8094 16034 8146 16046
rect 15934 16034 15986 16046
rect 17054 16098 17106 16110
rect 17054 16034 17106 16046
rect 17838 16098 17890 16110
rect 17838 16034 17890 16046
rect 18958 16098 19010 16110
rect 26462 16098 26514 16110
rect 32510 16098 32562 16110
rect 38894 16098 38946 16110
rect 42478 16098 42530 16110
rect 43486 16098 43538 16110
rect 47630 16098 47682 16110
rect 50990 16098 51042 16110
rect 57934 16098 57986 16110
rect 73838 16098 73890 16110
rect 24994 16046 25006 16098
rect 25058 16046 25070 16098
rect 29922 16046 29934 16098
rect 29986 16046 29998 16098
rect 31042 16046 31054 16098
rect 31106 16046 31118 16098
rect 35858 16046 35870 16098
rect 35922 16046 35934 16098
rect 36978 16046 36990 16098
rect 37042 16046 37054 16098
rect 38210 16046 38222 16098
rect 38274 16046 38286 16098
rect 39106 16046 39118 16098
rect 39170 16046 39182 16098
rect 41234 16046 41246 16098
rect 41298 16046 41310 16098
rect 43026 16046 43038 16098
rect 43090 16046 43102 16098
rect 43810 16046 43822 16098
rect 43874 16046 43886 16098
rect 44818 16046 44830 16098
rect 44882 16046 44894 16098
rect 48850 16046 48862 16098
rect 48914 16046 48926 16098
rect 53666 16046 53678 16098
rect 53730 16046 53742 16098
rect 54002 16046 54014 16098
rect 54066 16046 54078 16098
rect 54338 16046 54350 16098
rect 54402 16046 54414 16098
rect 54674 16046 54686 16098
rect 54738 16046 54750 16098
rect 57250 16046 57262 16098
rect 57314 16046 57326 16098
rect 68450 16046 68462 16098
rect 68514 16046 68526 16098
rect 74386 16046 74398 16098
rect 74450 16046 74462 16098
rect 76962 16046 76974 16098
rect 77026 16046 77038 16098
rect 18958 16034 19010 16046
rect 26462 16034 26514 16046
rect 32510 16034 32562 16046
rect 38894 16034 38946 16046
rect 42478 16034 42530 16046
rect 43486 16034 43538 16046
rect 47630 16034 47682 16046
rect 50990 16034 51042 16046
rect 57934 16034 57986 16046
rect 73838 16034 73890 16046
rect 3390 15986 3442 15998
rect 3390 15922 3442 15934
rect 4398 15986 4450 15998
rect 12238 15986 12290 15998
rect 8866 15934 8878 15986
rect 8930 15934 8942 15986
rect 11330 15934 11342 15986
rect 11394 15934 11406 15986
rect 11554 15934 11566 15986
rect 11618 15934 11630 15986
rect 4398 15922 4450 15934
rect 12238 15922 12290 15934
rect 14478 15986 14530 15998
rect 14478 15922 14530 15934
rect 15262 15986 15314 15998
rect 15262 15922 15314 15934
rect 16158 15986 16210 15998
rect 27022 15986 27074 15998
rect 19842 15934 19854 15986
rect 19906 15934 19918 15986
rect 24210 15934 24222 15986
rect 24274 15934 24286 15986
rect 16158 15922 16210 15934
rect 27022 15922 27074 15934
rect 27470 15986 27522 15998
rect 32286 15986 32338 15998
rect 44046 15986 44098 15998
rect 30258 15934 30270 15986
rect 30322 15934 30334 15986
rect 31378 15934 31390 15986
rect 31442 15934 31454 15986
rect 31714 15934 31726 15986
rect 31778 15934 31790 15986
rect 36418 15934 36430 15986
rect 36482 15934 36494 15986
rect 42130 15934 42142 15986
rect 42194 15934 42206 15986
rect 27470 15922 27522 15934
rect 32286 15922 32338 15934
rect 44046 15922 44098 15934
rect 49310 15986 49362 15998
rect 49310 15922 49362 15934
rect 52222 15986 52274 15998
rect 56130 15934 56142 15986
rect 56194 15934 56206 15986
rect 66546 15934 66558 15986
rect 66610 15934 66622 15986
rect 52222 15922 52274 15934
rect 4062 15874 4114 15886
rect 4062 15810 4114 15822
rect 10446 15874 10498 15886
rect 10446 15810 10498 15822
rect 14254 15874 14306 15886
rect 14254 15810 14306 15822
rect 14702 15874 14754 15886
rect 14702 15810 14754 15822
rect 14926 15874 14978 15886
rect 14926 15810 14978 15822
rect 15150 15874 15202 15886
rect 15150 15810 15202 15822
rect 16270 15874 16322 15886
rect 16270 15810 16322 15822
rect 20190 15874 20242 15886
rect 20190 15810 20242 15822
rect 20638 15874 20690 15886
rect 44158 15874 44210 15886
rect 35970 15822 35982 15874
rect 36034 15822 36046 15874
rect 42802 15822 42814 15874
rect 42866 15822 42878 15874
rect 20638 15810 20690 15822
rect 44158 15810 44210 15822
rect 46398 15874 46450 15886
rect 46398 15810 46450 15822
rect 64990 15874 65042 15886
rect 64990 15810 65042 15822
rect 65438 15874 65490 15886
rect 65438 15810 65490 15822
rect 65662 15874 65714 15886
rect 76750 15874 76802 15886
rect 74162 15822 74174 15874
rect 74226 15822 74238 15874
rect 65662 15810 65714 15822
rect 76750 15810 76802 15822
rect 1344 15706 78784 15740
rect 1344 15654 20534 15706
rect 20586 15654 20638 15706
rect 20690 15654 20742 15706
rect 20794 15654 39854 15706
rect 39906 15654 39958 15706
rect 40010 15654 40062 15706
rect 40114 15654 59174 15706
rect 59226 15654 59278 15706
rect 59330 15654 59382 15706
rect 59434 15654 78494 15706
rect 78546 15654 78598 15706
rect 78650 15654 78702 15706
rect 78754 15654 78784 15706
rect 1344 15620 78784 15654
rect 5294 15538 5346 15550
rect 5294 15474 5346 15486
rect 7646 15538 7698 15550
rect 7646 15474 7698 15486
rect 21758 15538 21810 15550
rect 21758 15474 21810 15486
rect 22206 15538 22258 15550
rect 22206 15474 22258 15486
rect 23438 15538 23490 15550
rect 23438 15474 23490 15486
rect 26686 15538 26738 15550
rect 26686 15474 26738 15486
rect 30830 15538 30882 15550
rect 30830 15474 30882 15486
rect 31278 15538 31330 15550
rect 31278 15474 31330 15486
rect 32286 15538 32338 15550
rect 32286 15474 32338 15486
rect 32958 15538 33010 15550
rect 32958 15474 33010 15486
rect 33854 15538 33906 15550
rect 33854 15474 33906 15486
rect 34526 15538 34578 15550
rect 35198 15538 35250 15550
rect 34850 15486 34862 15538
rect 34914 15486 34926 15538
rect 34526 15474 34578 15486
rect 35198 15474 35250 15486
rect 39230 15538 39282 15550
rect 39230 15474 39282 15486
rect 43486 15538 43538 15550
rect 43486 15474 43538 15486
rect 43598 15538 43650 15550
rect 43598 15474 43650 15486
rect 44158 15538 44210 15550
rect 44158 15474 44210 15486
rect 44382 15538 44434 15550
rect 44382 15474 44434 15486
rect 46062 15538 46114 15550
rect 50990 15538 51042 15550
rect 48850 15486 48862 15538
rect 48914 15486 48926 15538
rect 49074 15486 49086 15538
rect 49138 15486 49150 15538
rect 46062 15474 46114 15486
rect 50990 15474 51042 15486
rect 52558 15538 52610 15550
rect 52558 15474 52610 15486
rect 54798 15538 54850 15550
rect 54798 15474 54850 15486
rect 55134 15538 55186 15550
rect 55134 15474 55186 15486
rect 56590 15538 56642 15550
rect 57262 15538 57314 15550
rect 56914 15486 56926 15538
rect 56978 15486 56990 15538
rect 56590 15474 56642 15486
rect 57262 15474 57314 15486
rect 58046 15538 58098 15550
rect 58046 15474 58098 15486
rect 63870 15538 63922 15550
rect 63870 15474 63922 15486
rect 67566 15538 67618 15550
rect 67566 15474 67618 15486
rect 68238 15538 68290 15550
rect 68238 15474 68290 15486
rect 68686 15538 68738 15550
rect 68686 15474 68738 15486
rect 69134 15538 69186 15550
rect 69134 15474 69186 15486
rect 16158 15426 16210 15438
rect 2706 15374 2718 15426
rect 2770 15374 2782 15426
rect 5954 15374 5966 15426
rect 6018 15374 6030 15426
rect 6402 15374 6414 15426
rect 6466 15374 6478 15426
rect 6850 15374 6862 15426
rect 6914 15374 6926 15426
rect 16158 15362 16210 15374
rect 17390 15426 17442 15438
rect 17390 15362 17442 15374
rect 24446 15426 24498 15438
rect 32062 15426 32114 15438
rect 29698 15374 29710 15426
rect 29762 15374 29774 15426
rect 24446 15362 24498 15374
rect 32062 15362 32114 15374
rect 32510 15426 32562 15438
rect 32510 15362 32562 15374
rect 33182 15426 33234 15438
rect 33182 15362 33234 15374
rect 33630 15426 33682 15438
rect 33630 15362 33682 15374
rect 34078 15426 34130 15438
rect 42702 15426 42754 15438
rect 64654 15426 64706 15438
rect 70030 15426 70082 15438
rect 36754 15374 36766 15426
rect 36818 15374 36830 15426
rect 50082 15374 50094 15426
rect 50146 15374 50158 15426
rect 55458 15374 55470 15426
rect 55522 15374 55534 15426
rect 57586 15374 57598 15426
rect 57650 15374 57662 15426
rect 59266 15374 59278 15426
rect 59330 15374 59342 15426
rect 65202 15374 65214 15426
rect 65266 15374 65278 15426
rect 65538 15374 65550 15426
rect 65602 15374 65614 15426
rect 66770 15374 66782 15426
rect 66834 15374 66846 15426
rect 74498 15374 74510 15426
rect 74562 15374 74574 15426
rect 34078 15362 34130 15374
rect 42702 15362 42754 15374
rect 64654 15362 64706 15374
rect 70030 15362 70082 15374
rect 5630 15314 5682 15326
rect 2034 15262 2046 15314
rect 2098 15262 2110 15314
rect 5630 15250 5682 15262
rect 7198 15314 7250 15326
rect 17950 15314 18002 15326
rect 11554 15262 11566 15314
rect 11618 15262 11630 15314
rect 12786 15262 12798 15314
rect 12850 15262 12862 15314
rect 13122 15262 13134 15314
rect 13186 15262 13198 15314
rect 14578 15262 14590 15314
rect 14642 15262 14654 15314
rect 17602 15262 17614 15314
rect 17666 15262 17678 15314
rect 7198 15250 7250 15262
rect 17950 15250 18002 15262
rect 18286 15314 18338 15326
rect 18286 15250 18338 15262
rect 18622 15314 18674 15326
rect 23662 15314 23714 15326
rect 21522 15262 21534 15314
rect 21586 15262 21598 15314
rect 18622 15250 18674 15262
rect 23662 15250 23714 15262
rect 24110 15314 24162 15326
rect 24110 15250 24162 15262
rect 24558 15314 24610 15326
rect 24558 15250 24610 15262
rect 25342 15314 25394 15326
rect 25342 15250 25394 15262
rect 25566 15314 25618 15326
rect 25566 15250 25618 15262
rect 25790 15314 25842 15326
rect 25790 15250 25842 15262
rect 26350 15314 26402 15326
rect 26350 15250 26402 15262
rect 26462 15314 26514 15326
rect 26462 15250 26514 15262
rect 28142 15314 28194 15326
rect 31726 15314 31778 15326
rect 29586 15262 29598 15314
rect 29650 15262 29662 15314
rect 28142 15250 28194 15262
rect 31726 15250 31778 15262
rect 33294 15314 33346 15326
rect 33294 15250 33346 15262
rect 35758 15314 35810 15326
rect 40014 15314 40066 15326
rect 40910 15314 40962 15326
rect 43710 15314 43762 15326
rect 36642 15262 36654 15314
rect 36706 15262 36718 15314
rect 37426 15262 37438 15314
rect 37490 15262 37502 15314
rect 40226 15262 40238 15314
rect 40290 15262 40302 15314
rect 41122 15262 41134 15314
rect 41186 15262 41198 15314
rect 35758 15250 35810 15262
rect 40014 15250 40066 15262
rect 40910 15250 40962 15262
rect 43710 15250 43762 15262
rect 44046 15314 44098 15326
rect 56030 15314 56082 15326
rect 64766 15314 64818 15326
rect 73950 15314 74002 15326
rect 44706 15262 44718 15314
rect 44770 15262 44782 15314
rect 47730 15262 47742 15314
rect 47794 15262 47806 15314
rect 48738 15262 48750 15314
rect 48802 15262 48814 15314
rect 49634 15262 49646 15314
rect 49698 15262 49710 15314
rect 51426 15262 51438 15314
rect 51490 15262 51502 15314
rect 59714 15262 59726 15314
rect 59778 15262 59790 15314
rect 60274 15262 60286 15314
rect 60338 15262 60350 15314
rect 66322 15262 66334 15314
rect 66386 15262 66398 15314
rect 67218 15262 67230 15314
rect 67282 15262 67294 15314
rect 69794 15262 69806 15314
rect 69858 15262 69870 15314
rect 74386 15262 74398 15314
rect 74450 15262 74462 15314
rect 76066 15262 76078 15314
rect 76130 15262 76142 15314
rect 44046 15250 44098 15262
rect 56030 15250 56082 15262
rect 64766 15250 64818 15262
rect 73950 15250 74002 15262
rect 16606 15202 16658 15214
rect 4834 15150 4846 15202
rect 4898 15150 4910 15202
rect 14690 15150 14702 15202
rect 14754 15150 14766 15202
rect 16606 15138 16658 15150
rect 18398 15202 18450 15214
rect 23550 15202 23602 15214
rect 19170 15150 19182 15202
rect 19234 15150 19246 15202
rect 18398 15138 18450 15150
rect 23550 15138 23602 15150
rect 27134 15202 27186 15214
rect 27134 15138 27186 15150
rect 27582 15202 27634 15214
rect 27582 15138 27634 15150
rect 35534 15202 35586 15214
rect 40350 15202 40402 15214
rect 36754 15150 36766 15202
rect 36818 15150 36830 15202
rect 38210 15150 38222 15202
rect 38274 15150 38286 15202
rect 35534 15138 35586 15150
rect 40350 15138 40402 15150
rect 45166 15202 45218 15214
rect 48190 15202 48242 15214
rect 53006 15202 53058 15214
rect 73166 15202 73218 15214
rect 45602 15150 45614 15202
rect 45666 15150 45678 15202
rect 51762 15150 51774 15202
rect 51826 15150 51838 15202
rect 59602 15150 59614 15202
rect 59666 15150 59678 15202
rect 66882 15150 66894 15202
rect 66946 15150 66958 15202
rect 45166 15138 45218 15150
rect 48190 15138 48242 15150
rect 53006 15138 53058 15150
rect 73166 15138 73218 15150
rect 77982 15202 78034 15214
rect 77982 15138 78034 15150
rect 17726 15090 17778 15102
rect 15026 15038 15038 15090
rect 15090 15038 15102 15090
rect 15922 15038 15934 15090
rect 15986 15087 15998 15090
rect 16482 15087 16494 15090
rect 15986 15041 16494 15087
rect 15986 15038 15998 15041
rect 16482 15038 16494 15041
rect 16546 15038 16558 15090
rect 17726 15026 17778 15038
rect 26014 15090 26066 15102
rect 32174 15090 32226 15102
rect 28578 15038 28590 15090
rect 28642 15038 28654 15090
rect 26014 15026 26066 15038
rect 32174 15026 32226 15038
rect 33742 15090 33794 15102
rect 73614 15090 73666 15102
rect 36082 15038 36094 15090
rect 36146 15038 36158 15090
rect 33742 15026 33794 15038
rect 73614 15026 73666 15038
rect 1344 14922 78624 14956
rect 1344 14870 10874 14922
rect 10926 14870 10978 14922
rect 11030 14870 11082 14922
rect 11134 14870 30194 14922
rect 30246 14870 30298 14922
rect 30350 14870 30402 14922
rect 30454 14870 49514 14922
rect 49566 14870 49618 14922
rect 49670 14870 49722 14922
rect 49774 14870 68834 14922
rect 68886 14870 68938 14922
rect 68990 14870 69042 14922
rect 69094 14870 78624 14922
rect 1344 14836 78624 14870
rect 38558 14754 38610 14766
rect 26898 14702 26910 14754
rect 26962 14751 26974 14754
rect 27346 14751 27358 14754
rect 26962 14705 27358 14751
rect 26962 14702 26974 14705
rect 27346 14702 27358 14705
rect 27410 14702 27422 14754
rect 38558 14690 38610 14702
rect 57262 14754 57314 14766
rect 57262 14690 57314 14702
rect 1934 14642 1986 14654
rect 18286 14642 18338 14654
rect 13906 14590 13918 14642
rect 13970 14590 13982 14642
rect 17154 14590 17166 14642
rect 17218 14590 17230 14642
rect 1934 14578 1986 14590
rect 18286 14578 18338 14590
rect 22094 14642 22146 14654
rect 22094 14578 22146 14590
rect 26910 14642 26962 14654
rect 37998 14642 38050 14654
rect 42030 14642 42082 14654
rect 32722 14590 32734 14642
rect 32786 14590 32798 14642
rect 37650 14590 37662 14642
rect 37714 14590 37726 14642
rect 40898 14590 40910 14642
rect 40962 14590 40974 14642
rect 26910 14578 26962 14590
rect 37998 14578 38050 14590
rect 42030 14578 42082 14590
rect 49198 14642 49250 14654
rect 49198 14578 49250 14590
rect 51662 14642 51714 14654
rect 51662 14578 51714 14590
rect 54350 14642 54402 14654
rect 54350 14578 54402 14590
rect 56142 14642 56194 14654
rect 59266 14590 59278 14642
rect 59330 14590 59342 14642
rect 64418 14590 64430 14642
rect 64482 14590 64494 14642
rect 65986 14590 65998 14642
rect 66050 14590 66062 14642
rect 68898 14590 68910 14642
rect 68962 14590 68974 14642
rect 71026 14590 71038 14642
rect 71090 14590 71102 14642
rect 56142 14578 56194 14590
rect 6078 14530 6130 14542
rect 18622 14530 18674 14542
rect 4274 14478 4286 14530
rect 4338 14478 4350 14530
rect 6850 14478 6862 14530
rect 6914 14478 6926 14530
rect 14690 14478 14702 14530
rect 14754 14478 14766 14530
rect 16706 14478 16718 14530
rect 16770 14478 16782 14530
rect 17378 14478 17390 14530
rect 17442 14478 17454 14530
rect 18386 14478 18398 14530
rect 18450 14478 18462 14530
rect 6078 14466 6130 14478
rect 18622 14466 18674 14478
rect 18958 14530 19010 14542
rect 27918 14530 27970 14542
rect 21522 14478 21534 14530
rect 21586 14478 21598 14530
rect 18958 14466 19010 14478
rect 27918 14466 27970 14478
rect 28590 14530 28642 14542
rect 28590 14466 28642 14478
rect 29150 14530 29202 14542
rect 29150 14466 29202 14478
rect 29710 14530 29762 14542
rect 35646 14530 35698 14542
rect 30258 14478 30270 14530
rect 30322 14478 30334 14530
rect 31266 14478 31278 14530
rect 31330 14478 31342 14530
rect 32386 14478 32398 14530
rect 32450 14478 32462 14530
rect 33618 14478 33630 14530
rect 33682 14478 33694 14530
rect 34626 14478 34638 14530
rect 34690 14478 34702 14530
rect 29710 14466 29762 14478
rect 35646 14466 35698 14478
rect 36206 14530 36258 14542
rect 38334 14530 38386 14542
rect 37426 14478 37438 14530
rect 37490 14478 37502 14530
rect 36206 14466 36258 14478
rect 38334 14466 38386 14478
rect 39678 14530 39730 14542
rect 51102 14530 51154 14542
rect 39890 14478 39902 14530
rect 39954 14478 39966 14530
rect 41010 14478 41022 14530
rect 41074 14478 41086 14530
rect 46946 14478 46958 14530
rect 47010 14478 47022 14530
rect 48290 14478 48302 14530
rect 48354 14478 48366 14530
rect 50306 14478 50318 14530
rect 50370 14478 50382 14530
rect 39678 14466 39730 14478
rect 51102 14466 51154 14478
rect 52110 14530 52162 14542
rect 54686 14530 54738 14542
rect 52882 14478 52894 14530
rect 52946 14478 52958 14530
rect 52110 14466 52162 14478
rect 54686 14466 54738 14478
rect 55246 14530 55298 14542
rect 55246 14466 55298 14478
rect 56590 14530 56642 14542
rect 56590 14466 56642 14478
rect 56702 14530 56754 14542
rect 56702 14466 56754 14478
rect 57038 14530 57090 14542
rect 57038 14466 57090 14478
rect 57374 14530 57426 14542
rect 59614 14530 59666 14542
rect 57922 14478 57934 14530
rect 57986 14478 57998 14530
rect 58818 14478 58830 14530
rect 58882 14478 58894 14530
rect 57374 14466 57426 14478
rect 59614 14466 59666 14478
rect 63982 14530 64034 14542
rect 63982 14466 64034 14478
rect 64094 14530 64146 14542
rect 76190 14530 76242 14542
rect 64530 14478 64542 14530
rect 64594 14478 64606 14530
rect 66098 14478 66110 14530
rect 66162 14478 66174 14530
rect 66882 14478 66894 14530
rect 66946 14478 66958 14530
rect 71810 14478 71822 14530
rect 71874 14478 71886 14530
rect 75618 14478 75630 14530
rect 75682 14478 75694 14530
rect 64094 14466 64146 14478
rect 76190 14466 76242 14478
rect 7870 14418 7922 14430
rect 6738 14366 6750 14418
rect 6802 14366 6814 14418
rect 7870 14354 7922 14366
rect 18846 14418 18898 14430
rect 18846 14354 18898 14366
rect 41582 14418 41634 14430
rect 56926 14418 56978 14430
rect 59838 14418 59890 14430
rect 76862 14418 76914 14430
rect 47506 14366 47518 14418
rect 47570 14366 47582 14418
rect 50754 14366 50766 14418
rect 50818 14366 50830 14418
rect 53778 14366 53790 14418
rect 53842 14366 53854 14418
rect 57586 14366 57598 14418
rect 57650 14366 57662 14418
rect 65874 14366 65886 14418
rect 65938 14366 65950 14418
rect 41582 14354 41634 14366
rect 56926 14354 56978 14366
rect 59838 14354 59890 14366
rect 76862 14354 76914 14366
rect 77198 14418 77250 14430
rect 77198 14354 77250 14366
rect 77646 14418 77698 14430
rect 77646 14354 77698 14366
rect 4846 14306 4898 14318
rect 4846 14242 4898 14254
rect 5742 14306 5794 14318
rect 5742 14242 5794 14254
rect 7534 14306 7586 14318
rect 7534 14242 7586 14254
rect 12350 14306 12402 14318
rect 12350 14242 12402 14254
rect 15150 14306 15202 14318
rect 15150 14242 15202 14254
rect 16942 14306 16994 14318
rect 16942 14242 16994 14254
rect 17166 14306 17218 14318
rect 17166 14242 17218 14254
rect 17950 14306 18002 14318
rect 17950 14242 18002 14254
rect 18174 14306 18226 14318
rect 39790 14306 39842 14318
rect 21298 14254 21310 14306
rect 21362 14254 21374 14306
rect 27570 14254 27582 14306
rect 27634 14254 27646 14306
rect 38882 14254 38894 14306
rect 38946 14254 38958 14306
rect 18174 14242 18226 14254
rect 39790 14242 39842 14254
rect 42590 14306 42642 14318
rect 42590 14242 42642 14254
rect 55582 14306 55634 14318
rect 55582 14242 55634 14254
rect 59278 14306 59330 14318
rect 59278 14242 59330 14254
rect 59390 14306 59442 14318
rect 59390 14242 59442 14254
rect 63534 14306 63586 14318
rect 63534 14242 63586 14254
rect 64318 14306 64370 14318
rect 64318 14242 64370 14254
rect 72270 14306 72322 14318
rect 72270 14242 72322 14254
rect 74622 14306 74674 14318
rect 74622 14242 74674 14254
rect 76526 14306 76578 14318
rect 76526 14242 76578 14254
rect 1344 14138 78784 14172
rect 1344 14086 20534 14138
rect 20586 14086 20638 14138
rect 20690 14086 20742 14138
rect 20794 14086 39854 14138
rect 39906 14086 39958 14138
rect 40010 14086 40062 14138
rect 40114 14086 59174 14138
rect 59226 14086 59278 14138
rect 59330 14086 59382 14138
rect 59434 14086 78494 14138
rect 78546 14086 78598 14138
rect 78650 14086 78702 14138
rect 78754 14086 78784 14138
rect 1344 14052 78784 14086
rect 11902 13970 11954 13982
rect 11902 13906 11954 13918
rect 13022 13970 13074 13982
rect 17838 13970 17890 13982
rect 16482 13918 16494 13970
rect 16546 13918 16558 13970
rect 13022 13906 13074 13918
rect 17838 13906 17890 13918
rect 24334 13970 24386 13982
rect 24334 13906 24386 13918
rect 25454 13970 25506 13982
rect 25454 13906 25506 13918
rect 30046 13970 30098 13982
rect 30046 13906 30098 13918
rect 33406 13970 33458 13982
rect 33406 13906 33458 13918
rect 34190 13970 34242 13982
rect 34190 13906 34242 13918
rect 34862 13970 34914 13982
rect 34862 13906 34914 13918
rect 37550 13970 37602 13982
rect 37550 13906 37602 13918
rect 39230 13970 39282 13982
rect 39230 13906 39282 13918
rect 43038 13970 43090 13982
rect 43038 13906 43090 13918
rect 46398 13970 46450 13982
rect 47966 13970 48018 13982
rect 47842 13918 47854 13970
rect 47906 13918 47918 13970
rect 46398 13906 46450 13918
rect 47966 13906 48018 13918
rect 52894 13970 52946 13982
rect 56142 13970 56194 13982
rect 63310 13970 63362 13982
rect 55570 13918 55582 13970
rect 55634 13918 55646 13970
rect 59714 13918 59726 13970
rect 59778 13918 59790 13970
rect 52894 13906 52946 13918
rect 56142 13906 56194 13918
rect 63310 13906 63362 13918
rect 63534 13970 63586 13982
rect 63534 13906 63586 13918
rect 63646 13970 63698 13982
rect 70030 13970 70082 13982
rect 66098 13918 66110 13970
rect 66162 13918 66174 13970
rect 63646 13906 63698 13918
rect 70030 13906 70082 13918
rect 8430 13858 8482 13870
rect 13918 13858 13970 13870
rect 10322 13806 10334 13858
rect 10386 13806 10398 13858
rect 10546 13806 10558 13858
rect 10610 13806 10622 13858
rect 8430 13794 8482 13806
rect 13918 13794 13970 13806
rect 14030 13858 14082 13870
rect 14030 13794 14082 13806
rect 15934 13858 15986 13870
rect 15934 13794 15986 13806
rect 23102 13858 23154 13870
rect 28366 13858 28418 13870
rect 31838 13858 31890 13870
rect 23986 13806 23998 13858
rect 24050 13806 24062 13858
rect 30482 13806 30494 13858
rect 30546 13806 30558 13858
rect 23102 13794 23154 13806
rect 28366 13794 28418 13806
rect 31838 13794 31890 13806
rect 33070 13858 33122 13870
rect 33070 13794 33122 13806
rect 33966 13858 34018 13870
rect 33966 13794 34018 13806
rect 34414 13858 34466 13870
rect 34414 13794 34466 13806
rect 35646 13858 35698 13870
rect 35646 13794 35698 13806
rect 37886 13858 37938 13870
rect 37886 13794 37938 13806
rect 40910 13858 40962 13870
rect 41694 13858 41746 13870
rect 41234 13806 41246 13858
rect 41298 13806 41310 13858
rect 40910 13794 40962 13806
rect 41694 13794 41746 13806
rect 43262 13858 43314 13870
rect 43262 13794 43314 13806
rect 43598 13858 43650 13870
rect 43598 13794 43650 13806
rect 45166 13858 45218 13870
rect 54462 13858 54514 13870
rect 61966 13858 62018 13870
rect 46722 13806 46734 13858
rect 46786 13806 46798 13858
rect 50418 13806 50430 13858
rect 50482 13806 50494 13858
rect 60722 13806 60734 13858
rect 60786 13806 60798 13858
rect 45166 13794 45218 13806
rect 54462 13794 54514 13806
rect 61966 13794 62018 13806
rect 62862 13858 62914 13870
rect 62862 13794 62914 13806
rect 63870 13858 63922 13870
rect 63870 13794 63922 13806
rect 65438 13858 65490 13870
rect 74062 13858 74114 13870
rect 66210 13806 66222 13858
rect 66274 13806 66286 13858
rect 70578 13806 70590 13858
rect 70642 13806 70654 13858
rect 71138 13806 71150 13858
rect 71202 13806 71214 13858
rect 73266 13806 73278 13858
rect 73330 13806 73342 13858
rect 65438 13794 65490 13806
rect 74062 13794 74114 13806
rect 74398 13858 74450 13870
rect 76850 13806 76862 13858
rect 76914 13806 76926 13858
rect 74398 13794 74450 13806
rect 8766 13746 8818 13758
rect 2146 13694 2158 13746
rect 2210 13694 2222 13746
rect 8766 13682 8818 13694
rect 9662 13746 9714 13758
rect 9662 13682 9714 13694
rect 9998 13746 10050 13758
rect 12350 13746 12402 13758
rect 11666 13694 11678 13746
rect 11730 13694 11742 13746
rect 12114 13694 12126 13746
rect 12178 13694 12190 13746
rect 9998 13682 10050 13694
rect 12350 13682 12402 13694
rect 12686 13746 12738 13758
rect 12686 13682 12738 13694
rect 15822 13746 15874 13758
rect 15822 13682 15874 13694
rect 16046 13746 16098 13758
rect 17614 13746 17666 13758
rect 17378 13694 17390 13746
rect 17442 13694 17454 13746
rect 16046 13682 16098 13694
rect 17614 13682 17666 13694
rect 17726 13746 17778 13758
rect 17726 13682 17778 13694
rect 17950 13746 18002 13758
rect 22990 13746 23042 13758
rect 22754 13694 22766 13746
rect 22818 13694 22830 13746
rect 17950 13682 18002 13694
rect 22990 13682 23042 13694
rect 27134 13746 27186 13758
rect 27134 13682 27186 13694
rect 28254 13746 28306 13758
rect 28254 13682 28306 13694
rect 28478 13746 28530 13758
rect 28478 13682 28530 13694
rect 29038 13746 29090 13758
rect 29038 13682 29090 13694
rect 31502 13746 31554 13758
rect 33294 13746 33346 13758
rect 32050 13694 32062 13746
rect 32114 13694 32126 13746
rect 31502 13682 31554 13694
rect 33294 13682 33346 13694
rect 33630 13746 33682 13758
rect 33630 13682 33682 13694
rect 38110 13746 38162 13758
rect 42814 13746 42866 13758
rect 42578 13694 42590 13746
rect 42642 13694 42654 13746
rect 38110 13682 38162 13694
rect 42814 13682 42866 13694
rect 42926 13746 42978 13758
rect 51662 13746 51714 13758
rect 43810 13694 43822 13746
rect 43874 13694 43886 13746
rect 44034 13694 44046 13746
rect 44098 13694 44110 13746
rect 45378 13694 45390 13746
rect 45442 13694 45454 13746
rect 47282 13694 47294 13746
rect 47346 13694 47358 13746
rect 47618 13694 47630 13746
rect 47682 13694 47694 13746
rect 49074 13694 49086 13746
rect 49138 13694 49150 13746
rect 50194 13694 50206 13746
rect 50258 13694 50270 13746
rect 42926 13682 42978 13694
rect 51662 13682 51714 13694
rect 53342 13746 53394 13758
rect 53342 13682 53394 13694
rect 54910 13746 54962 13758
rect 54910 13682 54962 13694
rect 55246 13746 55298 13758
rect 63422 13746 63474 13758
rect 70366 13746 70418 13758
rect 56690 13694 56702 13746
rect 56754 13694 56766 13746
rect 58034 13694 58046 13746
rect 58098 13694 58110 13746
rect 58370 13694 58382 13746
rect 58434 13694 58446 13746
rect 58818 13694 58830 13746
rect 58882 13694 58894 13746
rect 61282 13694 61294 13746
rect 61346 13694 61358 13746
rect 62178 13694 62190 13746
rect 62242 13694 62254 13746
rect 64418 13694 64430 13746
rect 64482 13694 64494 13746
rect 66882 13694 66894 13746
rect 66946 13694 66958 13746
rect 67890 13694 67902 13746
rect 67954 13694 67966 13746
rect 68226 13694 68238 13746
rect 68290 13694 68302 13746
rect 55246 13682 55298 13694
rect 63422 13682 63474 13694
rect 70366 13682 70418 13694
rect 71710 13746 71762 13758
rect 71710 13682 71762 13694
rect 72718 13746 72770 13758
rect 73378 13694 73390 13746
rect 73442 13694 73454 13746
rect 77634 13694 77646 13746
rect 77698 13694 77710 13746
rect 72718 13682 72770 13694
rect 7198 13634 7250 13646
rect 2930 13582 2942 13634
rect 2994 13582 3006 13634
rect 5058 13582 5070 13634
rect 5122 13582 5134 13634
rect 7198 13570 7250 13582
rect 11342 13634 11394 13646
rect 11342 13570 11394 13582
rect 12910 13634 12962 13646
rect 12910 13570 12962 13582
rect 21086 13634 21138 13646
rect 21086 13570 21138 13582
rect 25342 13634 25394 13646
rect 25342 13570 25394 13582
rect 26014 13634 26066 13646
rect 26014 13570 26066 13582
rect 26686 13634 26738 13646
rect 29486 13634 29538 13646
rect 27794 13582 27806 13634
rect 27858 13582 27870 13634
rect 26686 13570 26738 13582
rect 29486 13570 29538 13582
rect 34078 13634 34130 13646
rect 34078 13570 34130 13582
rect 36094 13634 36146 13646
rect 36094 13570 36146 13582
rect 36654 13634 36706 13646
rect 36654 13570 36706 13582
rect 37102 13634 37154 13646
rect 40014 13634 40066 13646
rect 38434 13582 38446 13634
rect 38498 13582 38510 13634
rect 37102 13570 37154 13582
rect 40014 13570 40066 13582
rect 42142 13634 42194 13646
rect 42142 13570 42194 13582
rect 43934 13634 43986 13646
rect 43934 13570 43986 13582
rect 45950 13634 46002 13646
rect 49858 13582 49870 13634
rect 49922 13582 49934 13634
rect 74722 13582 74734 13634
rect 74786 13582 74798 13634
rect 45950 13570 46002 13582
rect 13918 13522 13970 13534
rect 26910 13522 26962 13534
rect 23538 13470 23550 13522
rect 23602 13470 23614 13522
rect 13918 13458 13970 13470
rect 26910 13458 26962 13470
rect 27582 13522 27634 13534
rect 40126 13522 40178 13534
rect 30706 13470 30718 13522
rect 30770 13470 30782 13522
rect 27582 13458 27634 13470
rect 40126 13458 40178 13470
rect 52446 13522 52498 13534
rect 52446 13458 52498 13470
rect 72382 13522 72434 13534
rect 72382 13458 72434 13470
rect 1344 13354 78624 13388
rect 1344 13302 10874 13354
rect 10926 13302 10978 13354
rect 11030 13302 11082 13354
rect 11134 13302 30194 13354
rect 30246 13302 30298 13354
rect 30350 13302 30402 13354
rect 30454 13302 49514 13354
rect 49566 13302 49618 13354
rect 49670 13302 49722 13354
rect 49774 13302 68834 13354
rect 68886 13302 68938 13354
rect 68990 13302 69042 13354
rect 69094 13302 78624 13354
rect 1344 13268 78624 13302
rect 18622 13186 18674 13198
rect 18622 13122 18674 13134
rect 31278 13186 31330 13198
rect 31278 13122 31330 13134
rect 31838 13186 31890 13198
rect 31838 13122 31890 13134
rect 33070 13186 33122 13198
rect 33070 13122 33122 13134
rect 45390 13186 45442 13198
rect 45390 13122 45442 13134
rect 45726 13186 45778 13198
rect 74510 13186 74562 13198
rect 55458 13134 55470 13186
rect 55522 13183 55534 13186
rect 56242 13183 56254 13186
rect 55522 13137 56254 13183
rect 55522 13134 55534 13137
rect 56242 13134 56254 13137
rect 56306 13134 56318 13186
rect 45726 13122 45778 13134
rect 74510 13122 74562 13134
rect 16942 13074 16994 13086
rect 8082 13022 8094 13074
rect 8146 13022 8158 13074
rect 10210 13022 10222 13074
rect 10274 13022 10286 13074
rect 16942 13010 16994 13022
rect 20078 13074 20130 13086
rect 25118 13074 25170 13086
rect 29262 13074 29314 13086
rect 37214 13074 37266 13086
rect 44270 13074 44322 13086
rect 20402 13022 20414 13074
rect 20466 13022 20478 13074
rect 24210 13022 24222 13074
rect 24274 13022 24286 13074
rect 27570 13022 27582 13074
rect 27634 13022 27646 13074
rect 32722 13022 32734 13074
rect 32786 13022 32798 13074
rect 39106 13022 39118 13074
rect 39170 13022 39182 13074
rect 41906 13022 41918 13074
rect 41970 13022 41982 13074
rect 42242 13022 42254 13074
rect 42306 13022 42318 13074
rect 20078 13010 20130 13022
rect 25118 13010 25170 13022
rect 29262 13010 29314 13022
rect 37214 13010 37266 13022
rect 44270 13010 44322 13022
rect 44942 13074 44994 13086
rect 44942 13010 44994 13022
rect 50206 13074 50258 13086
rect 50206 13010 50258 13022
rect 55806 13074 55858 13086
rect 55806 13010 55858 13022
rect 56254 13074 56306 13086
rect 59726 13074 59778 13086
rect 64206 13074 64258 13086
rect 57026 13022 57038 13074
rect 57090 13022 57102 13074
rect 58482 13022 58494 13074
rect 58546 13022 58558 13074
rect 61618 13022 61630 13074
rect 61682 13022 61694 13074
rect 63746 13022 63758 13074
rect 63810 13022 63822 13074
rect 65314 13022 65326 13074
rect 65378 13022 65390 13074
rect 72594 13022 72606 13074
rect 72658 13022 72670 13074
rect 56254 13010 56306 13022
rect 59726 13010 59778 13022
rect 64206 13010 64258 13022
rect 2718 12962 2770 12974
rect 2718 12898 2770 12910
rect 3614 12962 3666 12974
rect 14590 12962 14642 12974
rect 7410 12910 7422 12962
rect 7474 12910 7486 12962
rect 3614 12898 3666 12910
rect 14590 12898 14642 12910
rect 15934 12962 15986 12974
rect 15934 12898 15986 12910
rect 16270 12962 16322 12974
rect 16270 12898 16322 12910
rect 16382 12962 16434 12974
rect 19518 12962 19570 12974
rect 20862 12962 20914 12974
rect 22990 12962 23042 12974
rect 17490 12910 17502 12962
rect 17554 12910 17566 12962
rect 18274 12910 18286 12962
rect 18338 12910 18350 12962
rect 20514 12910 20526 12962
rect 20578 12910 20590 12962
rect 21522 12910 21534 12962
rect 21586 12910 21598 12962
rect 16382 12898 16434 12910
rect 19518 12898 19570 12910
rect 20862 12898 20914 12910
rect 22990 12898 23042 12910
rect 24446 12962 24498 12974
rect 24446 12898 24498 12910
rect 24894 12962 24946 12974
rect 26126 12962 26178 12974
rect 32286 12962 32338 12974
rect 35198 12962 35250 12974
rect 25218 12910 25230 12962
rect 25282 12910 25294 12962
rect 26450 12910 26462 12962
rect 26514 12910 26526 12962
rect 26674 12910 26686 12962
rect 26738 12910 26750 12962
rect 27906 12910 27918 12962
rect 27970 12910 27982 12962
rect 28690 12910 28702 12962
rect 28754 12910 28766 12962
rect 32834 12910 32846 12962
rect 32898 12910 32910 12962
rect 33282 12910 33294 12962
rect 33346 12910 33358 12962
rect 33730 12910 33742 12962
rect 33794 12910 33806 12962
rect 34626 12910 34638 12962
rect 34690 12910 34702 12962
rect 34962 12910 34974 12962
rect 35026 12910 35038 12962
rect 24894 12898 24946 12910
rect 26126 12898 26178 12910
rect 32286 12898 32338 12910
rect 35198 12898 35250 12910
rect 35310 12962 35362 12974
rect 35310 12898 35362 12910
rect 35422 12962 35474 12974
rect 55358 12962 55410 12974
rect 37650 12910 37662 12962
rect 37714 12910 37726 12962
rect 39666 12910 39678 12962
rect 39730 12910 39742 12962
rect 40338 12910 40350 12962
rect 40402 12910 40414 12962
rect 41458 12910 41470 12962
rect 41522 12910 41534 12962
rect 42354 12910 42366 12962
rect 42418 12910 42430 12962
rect 46386 12910 46398 12962
rect 46450 12910 46462 12962
rect 47058 12910 47070 12962
rect 47122 12910 47134 12962
rect 48290 12910 48302 12962
rect 48354 12910 48366 12962
rect 48626 12910 48638 12962
rect 48690 12910 48702 12962
rect 48962 12910 48974 12962
rect 49026 12910 49038 12962
rect 51538 12910 51550 12962
rect 51602 12910 51614 12962
rect 35422 12898 35474 12910
rect 55358 12898 55410 12910
rect 56702 12962 56754 12974
rect 56702 12898 56754 12910
rect 56814 12962 56866 12974
rect 56814 12898 56866 12910
rect 57150 12962 57202 12974
rect 57810 12910 57822 12962
rect 57874 12910 57886 12962
rect 59266 12910 59278 12962
rect 59330 12910 59342 12962
rect 60834 12910 60846 12962
rect 60898 12910 60910 12962
rect 65538 12910 65550 12962
rect 65602 12910 65614 12962
rect 66210 12910 66222 12962
rect 66274 12910 66286 12962
rect 66658 12910 66670 12962
rect 66722 12910 66734 12962
rect 69682 12910 69694 12962
rect 69746 12910 69758 12962
rect 73154 12910 73166 12962
rect 73218 12910 73230 12962
rect 73938 12910 73950 12962
rect 74002 12910 74014 12962
rect 57150 12898 57202 12910
rect 2382 12850 2434 12862
rect 2382 12786 2434 12798
rect 3278 12850 3330 12862
rect 3278 12786 3330 12798
rect 6526 12850 6578 12862
rect 6526 12786 6578 12798
rect 11790 12850 11842 12862
rect 11790 12786 11842 12798
rect 12798 12850 12850 12862
rect 17278 12850 17330 12862
rect 13794 12798 13806 12850
rect 13858 12798 13870 12850
rect 14018 12798 14030 12850
rect 14082 12798 14094 12850
rect 12798 12786 12850 12798
rect 17278 12786 17330 12798
rect 17726 12850 17778 12862
rect 17726 12786 17778 12798
rect 17838 12850 17890 12862
rect 17838 12786 17890 12798
rect 18062 12850 18114 12862
rect 18062 12786 18114 12798
rect 18846 12850 18898 12862
rect 18846 12786 18898 12798
rect 18958 12850 19010 12862
rect 18958 12786 19010 12798
rect 20302 12850 20354 12862
rect 20302 12786 20354 12798
rect 21758 12850 21810 12862
rect 21758 12786 21810 12798
rect 24222 12850 24274 12862
rect 24222 12786 24274 12798
rect 24670 12850 24722 12862
rect 31390 12850 31442 12862
rect 27234 12798 27246 12850
rect 27298 12798 27310 12850
rect 24670 12786 24722 12798
rect 31390 12786 31442 12798
rect 31726 12850 31778 12862
rect 50878 12850 50930 12862
rect 34514 12798 34526 12850
rect 34578 12798 34590 12850
rect 46274 12798 46286 12850
rect 46338 12798 46350 12850
rect 31726 12786 31778 12798
rect 50878 12786 50930 12798
rect 57038 12850 57090 12862
rect 57922 12798 57934 12850
rect 57986 12798 57998 12850
rect 64866 12798 64878 12850
rect 64930 12798 64942 12850
rect 66882 12798 66894 12850
rect 66946 12798 66958 12850
rect 70354 12798 70366 12850
rect 70418 12798 70430 12850
rect 72930 12798 72942 12850
rect 72994 12847 73006 12850
rect 73169 12847 73215 12910
rect 74846 12850 74898 12862
rect 72994 12801 73215 12847
rect 72994 12798 73006 12801
rect 73714 12798 73726 12850
rect 73778 12798 73790 12850
rect 57038 12786 57090 12798
rect 74846 12786 74898 12798
rect 75294 12850 75346 12862
rect 75294 12786 75346 12798
rect 6190 12738 6242 12750
rect 6190 12674 6242 12686
rect 11902 12738 11954 12750
rect 11902 12674 11954 12686
rect 12910 12738 12962 12750
rect 15038 12738 15090 12750
rect 14242 12686 14254 12738
rect 14306 12686 14318 12738
rect 12910 12674 12962 12686
rect 15038 12674 15090 12686
rect 15486 12738 15538 12750
rect 15486 12674 15538 12686
rect 16046 12738 16098 12750
rect 16046 12674 16098 12686
rect 16158 12738 16210 12750
rect 16158 12674 16210 12686
rect 18510 12738 18562 12750
rect 18510 12674 18562 12686
rect 19182 12738 19234 12750
rect 19182 12674 19234 12686
rect 21198 12738 21250 12750
rect 21198 12674 21250 12686
rect 21310 12738 21362 12750
rect 21310 12674 21362 12686
rect 23774 12738 23826 12750
rect 23774 12674 23826 12686
rect 24110 12738 24162 12750
rect 24110 12674 24162 12686
rect 25454 12738 25506 12750
rect 25454 12674 25506 12686
rect 26910 12738 26962 12750
rect 26910 12674 26962 12686
rect 27022 12738 27074 12750
rect 27022 12674 27074 12686
rect 32398 12738 32450 12750
rect 32398 12674 32450 12686
rect 32622 12738 32674 12750
rect 32622 12674 32674 12686
rect 35534 12738 35586 12750
rect 35534 12674 35586 12686
rect 36094 12738 36146 12750
rect 59054 12738 59106 12750
rect 36418 12686 36430 12738
rect 36482 12686 36494 12738
rect 37426 12686 37438 12738
rect 37490 12686 37502 12738
rect 36094 12674 36146 12686
rect 59054 12674 59106 12686
rect 64654 12738 64706 12750
rect 64654 12674 64706 12686
rect 73278 12738 73330 12750
rect 73278 12674 73330 12686
rect 75630 12738 75682 12750
rect 75630 12674 75682 12686
rect 1344 12570 78784 12604
rect 1344 12518 20534 12570
rect 20586 12518 20638 12570
rect 20690 12518 20742 12570
rect 20794 12518 39854 12570
rect 39906 12518 39958 12570
rect 40010 12518 40062 12570
rect 40114 12518 59174 12570
rect 59226 12518 59278 12570
rect 59330 12518 59382 12570
rect 59434 12518 78494 12570
rect 78546 12518 78598 12570
rect 78650 12518 78702 12570
rect 78754 12518 78784 12570
rect 1344 12484 78784 12518
rect 23214 12402 23266 12414
rect 32062 12402 32114 12414
rect 25218 12350 25230 12402
rect 25282 12350 25294 12402
rect 23214 12338 23266 12350
rect 32062 12338 32114 12350
rect 33518 12402 33570 12414
rect 33518 12338 33570 12350
rect 33630 12402 33682 12414
rect 33630 12338 33682 12350
rect 33854 12402 33906 12414
rect 33854 12338 33906 12350
rect 34526 12402 34578 12414
rect 34526 12338 34578 12350
rect 38670 12402 38722 12414
rect 38670 12338 38722 12350
rect 39454 12402 39506 12414
rect 39454 12338 39506 12350
rect 41470 12402 41522 12414
rect 41470 12338 41522 12350
rect 41694 12402 41746 12414
rect 41694 12338 41746 12350
rect 42366 12402 42418 12414
rect 42366 12338 42418 12350
rect 43598 12402 43650 12414
rect 43598 12338 43650 12350
rect 47854 12402 47906 12414
rect 55806 12402 55858 12414
rect 53554 12350 53566 12402
rect 53618 12350 53630 12402
rect 47854 12338 47906 12350
rect 55806 12338 55858 12350
rect 56814 12402 56866 12414
rect 56814 12338 56866 12350
rect 57374 12402 57426 12414
rect 57374 12338 57426 12350
rect 58158 12402 58210 12414
rect 58158 12338 58210 12350
rect 58382 12402 58434 12414
rect 61070 12402 61122 12414
rect 60162 12350 60174 12402
rect 60226 12350 60238 12402
rect 60386 12350 60398 12402
rect 60450 12350 60462 12402
rect 58382 12338 58434 12350
rect 61070 12338 61122 12350
rect 61742 12402 61794 12414
rect 61742 12338 61794 12350
rect 64542 12402 64594 12414
rect 64542 12338 64594 12350
rect 65102 12402 65154 12414
rect 69806 12402 69858 12414
rect 65650 12350 65662 12402
rect 65714 12350 65726 12402
rect 65874 12350 65886 12402
rect 65938 12350 65950 12402
rect 65102 12338 65154 12350
rect 69806 12338 69858 12350
rect 70478 12402 70530 12414
rect 70478 12338 70530 12350
rect 2830 12290 2882 12302
rect 18958 12290 19010 12302
rect 6290 12238 6302 12290
rect 6354 12238 6366 12290
rect 17602 12238 17614 12290
rect 17666 12238 17678 12290
rect 2830 12226 2882 12238
rect 18958 12226 19010 12238
rect 20638 12290 20690 12302
rect 20638 12226 20690 12238
rect 20974 12290 21026 12302
rect 20974 12226 21026 12238
rect 22430 12290 22482 12302
rect 22430 12226 22482 12238
rect 23998 12290 24050 12302
rect 28702 12290 28754 12302
rect 26786 12238 26798 12290
rect 26850 12238 26862 12290
rect 28130 12238 28142 12290
rect 28194 12238 28206 12290
rect 23998 12226 24050 12238
rect 28702 12226 28754 12238
rect 33294 12290 33346 12302
rect 41246 12290 41298 12302
rect 38994 12238 39006 12290
rect 39058 12238 39070 12290
rect 40114 12238 40126 12290
rect 40178 12238 40190 12290
rect 33294 12226 33346 12238
rect 41246 12226 41298 12238
rect 41806 12290 41858 12302
rect 54238 12290 54290 12302
rect 70814 12290 70866 12302
rect 45154 12238 45166 12290
rect 45218 12238 45230 12290
rect 53442 12238 53454 12290
rect 53506 12238 53518 12290
rect 59378 12238 59390 12290
rect 59442 12238 59454 12290
rect 62402 12238 62414 12290
rect 62466 12238 62478 12290
rect 62850 12238 62862 12290
rect 62914 12238 62926 12290
rect 66546 12238 66558 12290
rect 66610 12238 66622 12290
rect 77074 12238 77086 12290
rect 77138 12238 77150 12290
rect 41806 12226 41858 12238
rect 54238 12226 54290 12238
rect 70814 12226 70866 12238
rect 3166 12178 3218 12190
rect 18622 12178 18674 12190
rect 5506 12126 5518 12178
rect 5570 12126 5582 12178
rect 12338 12126 12350 12178
rect 12402 12126 12414 12178
rect 12674 12126 12686 12178
rect 12738 12126 12750 12178
rect 14242 12126 14254 12178
rect 14306 12126 14318 12178
rect 15698 12126 15710 12178
rect 15762 12126 15774 12178
rect 3166 12114 3218 12126
rect 18622 12114 18674 12126
rect 18846 12178 18898 12190
rect 18846 12114 18898 12126
rect 19406 12178 19458 12190
rect 19406 12114 19458 12126
rect 19854 12178 19906 12190
rect 19854 12114 19906 12126
rect 20414 12178 20466 12190
rect 20414 12114 20466 12126
rect 22878 12178 22930 12190
rect 22878 12114 22930 12126
rect 24222 12178 24274 12190
rect 24222 12114 24274 12126
rect 24334 12178 24386 12190
rect 24334 12114 24386 12126
rect 24446 12178 24498 12190
rect 25678 12178 25730 12190
rect 24658 12126 24670 12178
rect 24722 12126 24734 12178
rect 24446 12114 24498 12126
rect 25678 12114 25730 12126
rect 25790 12178 25842 12190
rect 28926 12178 28978 12190
rect 26002 12126 26014 12178
rect 26066 12126 26078 12178
rect 27010 12126 27022 12178
rect 27074 12126 27086 12178
rect 27906 12126 27918 12178
rect 27970 12126 27982 12178
rect 25790 12114 25842 12126
rect 28926 12114 28978 12126
rect 33742 12178 33794 12190
rect 42478 12178 42530 12190
rect 36194 12126 36206 12178
rect 36258 12126 36270 12178
rect 38098 12126 38110 12178
rect 38162 12126 38174 12178
rect 39890 12126 39902 12178
rect 39954 12126 39966 12178
rect 33742 12114 33794 12126
rect 42478 12114 42530 12126
rect 42814 12178 42866 12190
rect 43486 12178 43538 12190
rect 57934 12178 57986 12190
rect 43026 12126 43038 12178
rect 43090 12126 43102 12178
rect 44482 12126 44494 12178
rect 44546 12126 44558 12178
rect 50642 12126 50654 12178
rect 50706 12126 50718 12178
rect 51762 12126 51774 12178
rect 51826 12126 51838 12178
rect 52322 12126 52334 12178
rect 52386 12126 52398 12178
rect 54898 12126 54910 12178
rect 54962 12126 54974 12178
rect 42814 12114 42866 12126
rect 43486 12114 43538 12126
rect 57934 12114 57986 12126
rect 58046 12178 58098 12190
rect 58046 12114 58098 12126
rect 58270 12178 58322 12190
rect 62078 12178 62130 12190
rect 59042 12126 59054 12178
rect 59106 12126 59118 12178
rect 60386 12126 60398 12178
rect 60450 12126 60462 12178
rect 58270 12114 58322 12126
rect 62078 12114 62130 12126
rect 63422 12178 63474 12190
rect 63422 12114 63474 12126
rect 63870 12178 63922 12190
rect 70142 12178 70194 12190
rect 65538 12126 65550 12178
rect 65602 12126 65614 12178
rect 66882 12126 66894 12178
rect 66946 12126 66958 12178
rect 77746 12126 77758 12178
rect 77810 12126 77822 12178
rect 63870 12114 63922 12126
rect 70142 12114 70194 12126
rect 12126 12066 12178 12078
rect 22206 12066 22258 12078
rect 8418 12014 8430 12066
rect 8482 12014 8494 12066
rect 15810 12014 15822 12066
rect 15874 12014 15886 12066
rect 21298 12014 21310 12066
rect 21362 12014 21374 12066
rect 12126 12002 12178 12014
rect 22206 12002 22258 12014
rect 23662 12066 23714 12078
rect 32510 12066 32562 12078
rect 39342 12066 39394 12078
rect 43150 12066 43202 12078
rect 27682 12014 27694 12066
rect 27746 12014 27758 12066
rect 35410 12014 35422 12066
rect 35474 12014 35486 12066
rect 36978 12014 36990 12066
rect 37042 12014 37054 12066
rect 41794 12014 41806 12066
rect 41858 12014 41870 12066
rect 23662 12002 23714 12014
rect 32510 12002 32562 12014
rect 39342 12002 39394 12014
rect 43150 12002 43202 12014
rect 43934 12066 43986 12078
rect 50094 12066 50146 12078
rect 47282 12014 47294 12066
rect 47346 12014 47358 12066
rect 74946 12014 74958 12066
rect 75010 12014 75022 12066
rect 43934 12002 43986 12014
rect 50094 12002 50146 12014
rect 20078 11954 20130 11966
rect 16258 11902 16270 11954
rect 16322 11902 16334 11954
rect 20078 11890 20130 11902
rect 20526 11954 20578 11966
rect 20526 11890 20578 11902
rect 29262 11954 29314 11966
rect 31938 11902 31950 11954
rect 32002 11951 32014 11954
rect 32610 11951 32622 11954
rect 32002 11905 32622 11951
rect 32002 11902 32014 11905
rect 32610 11902 32622 11905
rect 32674 11902 32686 11954
rect 29262 11890 29314 11902
rect 1344 11786 78624 11820
rect 1344 11734 10874 11786
rect 10926 11734 10978 11786
rect 11030 11734 11082 11786
rect 11134 11734 30194 11786
rect 30246 11734 30298 11786
rect 30350 11734 30402 11786
rect 30454 11734 49514 11786
rect 49566 11734 49618 11786
rect 49670 11734 49722 11786
rect 49774 11734 68834 11786
rect 68886 11734 68938 11786
rect 68990 11734 69042 11786
rect 69094 11734 78624 11786
rect 1344 11700 78624 11734
rect 6638 11618 6690 11630
rect 19182 11618 19234 11630
rect 18386 11566 18398 11618
rect 18450 11566 18462 11618
rect 6638 11554 6690 11566
rect 19182 11554 19234 11566
rect 19294 11618 19346 11630
rect 19294 11554 19346 11566
rect 19518 11618 19570 11630
rect 19518 11554 19570 11566
rect 21758 11618 21810 11630
rect 21758 11554 21810 11566
rect 48190 11618 48242 11630
rect 48190 11554 48242 11566
rect 5070 11506 5122 11518
rect 2482 11454 2494 11506
rect 2546 11454 2558 11506
rect 4610 11454 4622 11506
rect 4674 11454 4686 11506
rect 5070 11442 5122 11454
rect 6974 11506 7026 11518
rect 6974 11442 7026 11454
rect 8318 11506 8370 11518
rect 8318 11442 8370 11454
rect 16494 11506 16546 11518
rect 16494 11442 16546 11454
rect 17278 11506 17330 11518
rect 21310 11506 21362 11518
rect 18274 11454 18286 11506
rect 18338 11454 18350 11506
rect 17278 11442 17330 11454
rect 21310 11442 21362 11454
rect 22206 11506 22258 11518
rect 22206 11442 22258 11454
rect 26798 11506 26850 11518
rect 26798 11442 26850 11454
rect 27246 11506 27298 11518
rect 27246 11442 27298 11454
rect 27470 11506 27522 11518
rect 27470 11442 27522 11454
rect 31950 11506 32002 11518
rect 31950 11442 32002 11454
rect 34190 11506 34242 11518
rect 34190 11442 34242 11454
rect 35982 11506 36034 11518
rect 35982 11442 36034 11454
rect 39006 11506 39058 11518
rect 39006 11442 39058 11454
rect 40014 11506 40066 11518
rect 40014 11442 40066 11454
rect 40350 11506 40402 11518
rect 40350 11442 40402 11454
rect 40798 11506 40850 11518
rect 40798 11442 40850 11454
rect 42142 11506 42194 11518
rect 42142 11442 42194 11454
rect 42366 11506 42418 11518
rect 46734 11506 46786 11518
rect 43586 11454 43598 11506
rect 43650 11454 43662 11506
rect 42366 11442 42418 11454
rect 46734 11442 46786 11454
rect 50206 11506 50258 11518
rect 50206 11442 50258 11454
rect 56030 11506 56082 11518
rect 56030 11442 56082 11454
rect 57374 11506 57426 11518
rect 57374 11442 57426 11454
rect 60734 11506 60786 11518
rect 60734 11442 60786 11454
rect 61518 11506 61570 11518
rect 67778 11454 67790 11506
rect 67842 11454 67854 11506
rect 61518 11442 61570 11454
rect 14590 11394 14642 11406
rect 1810 11342 1822 11394
rect 1874 11342 1886 11394
rect 7746 11342 7758 11394
rect 7810 11342 7822 11394
rect 14590 11330 14642 11342
rect 15262 11394 15314 11406
rect 15262 11330 15314 11342
rect 15934 11394 15986 11406
rect 15934 11330 15986 11342
rect 16718 11394 16770 11406
rect 16718 11330 16770 11342
rect 16830 11394 16882 11406
rect 16830 11330 16882 11342
rect 21534 11394 21586 11406
rect 21534 11330 21586 11342
rect 22766 11394 22818 11406
rect 23550 11394 23602 11406
rect 23202 11342 23214 11394
rect 23266 11342 23278 11394
rect 22766 11330 22818 11342
rect 23550 11330 23602 11342
rect 23774 11394 23826 11406
rect 23774 11330 23826 11342
rect 24446 11394 24498 11406
rect 24446 11330 24498 11342
rect 25342 11394 25394 11406
rect 25342 11330 25394 11342
rect 25566 11394 25618 11406
rect 25566 11330 25618 11342
rect 25678 11394 25730 11406
rect 25678 11330 25730 11342
rect 27134 11394 27186 11406
rect 27134 11330 27186 11342
rect 27694 11394 27746 11406
rect 27694 11330 27746 11342
rect 28030 11394 28082 11406
rect 28030 11330 28082 11342
rect 28142 11394 28194 11406
rect 29262 11394 29314 11406
rect 28354 11342 28366 11394
rect 28418 11342 28430 11394
rect 28142 11330 28194 11342
rect 29262 11330 29314 11342
rect 30718 11394 30770 11406
rect 30718 11330 30770 11342
rect 31166 11394 31218 11406
rect 31166 11330 31218 11342
rect 31838 11394 31890 11406
rect 41694 11394 41746 11406
rect 43822 11394 43874 11406
rect 44942 11394 44994 11406
rect 38210 11342 38222 11394
rect 38274 11342 38286 11394
rect 43362 11342 43374 11394
rect 43426 11342 43438 11394
rect 44034 11342 44046 11394
rect 44098 11342 44110 11394
rect 31838 11330 31890 11342
rect 41694 11330 41746 11342
rect 43822 11330 43874 11342
rect 44942 11330 44994 11342
rect 49758 11394 49810 11406
rect 49758 11330 49810 11342
rect 53118 11394 53170 11406
rect 58382 11394 58434 11406
rect 53890 11342 53902 11394
rect 53954 11342 53966 11394
rect 55010 11342 55022 11394
rect 55074 11342 55086 11394
rect 57698 11342 57710 11394
rect 57762 11342 57774 11394
rect 53118 11330 53170 11342
rect 58382 11330 58434 11342
rect 58718 11394 58770 11406
rect 59378 11342 59390 11394
rect 59442 11342 59454 11394
rect 64978 11342 64990 11394
rect 65042 11342 65054 11394
rect 75618 11342 75630 11394
rect 75682 11342 75694 11394
rect 58718 11330 58770 11342
rect 12014 11282 12066 11294
rect 7522 11230 7534 11282
rect 7586 11230 7598 11282
rect 12014 11218 12066 11230
rect 12798 11282 12850 11294
rect 15486 11282 15538 11294
rect 13794 11230 13806 11282
rect 13858 11230 13870 11282
rect 14018 11230 14030 11282
rect 14082 11230 14094 11282
rect 12798 11218 12850 11230
rect 15486 11218 15538 11230
rect 16158 11282 16210 11294
rect 22542 11282 22594 11294
rect 18610 11230 18622 11282
rect 18674 11230 18686 11282
rect 16158 11218 16210 11230
rect 22542 11218 22594 11230
rect 24110 11282 24162 11294
rect 24110 11218 24162 11230
rect 24558 11282 24610 11294
rect 24558 11218 24610 11230
rect 25118 11282 25170 11294
rect 41806 11282 41858 11294
rect 52110 11282 52162 11294
rect 37986 11230 37998 11282
rect 38050 11230 38062 11282
rect 48514 11230 48526 11282
rect 48578 11230 48590 11282
rect 48850 11230 48862 11282
rect 48914 11230 48926 11282
rect 25118 11218 25170 11230
rect 41806 11218 41858 11230
rect 52110 11218 52162 11230
rect 52782 11282 52834 11294
rect 72494 11282 72546 11294
rect 53778 11230 53790 11282
rect 53842 11230 53854 11282
rect 59490 11230 59502 11282
rect 59554 11230 59566 11282
rect 65650 11230 65662 11282
rect 65714 11230 65726 11282
rect 52782 11218 52834 11230
rect 72494 11218 72546 11230
rect 72606 11282 72658 11294
rect 72606 11218 72658 11230
rect 76750 11282 76802 11294
rect 76750 11218 76802 11230
rect 77086 11282 77138 11294
rect 77086 11218 77138 11230
rect 8766 11170 8818 11182
rect 8766 11106 8818 11118
rect 11230 11170 11282 11182
rect 11230 11106 11282 11118
rect 11790 11170 11842 11182
rect 11790 11106 11842 11118
rect 12126 11170 12178 11182
rect 12126 11106 12178 11118
rect 12910 11170 12962 11182
rect 15374 11170 15426 11182
rect 14242 11118 14254 11170
rect 14306 11118 14318 11170
rect 12910 11106 12962 11118
rect 15374 11106 15426 11118
rect 16382 11170 16434 11182
rect 16382 11106 16434 11118
rect 19966 11170 20018 11182
rect 19966 11106 20018 11118
rect 22878 11170 22930 11182
rect 22878 11106 22930 11118
rect 22990 11170 23042 11182
rect 22990 11106 23042 11118
rect 23998 11170 24050 11182
rect 23998 11106 24050 11118
rect 24670 11170 24722 11182
rect 24670 11106 24722 11118
rect 25454 11170 25506 11182
rect 25454 11106 25506 11118
rect 26350 11170 26402 11182
rect 26350 11106 26402 11118
rect 29710 11170 29762 11182
rect 29710 11106 29762 11118
rect 30158 11170 30210 11182
rect 30158 11106 30210 11118
rect 30494 11170 30546 11182
rect 30494 11106 30546 11118
rect 30606 11170 30658 11182
rect 30606 11106 30658 11118
rect 33182 11170 33234 11182
rect 33182 11106 33234 11118
rect 36430 11170 36482 11182
rect 37326 11170 37378 11182
rect 36978 11118 36990 11170
rect 37042 11118 37054 11170
rect 36430 11106 36482 11118
rect 37326 11106 37378 11118
rect 39454 11170 39506 11182
rect 39454 11106 39506 11118
rect 41246 11170 41298 11182
rect 41246 11106 41298 11118
rect 41358 11170 41410 11182
rect 41358 11106 41410 11118
rect 41918 11170 41970 11182
rect 41918 11106 41970 11118
rect 42814 11170 42866 11182
rect 42814 11106 42866 11118
rect 43598 11170 43650 11182
rect 43598 11106 43650 11118
rect 47854 11170 47906 11182
rect 51774 11170 51826 11182
rect 49410 11118 49422 11170
rect 49474 11118 49486 11170
rect 47854 11106 47906 11118
rect 51774 11106 51826 11118
rect 54462 11170 54514 11182
rect 54462 11106 54514 11118
rect 54798 11170 54850 11182
rect 54798 11106 54850 11118
rect 56814 11170 56866 11182
rect 56814 11106 56866 11118
rect 57934 11170 57986 11182
rect 57934 11106 57986 11118
rect 61070 11170 61122 11182
rect 61070 11106 61122 11118
rect 72270 11170 72322 11182
rect 72270 11106 72322 11118
rect 72830 11170 72882 11182
rect 72830 11106 72882 11118
rect 74622 11170 74674 11182
rect 74622 11106 74674 11118
rect 76414 11170 76466 11182
rect 76414 11106 76466 11118
rect 1344 11002 78784 11036
rect 1344 10950 20534 11002
rect 20586 10950 20638 11002
rect 20690 10950 20742 11002
rect 20794 10950 39854 11002
rect 39906 10950 39958 11002
rect 40010 10950 40062 11002
rect 40114 10950 59174 11002
rect 59226 10950 59278 11002
rect 59330 10950 59382 11002
rect 59434 10950 78494 11002
rect 78546 10950 78598 11002
rect 78650 10950 78702 11002
rect 78754 10950 78784 11002
rect 1344 10916 78784 10950
rect 4734 10834 4786 10846
rect 4734 10770 4786 10782
rect 17278 10834 17330 10846
rect 17278 10770 17330 10782
rect 18062 10834 18114 10846
rect 18062 10770 18114 10782
rect 20190 10834 20242 10846
rect 20190 10770 20242 10782
rect 20974 10834 21026 10846
rect 20974 10770 21026 10782
rect 21198 10834 21250 10846
rect 21198 10770 21250 10782
rect 23214 10834 23266 10846
rect 25454 10834 25506 10846
rect 24658 10782 24670 10834
rect 24722 10782 24734 10834
rect 23214 10770 23266 10782
rect 25454 10770 25506 10782
rect 26126 10834 26178 10846
rect 26126 10770 26178 10782
rect 27806 10834 27858 10846
rect 27806 10770 27858 10782
rect 37886 10834 37938 10846
rect 37886 10770 37938 10782
rect 38222 10834 38274 10846
rect 38222 10770 38274 10782
rect 41694 10834 41746 10846
rect 41694 10770 41746 10782
rect 42702 10834 42754 10846
rect 42702 10770 42754 10782
rect 46398 10834 46450 10846
rect 46398 10770 46450 10782
rect 54350 10834 54402 10846
rect 54350 10770 54402 10782
rect 54798 10834 54850 10846
rect 54798 10770 54850 10782
rect 56702 10834 56754 10846
rect 56702 10770 56754 10782
rect 66446 10834 66498 10846
rect 66446 10770 66498 10782
rect 67230 10834 67282 10846
rect 67230 10770 67282 10782
rect 68126 10834 68178 10846
rect 68126 10770 68178 10782
rect 76526 10834 76578 10846
rect 76526 10770 76578 10782
rect 8878 10722 8930 10734
rect 5842 10670 5854 10722
rect 5906 10670 5918 10722
rect 8878 10658 8930 10670
rect 9550 10722 9602 10734
rect 9550 10658 9602 10670
rect 17502 10722 17554 10734
rect 17502 10658 17554 10670
rect 19966 10722 20018 10734
rect 19966 10658 20018 10670
rect 20414 10722 20466 10734
rect 20414 10658 20466 10670
rect 22654 10722 22706 10734
rect 33966 10722 34018 10734
rect 41918 10722 41970 10734
rect 22654 10658 22706 10670
rect 24222 10666 24274 10678
rect 30370 10670 30382 10722
rect 30434 10670 30446 10722
rect 39666 10670 39678 10722
rect 39730 10670 39742 10722
rect 40002 10670 40014 10722
rect 40066 10670 40078 10722
rect 10110 10610 10162 10622
rect 17614 10610 17666 10622
rect 4274 10558 4286 10610
rect 4338 10558 4350 10610
rect 5618 10558 5630 10610
rect 5682 10558 5694 10610
rect 8642 10558 8654 10610
rect 8706 10558 8718 10610
rect 12338 10558 12350 10610
rect 12402 10558 12414 10610
rect 12562 10558 12574 10610
rect 12626 10558 12638 10610
rect 14242 10558 14254 10610
rect 14306 10558 14318 10610
rect 15474 10558 15486 10610
rect 15538 10558 15550 10610
rect 10110 10546 10162 10558
rect 17614 10546 17666 10558
rect 20526 10610 20578 10622
rect 20526 10546 20578 10558
rect 20862 10610 20914 10622
rect 20862 10546 20914 10558
rect 22206 10610 22258 10622
rect 24110 10610 24162 10622
rect 23874 10558 23886 10610
rect 23938 10558 23950 10610
rect 33966 10658 34018 10670
rect 41918 10658 41970 10670
rect 47854 10722 47906 10734
rect 47854 10658 47906 10670
rect 48190 10722 48242 10734
rect 61742 10722 61794 10734
rect 69358 10722 69410 10734
rect 51650 10670 51662 10722
rect 51714 10670 51726 10722
rect 55906 10670 55918 10722
rect 55970 10670 55982 10722
rect 64978 10670 64990 10722
rect 65042 10670 65054 10722
rect 65426 10670 65438 10722
rect 65490 10670 65502 10722
rect 48190 10658 48242 10670
rect 61742 10658 61794 10670
rect 69358 10658 69410 10670
rect 69582 10722 69634 10734
rect 76738 10670 76750 10722
rect 76802 10670 76814 10722
rect 77410 10670 77422 10722
rect 77474 10670 77486 10722
rect 69582 10658 69634 10670
rect 24222 10602 24274 10614
rect 28590 10610 28642 10622
rect 34302 10610 34354 10622
rect 22206 10546 22258 10558
rect 24110 10546 24162 10558
rect 29698 10558 29710 10610
rect 29762 10558 29774 10610
rect 28590 10546 28642 10558
rect 34302 10546 34354 10558
rect 42254 10610 42306 10622
rect 43374 10610 43426 10622
rect 43138 10558 43150 10610
rect 43202 10558 43214 10610
rect 42254 10546 42306 10558
rect 43374 10546 43426 10558
rect 43598 10610 43650 10622
rect 65998 10610 66050 10622
rect 43810 10558 43822 10610
rect 43874 10558 43886 10610
rect 50866 10558 50878 10610
rect 50930 10558 50942 10610
rect 55794 10558 55806 10610
rect 55858 10558 55870 10610
rect 57922 10558 57934 10610
rect 57986 10558 57998 10610
rect 61954 10558 61966 10610
rect 62018 10558 62030 10610
rect 43598 10546 43650 10558
rect 65998 10546 66050 10558
rect 66782 10610 66834 10622
rect 66782 10546 66834 10558
rect 69134 10610 69186 10622
rect 72594 10558 72606 10610
rect 72658 10558 72670 10610
rect 76962 10558 76974 10610
rect 77026 10558 77038 10610
rect 77634 10558 77646 10610
rect 77698 10558 77710 10610
rect 69134 10546 69186 10558
rect 1934 10498 1986 10510
rect 1934 10434 1986 10446
rect 6414 10498 6466 10510
rect 6414 10434 6466 10446
rect 6974 10498 7026 10510
rect 6974 10434 7026 10446
rect 10558 10498 10610 10510
rect 18510 10498 18562 10510
rect 15698 10446 15710 10498
rect 15762 10446 15774 10498
rect 10558 10434 10610 10446
rect 18510 10434 18562 10446
rect 21758 10498 21810 10510
rect 21758 10434 21810 10446
rect 23662 10498 23714 10510
rect 23662 10434 23714 10446
rect 27694 10498 27746 10510
rect 38670 10498 38722 10510
rect 32498 10446 32510 10498
rect 32562 10446 32574 10498
rect 27694 10434 27746 10446
rect 38670 10434 38722 10446
rect 41134 10498 41186 10510
rect 41134 10434 41186 10446
rect 43486 10498 43538 10510
rect 43486 10434 43538 10446
rect 44270 10498 44322 10510
rect 63870 10498 63922 10510
rect 53778 10446 53790 10498
rect 53842 10446 53854 10498
rect 58594 10446 58606 10498
rect 58658 10446 58670 10498
rect 60722 10446 60734 10498
rect 60786 10446 60798 10498
rect 44270 10434 44322 10446
rect 63870 10434 63922 10446
rect 65662 10498 65714 10510
rect 65662 10434 65714 10446
rect 68574 10498 68626 10510
rect 68574 10434 68626 10446
rect 69246 10498 69298 10510
rect 76078 10498 76130 10510
rect 73378 10446 73390 10498
rect 73442 10446 73454 10498
rect 75506 10446 75518 10498
rect 75570 10446 75582 10498
rect 69246 10434 69298 10446
rect 76078 10434 76130 10446
rect 5070 10386 5122 10398
rect 39118 10386 39170 10398
rect 16034 10334 16046 10386
rect 16098 10334 16110 10386
rect 5070 10322 5122 10334
rect 39118 10322 39170 10334
rect 39454 10386 39506 10398
rect 41582 10386 41634 10398
rect 41122 10334 41134 10386
rect 41186 10383 41198 10386
rect 41458 10383 41470 10386
rect 41186 10337 41470 10383
rect 41186 10334 41198 10337
rect 41458 10334 41470 10337
rect 41522 10334 41534 10386
rect 39454 10322 39506 10334
rect 41582 10322 41634 10334
rect 55134 10386 55186 10398
rect 75730 10334 75742 10386
rect 75794 10383 75806 10386
rect 76514 10383 76526 10386
rect 75794 10337 76526 10383
rect 75794 10334 75806 10337
rect 76514 10334 76526 10337
rect 76578 10334 76590 10386
rect 55134 10322 55186 10334
rect 1344 10218 78624 10252
rect 1344 10166 10874 10218
rect 10926 10166 10978 10218
rect 11030 10166 11082 10218
rect 11134 10166 30194 10218
rect 30246 10166 30298 10218
rect 30350 10166 30402 10218
rect 30454 10166 49514 10218
rect 49566 10166 49618 10218
rect 49670 10166 49722 10218
rect 49774 10166 68834 10218
rect 68886 10166 68938 10218
rect 68990 10166 69042 10218
rect 69094 10166 78624 10218
rect 1344 10132 78624 10166
rect 16830 10050 16882 10062
rect 21310 10050 21362 10062
rect 17378 9998 17390 10050
rect 17442 10047 17454 10050
rect 17938 10047 17950 10050
rect 17442 10001 17950 10047
rect 17442 9998 17454 10001
rect 17938 9998 17950 10001
rect 18002 9998 18014 10050
rect 16830 9986 16882 9998
rect 21310 9986 21362 9998
rect 45278 10050 45330 10062
rect 45278 9986 45330 9998
rect 51662 10050 51714 10062
rect 51662 9986 51714 9998
rect 6190 9938 6242 9950
rect 16718 9938 16770 9950
rect 7410 9886 7422 9938
rect 7474 9886 7486 9938
rect 9538 9886 9550 9938
rect 9602 9886 9614 9938
rect 12786 9886 12798 9938
rect 12850 9886 12862 9938
rect 14242 9886 14254 9938
rect 14306 9886 14318 9938
rect 16370 9886 16382 9938
rect 16434 9886 16446 9938
rect 6190 9874 6242 9886
rect 16718 9874 16770 9886
rect 17390 9938 17442 9950
rect 17390 9874 17442 9886
rect 21422 9938 21474 9950
rect 21422 9874 21474 9886
rect 21870 9938 21922 9950
rect 21870 9874 21922 9886
rect 22766 9938 22818 9950
rect 22766 9874 22818 9886
rect 24894 9938 24946 9950
rect 24894 9874 24946 9886
rect 25342 9938 25394 9950
rect 25342 9874 25394 9886
rect 25790 9938 25842 9950
rect 25790 9874 25842 9886
rect 31950 9938 32002 9950
rect 42590 9938 42642 9950
rect 33730 9886 33742 9938
rect 33794 9886 33806 9938
rect 35858 9886 35870 9938
rect 35922 9886 35934 9938
rect 37202 9886 37214 9938
rect 37266 9886 37278 9938
rect 41234 9886 41246 9938
rect 41298 9886 41310 9938
rect 31950 9874 32002 9886
rect 42590 9874 42642 9886
rect 43150 9938 43202 9950
rect 53454 9938 53506 9950
rect 48290 9886 48302 9938
rect 48354 9886 48366 9938
rect 50418 9886 50430 9938
rect 50482 9886 50494 9938
rect 54786 9886 54798 9938
rect 54850 9886 54862 9938
rect 56914 9886 56926 9938
rect 56978 9886 56990 9938
rect 61842 9886 61854 9938
rect 61906 9886 61918 9938
rect 63970 9886 63982 9938
rect 64034 9886 64046 9938
rect 65426 9886 65438 9938
rect 65490 9886 65502 9938
rect 69234 9886 69246 9938
rect 69298 9886 69310 9938
rect 71362 9886 71374 9938
rect 71426 9886 71438 9938
rect 43150 9874 43202 9886
rect 53454 9874 53506 9886
rect 4174 9826 4226 9838
rect 5742 9826 5794 9838
rect 19854 9826 19906 9838
rect 20414 9826 20466 9838
rect 4722 9774 4734 9826
rect 4786 9774 4798 9826
rect 10322 9774 10334 9826
rect 10386 9774 10398 9826
rect 12450 9774 12462 9826
rect 12514 9774 12526 9826
rect 13570 9774 13582 9826
rect 13634 9774 13646 9826
rect 20178 9774 20190 9826
rect 20242 9774 20254 9826
rect 4174 9762 4226 9774
rect 5742 9762 5794 9774
rect 19854 9762 19906 9774
rect 20414 9762 20466 9774
rect 20750 9826 20802 9838
rect 20750 9762 20802 9774
rect 31166 9826 31218 9838
rect 46734 9826 46786 9838
rect 71710 9826 71762 9838
rect 32946 9774 32958 9826
rect 33010 9774 33022 9826
rect 37538 9774 37550 9826
rect 37602 9774 37614 9826
rect 38322 9774 38334 9826
rect 38386 9774 38398 9826
rect 46050 9774 46062 9826
rect 46114 9774 46126 9826
rect 47506 9774 47518 9826
rect 47570 9774 47582 9826
rect 52882 9774 52894 9826
rect 52946 9774 52958 9826
rect 54002 9774 54014 9826
rect 54066 9774 54078 9826
rect 61058 9774 61070 9826
rect 61122 9774 61134 9826
rect 68562 9774 68574 9826
rect 68626 9774 68638 9826
rect 31166 9762 31218 9774
rect 46734 9762 46786 9774
rect 71710 9762 71762 9774
rect 72830 9826 72882 9838
rect 72830 9762 72882 9774
rect 73502 9826 73554 9838
rect 76414 9826 76466 9838
rect 74274 9774 74286 9826
rect 74338 9774 74350 9826
rect 73502 9762 73554 9774
rect 76414 9762 76466 9774
rect 3166 9714 3218 9726
rect 3166 9650 3218 9662
rect 3838 9714 3890 9726
rect 17838 9714 17890 9726
rect 4946 9662 4958 9714
rect 5010 9662 5022 9714
rect 3838 9650 3890 9662
rect 17838 9650 17890 9662
rect 19294 9714 19346 9726
rect 19294 9650 19346 9662
rect 19630 9714 19682 9726
rect 19630 9650 19682 9662
rect 26574 9714 26626 9726
rect 26574 9650 26626 9662
rect 31390 9714 31442 9726
rect 31390 9650 31442 9662
rect 31502 9714 31554 9726
rect 31502 9650 31554 9662
rect 32398 9714 32450 9726
rect 47070 9714 47122 9726
rect 57822 9714 57874 9726
rect 39106 9662 39118 9714
rect 39170 9662 39182 9714
rect 45938 9662 45950 9714
rect 46002 9662 46014 9714
rect 51090 9662 51102 9714
rect 51154 9662 51166 9714
rect 51314 9662 51326 9714
rect 51378 9662 51390 9714
rect 32398 9650 32450 9662
rect 47070 9650 47122 9662
rect 57822 9650 57874 9662
rect 64990 9714 65042 9726
rect 64990 9650 65042 9662
rect 65886 9714 65938 9726
rect 65886 9650 65938 9662
rect 66558 9714 66610 9726
rect 73838 9714 73890 9726
rect 72034 9662 72046 9714
rect 72098 9662 72110 9714
rect 66558 9650 66610 9662
rect 73838 9650 73890 9662
rect 77086 9714 77138 9726
rect 77086 9650 77138 9662
rect 2830 9602 2882 9614
rect 2830 9538 2882 9550
rect 12126 9602 12178 9614
rect 12126 9538 12178 9550
rect 19742 9602 19794 9614
rect 19742 9538 19794 9550
rect 20638 9602 20690 9614
rect 20638 9538 20690 9550
rect 26910 9602 26962 9614
rect 26910 9538 26962 9550
rect 41694 9602 41746 9614
rect 41694 9538 41746 9550
rect 43598 9602 43650 9614
rect 43598 9538 43650 9550
rect 44942 9602 44994 9614
rect 44942 9538 44994 9550
rect 51998 9602 52050 9614
rect 51998 9538 52050 9550
rect 52670 9602 52722 9614
rect 52670 9538 52722 9550
rect 57486 9602 57538 9614
rect 57486 9538 57538 9550
rect 66222 9602 66274 9614
rect 66222 9538 66274 9550
rect 73278 9602 73330 9614
rect 73278 9538 73330 9550
rect 73390 9602 73442 9614
rect 73390 9538 73442 9550
rect 76750 9602 76802 9614
rect 76750 9538 76802 9550
rect 1344 9434 78784 9468
rect 1344 9382 20534 9434
rect 20586 9382 20638 9434
rect 20690 9382 20742 9434
rect 20794 9382 39854 9434
rect 39906 9382 39958 9434
rect 40010 9382 40062 9434
rect 40114 9382 59174 9434
rect 59226 9382 59278 9434
rect 59330 9382 59382 9434
rect 59434 9382 78494 9434
rect 78546 9382 78598 9434
rect 78650 9382 78702 9434
rect 78754 9382 78784 9434
rect 1344 9348 78784 9382
rect 6638 9266 6690 9278
rect 6638 9202 6690 9214
rect 7086 9266 7138 9278
rect 7870 9266 7922 9278
rect 7522 9214 7534 9266
rect 7586 9214 7598 9266
rect 7086 9202 7138 9214
rect 7870 9202 7922 9214
rect 9662 9266 9714 9278
rect 9662 9202 9714 9214
rect 13246 9266 13298 9278
rect 13246 9202 13298 9214
rect 14926 9266 14978 9278
rect 14926 9202 14978 9214
rect 34526 9266 34578 9278
rect 34526 9202 34578 9214
rect 39118 9266 39170 9278
rect 39118 9202 39170 9214
rect 49646 9266 49698 9278
rect 49646 9202 49698 9214
rect 56030 9266 56082 9278
rect 56030 9202 56082 9214
rect 61294 9266 61346 9278
rect 61294 9202 61346 9214
rect 61966 9266 62018 9278
rect 61966 9202 62018 9214
rect 68574 9266 68626 9278
rect 68574 9202 68626 9214
rect 68798 9266 68850 9278
rect 68798 9202 68850 9214
rect 69582 9266 69634 9278
rect 69582 9202 69634 9214
rect 69806 9266 69858 9278
rect 69806 9202 69858 9214
rect 71374 9266 71426 9278
rect 71374 9202 71426 9214
rect 72382 9266 72434 9278
rect 72382 9202 72434 9214
rect 73614 9266 73666 9278
rect 73614 9202 73666 9214
rect 73950 9266 74002 9278
rect 73950 9202 74002 9214
rect 8430 9154 8482 9166
rect 11454 9154 11506 9166
rect 13470 9154 13522 9166
rect 5170 9102 5182 9154
rect 5234 9102 5246 9154
rect 5506 9102 5518 9154
rect 5570 9102 5582 9154
rect 10770 9102 10782 9154
rect 10834 9102 10846 9154
rect 12338 9102 12350 9154
rect 12402 9102 12414 9154
rect 12674 9102 12686 9154
rect 12738 9102 12750 9154
rect 8430 9090 8482 9102
rect 11454 9090 11506 9102
rect 13470 9090 13522 9102
rect 13582 9154 13634 9166
rect 13582 9090 13634 9102
rect 14030 9154 14082 9166
rect 22990 9154 23042 9166
rect 30494 9154 30546 9166
rect 38446 9154 38498 9166
rect 48750 9154 48802 9166
rect 19506 9102 19518 9154
rect 19570 9102 19582 9154
rect 26898 9102 26910 9154
rect 26962 9102 26974 9154
rect 35410 9102 35422 9154
rect 35474 9102 35486 9154
rect 47170 9102 47182 9154
rect 47234 9102 47246 9154
rect 47506 9102 47518 9154
rect 47570 9102 47582 9154
rect 52546 9102 52558 9154
rect 52610 9102 52622 9154
rect 57586 9102 57598 9154
rect 57650 9102 57662 9154
rect 62514 9102 62526 9154
rect 62578 9102 62590 9154
rect 63074 9102 63086 9154
rect 63138 9102 63150 9154
rect 63522 9102 63534 9154
rect 63586 9102 63598 9154
rect 65762 9102 65774 9154
rect 65826 9102 65838 9154
rect 14030 9090 14082 9102
rect 22990 9090 23042 9102
rect 30494 9090 30546 9102
rect 38446 9090 38498 9102
rect 48750 9090 48802 9102
rect 5742 9042 5794 9054
rect 4274 8990 4286 9042
rect 4338 8990 4350 9042
rect 5742 8978 5794 8990
rect 8990 9042 9042 9054
rect 23326 9042 23378 9054
rect 30830 9042 30882 9054
rect 10658 8990 10670 9042
rect 10722 8990 10734 9042
rect 18834 8990 18846 9042
rect 18898 8990 18910 9042
rect 26114 8990 26126 9042
rect 26178 8990 26190 9042
rect 8990 8978 9042 8990
rect 23326 8978 23378 8990
rect 30830 8978 30882 8990
rect 34862 9042 34914 9054
rect 36206 9042 36258 9054
rect 47742 9042 47794 9054
rect 35634 8990 35646 9042
rect 35698 8990 35710 9042
rect 38658 8990 38670 9042
rect 38722 8990 38734 9042
rect 39330 8990 39342 9042
rect 39394 8990 39406 9042
rect 46162 8990 46174 9042
rect 46226 8990 46238 9042
rect 34862 8978 34914 8990
rect 36206 8978 36258 8990
rect 47742 8978 47794 8990
rect 48078 9042 48130 9054
rect 62302 9042 62354 9054
rect 69918 9042 69970 9054
rect 48962 8990 48974 9042
rect 49026 8990 49038 9042
rect 53218 8990 53230 9042
rect 53282 8990 53294 9042
rect 56802 8990 56814 9042
rect 56866 8990 56878 9042
rect 63746 8990 63758 9042
rect 63810 8990 63822 9042
rect 65090 8990 65102 9042
rect 65154 8990 65166 9042
rect 48078 8978 48130 8990
rect 62302 8978 62354 8990
rect 69918 8978 69970 8990
rect 70366 9042 70418 9054
rect 70366 8978 70418 8990
rect 72270 9042 72322 9054
rect 72270 8978 72322 8990
rect 72606 9042 72658 9054
rect 76066 8990 76078 9042
rect 76130 8990 76142 9042
rect 72606 8978 72658 8990
rect 34078 8930 34130 8942
rect 21634 8878 21646 8930
rect 21698 8878 21710 8930
rect 29026 8878 29038 8930
rect 29090 8878 29102 8930
rect 34078 8866 34130 8878
rect 37998 8930 38050 8942
rect 60846 8930 60898 8942
rect 72942 8930 72994 8942
rect 43250 8878 43262 8930
rect 43314 8878 43326 8930
rect 45378 8878 45390 8930
rect 45442 8878 45454 8930
rect 37998 8866 38050 8878
rect 50418 8851 50430 8903
rect 50482 8851 50494 8903
rect 59714 8878 59726 8930
rect 59778 8878 59790 8930
rect 67890 8878 67902 8930
rect 67954 8878 67966 8930
rect 69234 8878 69246 8930
rect 69298 8878 69310 8930
rect 60846 8866 60898 8878
rect 72942 8866 72994 8878
rect 1934 8818 1986 8830
rect 1934 8754 1986 8766
rect 6078 8818 6130 8830
rect 6078 8754 6130 8766
rect 9998 8818 10050 8830
rect 9998 8754 10050 8766
rect 11790 8818 11842 8830
rect 11790 8754 11842 8766
rect 12126 8818 12178 8830
rect 12126 8754 12178 8766
rect 77982 8818 78034 8830
rect 77982 8754 78034 8766
rect 1344 8650 78624 8684
rect 1344 8598 10874 8650
rect 10926 8598 10978 8650
rect 11030 8598 11082 8650
rect 11134 8598 30194 8650
rect 30246 8598 30298 8650
rect 30350 8598 30402 8650
rect 30454 8598 49514 8650
rect 49566 8598 49618 8650
rect 49670 8598 49722 8650
rect 49774 8598 68834 8650
rect 68886 8598 68938 8650
rect 68990 8598 69042 8650
rect 69094 8598 78624 8650
rect 1344 8564 78624 8598
rect 26462 8482 26514 8494
rect 26462 8418 26514 8430
rect 57822 8482 57874 8494
rect 5182 8370 5234 8382
rect 2482 8318 2494 8370
rect 2546 8318 2558 8370
rect 4610 8318 4622 8370
rect 4674 8318 4686 8370
rect 5182 8306 5234 8318
rect 9214 8370 9266 8382
rect 14030 8370 14082 8382
rect 18286 8370 18338 8382
rect 21422 8370 21474 8382
rect 32498 8374 32510 8426
rect 32562 8374 32574 8426
rect 57822 8418 57874 8430
rect 66558 8482 66610 8494
rect 66558 8418 66610 8430
rect 34414 8370 34466 8382
rect 12674 8318 12686 8370
rect 12738 8318 12750 8370
rect 17490 8318 17502 8370
rect 17554 8318 17566 8370
rect 19842 8318 19854 8370
rect 19906 8318 19918 8370
rect 22754 8318 22766 8370
rect 22818 8318 22830 8370
rect 24882 8318 24894 8370
rect 24946 8318 24958 8370
rect 30370 8318 30382 8370
rect 30434 8318 30446 8370
rect 9214 8306 9266 8318
rect 14030 8306 14082 8318
rect 18286 8306 18338 8318
rect 21422 8306 21474 8318
rect 34414 8306 34466 8318
rect 40574 8370 40626 8382
rect 49422 8370 49474 8382
rect 47282 8318 47294 8370
rect 47346 8318 47358 8370
rect 40574 8306 40626 8318
rect 49422 8306 49474 8318
rect 58158 8370 58210 8382
rect 58158 8306 58210 8318
rect 63310 8370 63362 8382
rect 63310 8306 63362 8318
rect 66222 8370 66274 8382
rect 66222 8306 66274 8318
rect 67118 8370 67170 8382
rect 73602 8318 73614 8370
rect 73666 8318 73678 8370
rect 67118 8306 67170 8318
rect 5966 8258 6018 8270
rect 20750 8258 20802 8270
rect 26798 8258 26850 8270
rect 28142 8258 28194 8270
rect 37438 8258 37490 8270
rect 56702 8258 56754 8270
rect 1810 8206 1822 8258
rect 1874 8206 1886 8258
rect 9874 8206 9886 8258
rect 9938 8206 9950 8258
rect 14578 8206 14590 8258
rect 14642 8206 14654 8258
rect 19058 8206 19070 8258
rect 19122 8206 19134 8258
rect 20066 8206 20078 8258
rect 20130 8206 20142 8258
rect 21970 8206 21982 8258
rect 22034 8206 22046 8258
rect 27458 8206 27470 8258
rect 27522 8206 27534 8258
rect 29698 8206 29710 8258
rect 29762 8206 29774 8258
rect 34962 8206 34974 8258
rect 35026 8206 35038 8258
rect 35634 8206 35646 8258
rect 35698 8206 35710 8258
rect 38210 8206 38222 8258
rect 38274 8206 38286 8258
rect 44930 8206 44942 8258
rect 44994 8206 45006 8258
rect 46498 8206 46510 8258
rect 46562 8206 46574 8258
rect 65650 8206 65662 8258
rect 65714 8206 65726 8258
rect 70690 8206 70702 8258
rect 70754 8206 70766 8258
rect 5966 8194 6018 8206
rect 20750 8194 20802 8206
rect 26798 8194 26850 8206
rect 28142 8194 28194 8206
rect 37438 8194 37490 8206
rect 56702 8194 56754 8206
rect 20414 8146 20466 8158
rect 37102 8146 37154 8158
rect 39566 8146 39618 8158
rect 10546 8094 10558 8146
rect 10610 8094 10622 8146
rect 15362 8094 15374 8146
rect 15426 8094 15438 8146
rect 18834 8094 18846 8146
rect 18898 8094 18910 8146
rect 20178 8094 20190 8146
rect 20242 8094 20254 8146
rect 27346 8094 27358 8146
rect 27410 8094 27422 8146
rect 38098 8094 38110 8146
rect 38162 8094 38174 8146
rect 20414 8082 20466 8094
rect 37102 8082 37154 8094
rect 39566 8082 39618 8094
rect 45166 8146 45218 8158
rect 45166 8082 45218 8094
rect 57150 8146 57202 8158
rect 58370 8094 58382 8146
rect 58434 8094 58446 8146
rect 58706 8094 58718 8146
rect 58770 8094 58782 8146
rect 65538 8094 65550 8146
rect 65602 8094 65614 8146
rect 71474 8094 71486 8146
rect 71538 8094 71550 8146
rect 57150 8082 57202 8094
rect 5630 8034 5682 8046
rect 5630 7970 5682 7982
rect 13582 8034 13634 8046
rect 13582 7970 13634 7982
rect 17950 8034 18002 8046
rect 17950 7970 18002 7982
rect 20638 8034 20690 8046
rect 20638 7970 20690 7982
rect 26014 8034 26066 8046
rect 35870 8034 35922 8046
rect 34738 7982 34750 8034
rect 34802 7982 34814 8034
rect 26014 7970 26066 7982
rect 35870 7970 35922 7982
rect 38782 8034 38834 8046
rect 38782 7970 38834 7982
rect 39902 8034 39954 8046
rect 39902 7970 39954 7982
rect 55246 8034 55298 8046
rect 55246 7970 55298 7982
rect 69806 8034 69858 8046
rect 69806 7970 69858 7982
rect 70366 8034 70418 8046
rect 70366 7970 70418 7982
rect 1344 7866 78784 7900
rect 1344 7814 20534 7866
rect 20586 7814 20638 7866
rect 20690 7814 20742 7866
rect 20794 7814 39854 7866
rect 39906 7814 39958 7866
rect 40010 7814 40062 7866
rect 40114 7814 59174 7866
rect 59226 7814 59278 7866
rect 59330 7814 59382 7866
rect 59434 7814 78494 7866
rect 78546 7814 78598 7866
rect 78650 7814 78702 7866
rect 78754 7814 78784 7866
rect 1344 7780 78784 7814
rect 9662 7698 9714 7710
rect 9662 7634 9714 7646
rect 10782 7698 10834 7710
rect 10782 7634 10834 7646
rect 15598 7698 15650 7710
rect 15598 7634 15650 7646
rect 17502 7698 17554 7710
rect 17502 7634 17554 7646
rect 19518 7698 19570 7710
rect 19518 7634 19570 7646
rect 20526 7698 20578 7710
rect 20526 7634 20578 7646
rect 23438 7698 23490 7710
rect 23438 7634 23490 7646
rect 25342 7698 25394 7710
rect 25342 7634 25394 7646
rect 31054 7698 31106 7710
rect 31054 7634 31106 7646
rect 33182 7698 33234 7710
rect 33182 7634 33234 7646
rect 41022 7698 41074 7710
rect 41022 7634 41074 7646
rect 41470 7698 41522 7710
rect 41470 7634 41522 7646
rect 44606 7698 44658 7710
rect 44606 7634 44658 7646
rect 72382 7698 72434 7710
rect 72382 7634 72434 7646
rect 72494 7698 72546 7710
rect 72494 7634 72546 7646
rect 72718 7698 72770 7710
rect 72718 7634 72770 7646
rect 2382 7586 2434 7598
rect 2382 7522 2434 7534
rect 2718 7586 2770 7598
rect 11118 7586 11170 7598
rect 3826 7534 3838 7586
rect 3890 7534 3902 7586
rect 8642 7534 8654 7586
rect 8706 7534 8718 7586
rect 2718 7522 2770 7534
rect 11118 7522 11170 7534
rect 15934 7586 15986 7598
rect 25902 7586 25954 7598
rect 42590 7586 42642 7598
rect 62974 7586 63026 7598
rect 23986 7534 23998 7586
rect 24050 7534 24062 7586
rect 24322 7534 24334 7586
rect 24386 7534 24398 7586
rect 31714 7534 31726 7586
rect 31778 7534 31790 7586
rect 32162 7534 32174 7586
rect 32226 7534 32238 7586
rect 36530 7534 36542 7586
rect 36594 7534 36606 7586
rect 40114 7534 40126 7586
rect 40178 7534 40190 7586
rect 43922 7534 43934 7586
rect 43986 7534 43998 7586
rect 55570 7534 55582 7586
rect 55634 7534 55646 7586
rect 15934 7522 15986 7534
rect 25902 7522 25954 7534
rect 42590 7522 42642 7534
rect 62974 7522 63026 7534
rect 69694 7586 69746 7598
rect 69694 7522 69746 7534
rect 70366 7586 70418 7598
rect 70366 7522 70418 7534
rect 76750 7586 76802 7598
rect 76750 7522 76802 7534
rect 8094 7474 8146 7486
rect 23774 7474 23826 7486
rect 3042 7422 3054 7474
rect 3106 7422 3118 7474
rect 8866 7422 8878 7474
rect 8930 7422 8942 7474
rect 8094 7410 8146 7422
rect 23774 7410 23826 7422
rect 31390 7474 31442 7486
rect 39454 7474 39506 7486
rect 62638 7474 62690 7486
rect 70702 7474 70754 7486
rect 72270 7474 72322 7486
rect 37314 7422 37326 7474
rect 37378 7422 37390 7474
rect 40226 7422 40238 7474
rect 40290 7422 40302 7474
rect 44034 7422 44046 7474
rect 44098 7422 44110 7474
rect 52434 7422 52446 7474
rect 52498 7422 52510 7474
rect 55794 7422 55806 7474
rect 55858 7422 55870 7474
rect 69906 7422 69918 7474
rect 69970 7422 69982 7474
rect 71138 7422 71150 7474
rect 71202 7422 71214 7474
rect 76962 7422 76974 7474
rect 77026 7422 77038 7474
rect 31390 7410 31442 7422
rect 39454 7410 39506 7422
rect 62638 7410 62690 7422
rect 70702 7410 70754 7422
rect 72270 7410 72322 7422
rect 7422 7362 7474 7374
rect 68910 7362 68962 7374
rect 5954 7310 5966 7362
rect 6018 7310 6030 7362
rect 34402 7310 34414 7362
rect 34466 7310 34478 7362
rect 53106 7310 53118 7362
rect 53170 7310 53182 7362
rect 55234 7310 55246 7362
rect 55298 7310 55310 7362
rect 7422 7298 7474 7310
rect 68910 7298 68962 7310
rect 69246 7362 69298 7374
rect 73278 7362 73330 7374
rect 71474 7310 71486 7362
rect 71538 7310 71550 7362
rect 69246 7298 69298 7310
rect 73278 7298 73330 7310
rect 76526 7362 76578 7374
rect 76526 7298 76578 7310
rect 7758 7250 7810 7262
rect 7758 7186 7810 7198
rect 39118 7250 39170 7262
rect 39118 7186 39170 7198
rect 42926 7250 42978 7262
rect 42926 7186 42978 7198
rect 43262 7250 43314 7262
rect 43262 7186 43314 7198
rect 1344 7082 78624 7116
rect 1344 7030 10874 7082
rect 10926 7030 10978 7082
rect 11030 7030 11082 7082
rect 11134 7030 30194 7082
rect 30246 7030 30298 7082
rect 30350 7030 30402 7082
rect 30454 7030 49514 7082
rect 49566 7030 49618 7082
rect 49670 7030 49722 7082
rect 49774 7030 68834 7082
rect 68886 7030 68938 7082
rect 68990 7030 69042 7082
rect 69094 7030 78624 7082
rect 1344 6996 78624 7030
rect 48974 6914 49026 6926
rect 48974 6850 49026 6862
rect 54686 6914 54738 6926
rect 54686 6850 54738 6862
rect 58830 6914 58882 6926
rect 59490 6862 59502 6914
rect 59554 6911 59566 6914
rect 60050 6911 60062 6914
rect 59554 6865 60062 6911
rect 59554 6862 59566 6865
rect 60050 6862 60062 6865
rect 60114 6862 60126 6914
rect 58830 6850 58882 6862
rect 14254 6802 14306 6814
rect 14254 6738 14306 6750
rect 25006 6802 25058 6814
rect 25006 6738 25058 6750
rect 28142 6802 28194 6814
rect 39666 6750 39678 6802
rect 39730 6750 39742 6802
rect 41906 6750 41918 6802
rect 41970 6750 41982 6802
rect 61954 6750 61966 6802
rect 62018 6750 62030 6802
rect 28142 6738 28194 6750
rect 4846 6690 4898 6702
rect 4274 6638 4286 6690
rect 4338 6638 4350 6690
rect 4846 6626 4898 6638
rect 11342 6690 11394 6702
rect 32622 6690 32674 6702
rect 42926 6690 42978 6702
rect 13682 6638 13694 6690
rect 13746 6638 13758 6690
rect 25554 6638 25566 6690
rect 25618 6638 25630 6690
rect 38994 6638 39006 6690
rect 39058 6638 39070 6690
rect 11342 6626 11394 6638
rect 32622 6626 32674 6638
rect 42926 6626 42978 6638
rect 43262 6690 43314 6702
rect 56030 6690 56082 6702
rect 55458 6638 55470 6690
rect 55522 6638 55534 6690
rect 43262 6626 43314 6638
rect 56030 6626 56082 6638
rect 57262 6690 57314 6702
rect 59166 6690 59218 6702
rect 65326 6690 65378 6702
rect 58258 6638 58270 6690
rect 58322 6638 58334 6690
rect 64082 6638 64094 6690
rect 64146 6638 64158 6690
rect 64866 6638 64878 6690
rect 64930 6638 64942 6690
rect 57262 6626 57314 6638
rect 59166 6626 59218 6638
rect 65326 6626 65378 6638
rect 66222 6690 66274 6702
rect 66222 6626 66274 6638
rect 69694 6690 69746 6702
rect 69694 6626 69746 6638
rect 70702 6690 70754 6702
rect 70702 6626 70754 6638
rect 71710 6690 71762 6702
rect 71710 6626 71762 6638
rect 11006 6578 11058 6590
rect 2482 6526 2494 6578
rect 2546 6526 2558 6578
rect 11006 6514 11058 6526
rect 20078 6578 20130 6590
rect 20078 6514 20130 6526
rect 20414 6578 20466 6590
rect 20414 6514 20466 6526
rect 21646 6578 21698 6590
rect 21646 6514 21698 6526
rect 26574 6578 26626 6590
rect 26574 6514 26626 6526
rect 26910 6578 26962 6590
rect 35758 6578 35810 6590
rect 27458 6526 27470 6578
rect 27522 6526 27534 6578
rect 27906 6526 27918 6578
rect 27970 6526 27982 6578
rect 26910 6514 26962 6526
rect 35758 6514 35810 6526
rect 36094 6578 36146 6590
rect 50430 6578 50482 6590
rect 49186 6526 49198 6578
rect 49250 6526 49262 6578
rect 49746 6526 49758 6578
rect 49810 6526 49822 6578
rect 36094 6514 36146 6526
rect 50430 6514 50482 6526
rect 53342 6578 53394 6590
rect 53342 6514 53394 6526
rect 53678 6578 53730 6590
rect 53678 6514 53730 6526
rect 54350 6578 54402 6590
rect 65662 6578 65714 6590
rect 55234 6526 55246 6578
rect 55298 6526 55310 6578
rect 58034 6526 58046 6578
rect 58098 6526 58110 6578
rect 54350 6514 54402 6526
rect 65662 6514 65714 6526
rect 68686 6578 68738 6590
rect 68686 6514 68738 6526
rect 69022 6578 69074 6590
rect 69022 6514 69074 6526
rect 70926 6578 70978 6590
rect 70926 6514 70978 6526
rect 71262 6578 71314 6590
rect 71262 6514 71314 6526
rect 21310 6466 21362 6478
rect 28478 6466 28530 6478
rect 13458 6414 13470 6466
rect 13522 6414 13534 6466
rect 25330 6414 25342 6466
rect 25394 6414 25406 6466
rect 21310 6402 21362 6414
rect 28478 6402 28530 6414
rect 29374 6466 29426 6478
rect 29374 6402 29426 6414
rect 35422 6466 35474 6478
rect 35422 6402 35474 6414
rect 43598 6466 43650 6478
rect 43598 6402 43650 6414
rect 48638 6466 48690 6478
rect 48638 6402 48690 6414
rect 57598 6466 57650 6478
rect 57598 6402 57650 6414
rect 59726 6466 59778 6478
rect 59726 6402 59778 6414
rect 60622 6466 60674 6478
rect 60622 6402 60674 6414
rect 61742 6466 61794 6478
rect 61742 6402 61794 6414
rect 67342 6466 67394 6478
rect 67342 6402 67394 6414
rect 69358 6466 69410 6478
rect 69358 6402 69410 6414
rect 70030 6466 70082 6478
rect 70030 6402 70082 6414
rect 70142 6466 70194 6478
rect 70142 6402 70194 6414
rect 70254 6466 70306 6478
rect 70254 6402 70306 6414
rect 72270 6466 72322 6478
rect 72270 6402 72322 6414
rect 72606 6466 72658 6478
rect 72606 6402 72658 6414
rect 1344 6298 78784 6332
rect 1344 6246 20534 6298
rect 20586 6246 20638 6298
rect 20690 6246 20742 6298
rect 20794 6246 39854 6298
rect 39906 6246 39958 6298
rect 40010 6246 40062 6298
rect 40114 6246 59174 6298
rect 59226 6246 59278 6298
rect 59330 6246 59382 6298
rect 59434 6246 78494 6298
rect 78546 6246 78598 6298
rect 78650 6246 78702 6298
rect 78754 6246 78784 6298
rect 1344 6212 78784 6246
rect 10110 6130 10162 6142
rect 13134 6130 13186 6142
rect 10770 6078 10782 6130
rect 10834 6078 10846 6130
rect 10110 6066 10162 6078
rect 13134 6066 13186 6078
rect 14254 6130 14306 6142
rect 14254 6066 14306 6078
rect 19742 6130 19794 6142
rect 19742 6066 19794 6078
rect 21310 6130 21362 6142
rect 21310 6066 21362 6078
rect 26014 6130 26066 6142
rect 26014 6066 26066 6078
rect 36206 6130 36258 6142
rect 36206 6066 36258 6078
rect 37102 6130 37154 6142
rect 37102 6066 37154 6078
rect 37998 6130 38050 6142
rect 37998 6066 38050 6078
rect 42702 6130 42754 6142
rect 55358 6130 55410 6142
rect 51762 6078 51774 6130
rect 51826 6078 51838 6130
rect 42702 6066 42754 6078
rect 55358 6066 55410 6078
rect 55694 6130 55746 6142
rect 62638 6130 62690 6142
rect 71374 6130 71426 6142
rect 56578 6078 56590 6130
rect 56642 6078 56654 6130
rect 67106 6078 67118 6130
rect 67170 6078 67182 6130
rect 55694 6066 55746 6078
rect 62638 6066 62690 6078
rect 71374 6066 71426 6078
rect 72158 6130 72210 6142
rect 72158 6066 72210 6078
rect 72382 6130 72434 6142
rect 72382 6066 72434 6078
rect 72942 6130 72994 6142
rect 72942 6066 72994 6078
rect 73390 6130 73442 6142
rect 73390 6066 73442 6078
rect 11118 6018 11170 6030
rect 15822 6018 15874 6030
rect 12450 5966 12462 6018
rect 12514 5966 12526 6018
rect 11118 5954 11170 5966
rect 15822 5954 15874 5966
rect 16158 6018 16210 6030
rect 16158 5954 16210 5966
rect 16830 6018 16882 6030
rect 20414 6018 20466 6030
rect 18498 5966 18510 6018
rect 18562 5966 18574 6018
rect 16830 5954 16882 5966
rect 20414 5954 20466 5966
rect 21982 6018 22034 6030
rect 32174 6018 32226 6030
rect 23426 5966 23438 6018
rect 23490 5966 23502 6018
rect 21982 5954 22034 5966
rect 32174 5954 32226 5966
rect 32510 6018 32562 6030
rect 32510 5954 32562 5966
rect 33294 6018 33346 6030
rect 37438 6018 37490 6030
rect 48190 6018 48242 6030
rect 56030 6018 56082 6030
rect 61742 6018 61794 6030
rect 66334 6018 66386 6030
rect 35186 5966 35198 6018
rect 35250 5966 35262 6018
rect 42354 5966 42366 6018
rect 42418 5966 42430 6018
rect 43810 5966 43822 6018
rect 43874 5966 43886 6018
rect 49522 5966 49534 6018
rect 49586 5966 49598 6018
rect 58146 5966 58158 6018
rect 58210 5966 58222 6018
rect 63186 5966 63198 6018
rect 63250 5966 63262 6018
rect 63522 5966 63534 6018
rect 63586 5966 63598 6018
rect 65650 5966 65662 6018
rect 65714 5966 65726 6018
rect 33294 5954 33346 5966
rect 37438 5954 37490 5966
rect 48190 5954 48242 5966
rect 56030 5954 56082 5966
rect 61742 5954 61794 5966
rect 66334 5954 66386 5966
rect 14590 5906 14642 5918
rect 17838 5906 17890 5918
rect 26350 5906 26402 5918
rect 33630 5906 33682 5918
rect 8978 5854 8990 5906
rect 9042 5854 9054 5906
rect 10322 5854 10334 5906
rect 10386 5854 10398 5906
rect 12674 5854 12686 5906
rect 12738 5854 12750 5906
rect 16594 5854 16606 5906
rect 16658 5854 16670 5906
rect 18386 5854 18398 5906
rect 18450 5854 18462 5906
rect 19954 5854 19966 5906
rect 20018 5854 20030 5906
rect 20626 5854 20638 5906
rect 20690 5854 20702 5906
rect 21746 5854 21758 5906
rect 21810 5854 21822 5906
rect 23538 5854 23550 5906
rect 23602 5854 23614 5906
rect 29474 5854 29486 5906
rect 29538 5854 29550 5906
rect 14590 5842 14642 5854
rect 17838 5842 17890 5854
rect 26350 5842 26402 5854
rect 33630 5842 33682 5854
rect 34302 5906 34354 5918
rect 34302 5842 34354 5854
rect 34638 5906 34690 5918
rect 56926 5906 56978 5918
rect 60846 5906 60898 5918
rect 35298 5854 35310 5906
rect 35362 5854 35374 5906
rect 43026 5854 43038 5906
rect 43090 5854 43102 5906
rect 47954 5854 47966 5906
rect 48018 5854 48030 5906
rect 48850 5854 48862 5906
rect 48914 5854 48926 5906
rect 57474 5854 57486 5906
rect 57538 5854 57550 5906
rect 34638 5842 34690 5854
rect 56926 5842 56978 5854
rect 60846 5842 60898 5854
rect 62078 5906 62130 5918
rect 62078 5842 62130 5854
rect 62974 5906 63026 5918
rect 62974 5842 63026 5854
rect 65438 5906 65490 5918
rect 66670 5906 66722 5918
rect 72494 5906 72546 5918
rect 65874 5854 65886 5906
rect 65938 5854 65950 5906
rect 70018 5854 70030 5906
rect 70082 5854 70094 5906
rect 70578 5854 70590 5906
rect 70642 5854 70654 5906
rect 71586 5854 71598 5906
rect 71650 5854 71662 5906
rect 76066 5854 76078 5906
rect 76130 5854 76142 5906
rect 65438 5842 65490 5854
rect 66670 5842 66722 5854
rect 72494 5842 72546 5854
rect 15038 5794 15090 5806
rect 6066 5742 6078 5794
rect 6130 5742 6142 5794
rect 8194 5742 8206 5794
rect 8258 5742 8270 5794
rect 13570 5742 13582 5794
rect 13634 5742 13646 5794
rect 15038 5730 15090 5742
rect 19294 5794 19346 5806
rect 19294 5730 19346 5742
rect 24222 5794 24274 5806
rect 38670 5794 38722 5806
rect 55022 5794 55074 5806
rect 61406 5794 61458 5806
rect 77982 5794 78034 5806
rect 26674 5742 26686 5794
rect 26738 5742 26750 5794
rect 28802 5742 28814 5794
rect 28866 5742 28878 5794
rect 36642 5742 36654 5794
rect 36706 5742 36718 5794
rect 45938 5742 45950 5794
rect 46002 5742 46014 5794
rect 60274 5742 60286 5794
rect 60338 5742 60350 5794
rect 69346 5742 69358 5794
rect 69410 5742 69422 5794
rect 70914 5742 70926 5794
rect 70978 5742 70990 5794
rect 24222 5730 24274 5742
rect 38670 5730 38722 5742
rect 55022 5730 55074 5742
rect 61406 5730 61458 5742
rect 77982 5730 78034 5742
rect 11566 5682 11618 5694
rect 11566 5618 11618 5630
rect 11902 5682 11954 5694
rect 11902 5618 11954 5630
rect 17502 5682 17554 5694
rect 17502 5618 17554 5630
rect 22430 5682 22482 5694
rect 22430 5618 22482 5630
rect 22766 5682 22818 5694
rect 55010 5630 55022 5682
rect 55074 5679 55086 5682
rect 55346 5679 55358 5682
rect 55074 5633 55358 5679
rect 55074 5630 55086 5633
rect 55346 5630 55358 5633
rect 55410 5630 55422 5682
rect 22766 5618 22818 5630
rect 1344 5514 78624 5548
rect 1344 5462 10874 5514
rect 10926 5462 10978 5514
rect 11030 5462 11082 5514
rect 11134 5462 30194 5514
rect 30246 5462 30298 5514
rect 30350 5462 30402 5514
rect 30454 5462 49514 5514
rect 49566 5462 49618 5514
rect 49670 5462 49722 5514
rect 49774 5462 68834 5514
rect 68886 5462 68938 5514
rect 68990 5462 69042 5514
rect 69094 5462 78624 5514
rect 1344 5428 78624 5462
rect 45278 5346 45330 5358
rect 45278 5282 45330 5294
rect 54574 5346 54626 5358
rect 54574 5282 54626 5294
rect 62190 5346 62242 5358
rect 62190 5282 62242 5294
rect 62526 5346 62578 5358
rect 62526 5282 62578 5294
rect 66670 5346 66722 5358
rect 66670 5282 66722 5294
rect 13918 5234 13970 5246
rect 37438 5234 37490 5246
rect 46622 5234 46674 5246
rect 12898 5182 12910 5234
rect 12962 5182 12974 5234
rect 17042 5182 17054 5234
rect 17106 5182 17118 5234
rect 19170 5182 19182 5234
rect 19234 5182 19246 5234
rect 22194 5182 22206 5234
rect 22258 5182 22270 5234
rect 24322 5182 24334 5234
rect 24386 5182 24398 5234
rect 28466 5182 28478 5234
rect 28530 5182 28542 5234
rect 32722 5182 32734 5234
rect 32786 5182 32798 5234
rect 34850 5182 34862 5234
rect 34914 5182 34926 5234
rect 41794 5182 41806 5234
rect 41858 5182 41870 5234
rect 13918 5170 13970 5182
rect 37438 5170 37490 5182
rect 46622 5170 46674 5182
rect 47070 5234 47122 5246
rect 47070 5170 47122 5182
rect 50654 5234 50706 5246
rect 50654 5170 50706 5182
rect 59390 5234 59442 5246
rect 59390 5170 59442 5182
rect 59950 5234 60002 5246
rect 59950 5170 60002 5182
rect 68462 5234 68514 5246
rect 76974 5234 77026 5246
rect 70242 5182 70254 5234
rect 70306 5182 70318 5234
rect 72482 5182 72494 5234
rect 72546 5182 72558 5234
rect 68462 5170 68514 5182
rect 76974 5170 77026 5182
rect 15710 5122 15762 5134
rect 20750 5122 20802 5134
rect 29486 5122 29538 5134
rect 37102 5122 37154 5134
rect 44270 5122 44322 5134
rect 7522 5070 7534 5122
rect 7586 5070 7598 5122
rect 8978 5070 8990 5122
rect 9042 5070 9054 5122
rect 9986 5070 9998 5122
rect 10050 5070 10062 5122
rect 14690 5070 14702 5122
rect 14754 5070 14766 5122
rect 16258 5070 16270 5122
rect 16322 5070 16334 5122
rect 21522 5070 21534 5122
rect 21586 5070 21598 5122
rect 25666 5070 25678 5122
rect 25730 5070 25742 5122
rect 31938 5070 31950 5122
rect 32002 5070 32014 5122
rect 35410 5070 35422 5122
rect 35474 5070 35486 5122
rect 36194 5070 36206 5122
rect 36258 5070 36270 5122
rect 38210 5070 38222 5122
rect 38274 5070 38286 5122
rect 38994 5070 39006 5122
rect 39058 5070 39070 5122
rect 42690 5070 42702 5122
rect 42754 5070 42766 5122
rect 15710 5058 15762 5070
rect 20750 5058 20802 5070
rect 29486 5058 29538 5070
rect 37102 5058 37154 5070
rect 44270 5058 44322 5070
rect 44942 5122 44994 5134
rect 53006 5122 53058 5134
rect 54238 5122 54290 5134
rect 55918 5122 55970 5134
rect 57822 5122 57874 5134
rect 45714 5070 45726 5122
rect 45778 5070 45790 5122
rect 47842 5070 47854 5122
rect 47906 5070 47918 5122
rect 53554 5070 53566 5122
rect 53618 5070 53630 5122
rect 55346 5070 55358 5122
rect 55410 5070 55422 5122
rect 57138 5070 57150 5122
rect 57202 5070 57214 5122
rect 44942 5058 44994 5070
rect 53006 5058 53058 5070
rect 54238 5058 54290 5070
rect 55918 5058 55970 5070
rect 57822 5058 57874 5070
rect 58158 5122 58210 5134
rect 61182 5122 61234 5134
rect 63870 5122 63922 5134
rect 58818 5070 58830 5122
rect 58882 5070 58894 5122
rect 60722 5070 60734 5122
rect 60786 5070 60798 5122
rect 61618 5070 61630 5122
rect 61682 5070 61694 5122
rect 62962 5070 62974 5122
rect 63026 5070 63038 5122
rect 58158 5058 58210 5070
rect 61182 5058 61234 5070
rect 63870 5058 63922 5070
rect 65102 5122 65154 5134
rect 66334 5122 66386 5134
rect 65762 5070 65774 5122
rect 65826 5070 65838 5122
rect 65102 5058 65154 5070
rect 66334 5058 66386 5070
rect 67230 5122 67282 5134
rect 67230 5058 67282 5070
rect 67566 5122 67618 5134
rect 67566 5058 67618 5070
rect 67902 5122 67954 5134
rect 67902 5058 67954 5070
rect 68350 5122 68402 5134
rect 68350 5058 68402 5070
rect 69022 5122 69074 5134
rect 75742 5122 75794 5134
rect 69570 5070 69582 5122
rect 69634 5070 69646 5122
rect 69022 5058 69074 5070
rect 75742 5058 75794 5070
rect 76414 5122 76466 5134
rect 76414 5058 76466 5070
rect 7758 5010 7810 5022
rect 29150 5010 29202 5022
rect 10770 4958 10782 5010
rect 10834 4958 10846 5010
rect 14466 4958 14478 5010
rect 14530 4958 14542 5010
rect 26338 4958 26350 5010
rect 26402 4958 26414 5010
rect 7758 4946 7810 4958
rect 29150 4946 29202 4958
rect 31614 5010 31666 5022
rect 31614 4946 31666 4958
rect 35982 5010 36034 5022
rect 43262 5010 43314 5022
rect 38098 4958 38110 5010
rect 38162 4958 38174 5010
rect 39666 4958 39678 5010
rect 39730 4958 39742 5010
rect 35982 4946 36034 4958
rect 43262 4946 43314 4958
rect 43598 5010 43650 5022
rect 52670 5010 52722 5022
rect 60510 5010 60562 5022
rect 64766 5010 64818 5022
rect 67678 5010 67730 5022
rect 43922 4958 43934 5010
rect 43986 4958 43998 5010
rect 46050 4958 46062 5010
rect 46114 4958 46126 5010
rect 48514 4958 48526 5010
rect 48578 4958 48590 5010
rect 55234 4958 55246 5010
rect 55298 4958 55310 5010
rect 56242 4958 56254 5010
rect 56306 4958 56318 5010
rect 57250 4958 57262 5010
rect 57314 4958 57326 5010
rect 63298 4958 63310 5010
rect 63362 4958 63374 5010
rect 65538 4958 65550 5010
rect 65602 4958 65614 5010
rect 43598 4946 43650 4958
rect 52670 4946 52722 4958
rect 60510 4946 60562 4958
rect 64766 4946 64818 4958
rect 67678 4946 67730 4958
rect 68574 5010 68626 5022
rect 68574 4946 68626 4958
rect 9214 4898 9266 4910
rect 9214 4834 9266 4846
rect 13582 4898 13634 4910
rect 13582 4834 13634 4846
rect 15374 4898 15426 4910
rect 15374 4834 15426 4846
rect 20414 4898 20466 4910
rect 20414 4834 20466 4846
rect 31278 4898 31330 4910
rect 31278 4834 31330 4846
rect 35646 4898 35698 4910
rect 35646 4834 35698 4846
rect 42926 4898 42978 4910
rect 42926 4834 42978 4846
rect 53342 4898 53394 4910
rect 53342 4834 53394 4846
rect 58606 4898 58658 4910
rect 58606 4834 58658 4846
rect 1344 4730 78784 4764
rect 1344 4678 20534 4730
rect 20586 4678 20638 4730
rect 20690 4678 20742 4730
rect 20794 4678 39854 4730
rect 39906 4678 39958 4730
rect 40010 4678 40062 4730
rect 40114 4678 59174 4730
rect 59226 4678 59278 4730
rect 59330 4678 59382 4730
rect 59434 4678 78494 4730
rect 78546 4678 78598 4730
rect 78650 4678 78702 4730
rect 78754 4678 78784 4730
rect 1344 4644 78784 4678
rect 12798 4562 12850 4574
rect 12798 4498 12850 4510
rect 17614 4562 17666 4574
rect 17614 4498 17666 4510
rect 23326 4562 23378 4574
rect 23326 4498 23378 4510
rect 26126 4562 26178 4574
rect 26126 4498 26178 4510
rect 33294 4562 33346 4574
rect 33294 4498 33346 4510
rect 35086 4562 35138 4574
rect 35086 4498 35138 4510
rect 40014 4562 40066 4574
rect 40014 4498 40066 4510
rect 42814 4562 42866 4574
rect 42814 4498 42866 4510
rect 48190 4562 48242 4574
rect 48190 4498 48242 4510
rect 50654 4562 50706 4574
rect 50654 4498 50706 4510
rect 13134 4450 13186 4462
rect 25790 4450 25842 4462
rect 56030 4450 56082 4462
rect 10322 4398 10334 4450
rect 10386 4398 10398 4450
rect 14690 4398 14702 4450
rect 14754 4398 14766 4450
rect 18498 4398 18510 4450
rect 18562 4398 18574 4450
rect 20626 4398 20638 4450
rect 20690 4398 20702 4450
rect 23874 4398 23886 4450
rect 23938 4398 23950 4450
rect 24434 4398 24446 4450
rect 24498 4398 24510 4450
rect 27794 4398 27806 4450
rect 27858 4398 27870 4450
rect 30370 4398 30382 4450
rect 30434 4398 30446 4450
rect 34178 4398 34190 4450
rect 34242 4398 34254 4450
rect 37650 4398 37662 4450
rect 37714 4398 37726 4450
rect 42130 4398 42142 4450
rect 42194 4398 42206 4450
rect 44370 4398 44382 4450
rect 44434 4398 44446 4450
rect 49410 4398 49422 4450
rect 49474 4398 49486 4450
rect 49858 4398 49870 4450
rect 49922 4398 49934 4450
rect 52994 4398 53006 4450
rect 53058 4398 53070 4450
rect 57362 4398 57374 4450
rect 57426 4398 57438 4450
rect 61394 4398 61406 4450
rect 61458 4398 61470 4450
rect 65986 4398 65998 4450
rect 66050 4398 66062 4450
rect 13134 4386 13186 4398
rect 25790 4386 25842 4398
rect 56030 4386 56082 4398
rect 17950 4338 18002 4350
rect 19406 4338 19458 4350
rect 23662 4338 23714 4350
rect 4274 4286 4286 4338
rect 4338 4286 4350 4338
rect 9650 4286 9662 4338
rect 9714 4286 9726 4338
rect 14018 4286 14030 4338
rect 14082 4286 14094 4338
rect 18722 4286 18734 4338
rect 18786 4286 18798 4338
rect 19842 4286 19854 4338
rect 19906 4286 19918 4338
rect 17950 4274 18002 4286
rect 19406 4274 19458 4286
rect 23662 4274 23714 4286
rect 25454 4338 25506 4350
rect 25454 4274 25506 4286
rect 26462 4338 26514 4350
rect 26462 4274 26514 4286
rect 26910 4338 26962 4350
rect 26910 4274 26962 4286
rect 27246 4338 27298 4350
rect 33630 4338 33682 4350
rect 40350 4338 40402 4350
rect 28018 4286 28030 4338
rect 28082 4286 28094 4338
rect 29698 4286 29710 4338
rect 29762 4286 29774 4338
rect 34402 4286 34414 4338
rect 34466 4286 34478 4338
rect 38434 4286 38446 4338
rect 38498 4286 38510 4338
rect 27246 4274 27298 4286
rect 33630 4274 33682 4286
rect 40350 4274 40402 4286
rect 41022 4338 41074 4350
rect 41022 4274 41074 4286
rect 41358 4338 41410 4350
rect 48862 4338 48914 4350
rect 42018 4286 42030 4338
rect 42082 4286 42094 4338
rect 43698 4286 43710 4338
rect 43762 4286 43774 4338
rect 47954 4286 47966 4338
rect 48018 4286 48030 4338
rect 41358 4274 41410 4286
rect 48862 4274 48914 4286
rect 49198 4338 49250 4350
rect 52322 4286 52334 4338
rect 52386 4286 52398 4338
rect 55794 4286 55806 4338
rect 55858 4286 55870 4338
rect 56578 4286 56590 4338
rect 56642 4286 56654 4338
rect 60610 4286 60622 4338
rect 60674 4286 60686 4338
rect 65202 4286 65214 4338
rect 65266 4286 65278 4338
rect 68674 4286 68686 4338
rect 68738 4286 68750 4338
rect 75618 4286 75630 4338
rect 75682 4286 75694 4338
rect 49198 4274 49250 4286
rect 4734 4226 4786 4238
rect 4734 4162 4786 4174
rect 5182 4226 5234 4238
rect 46510 4226 46562 4238
rect 59502 4226 59554 4238
rect 12450 4174 12462 4226
rect 12514 4174 12526 4226
rect 16818 4174 16830 4226
rect 16882 4174 16894 4226
rect 22754 4174 22766 4226
rect 22818 4174 22830 4226
rect 32498 4174 32510 4226
rect 32562 4174 32574 4226
rect 35522 4174 35534 4226
rect 35586 4174 35598 4226
rect 55122 4174 55134 4226
rect 55186 4174 55198 4226
rect 63522 4174 63534 4226
rect 63586 4174 63598 4226
rect 68114 4174 68126 4226
rect 68178 4174 68190 4226
rect 5182 4162 5234 4174
rect 46510 4162 46562 4174
rect 59502 4162 59554 4174
rect 1934 4114 1986 4126
rect 1934 4050 1986 4062
rect 69470 4114 69522 4126
rect 69470 4050 69522 4062
rect 77982 4114 78034 4126
rect 77982 4050 78034 4062
rect 1344 3946 78624 3980
rect 1344 3894 10874 3946
rect 10926 3894 10978 3946
rect 11030 3894 11082 3946
rect 11134 3894 30194 3946
rect 30246 3894 30298 3946
rect 30350 3894 30402 3946
rect 30454 3894 49514 3946
rect 49566 3894 49618 3946
rect 49670 3894 49722 3946
rect 49774 3894 68834 3946
rect 68886 3894 68938 3946
rect 68990 3894 69042 3946
rect 69094 3894 78624 3946
rect 1344 3860 78624 3894
rect 1934 3666 1986 3678
rect 1934 3602 1986 3614
rect 5742 3666 5794 3678
rect 5742 3602 5794 3614
rect 36878 3666 36930 3678
rect 36878 3602 36930 3614
rect 57038 3666 57090 3678
rect 67118 3666 67170 3678
rect 64754 3614 64766 3666
rect 64818 3614 64830 3666
rect 57038 3602 57090 3614
rect 67118 3602 67170 3614
rect 68350 3666 68402 3678
rect 68350 3602 68402 3614
rect 68686 3666 68738 3678
rect 68686 3602 68738 3614
rect 20302 3554 20354 3566
rect 67902 3554 67954 3566
rect 4274 3502 4286 3554
rect 4338 3502 4350 3554
rect 4722 3502 4734 3554
rect 4786 3502 4798 3554
rect 20962 3502 20974 3554
rect 21026 3502 21038 3554
rect 24770 3502 24782 3554
rect 24834 3502 24846 3554
rect 72594 3502 72606 3554
rect 72658 3502 72670 3554
rect 77186 3502 77198 3554
rect 77250 3502 77262 3554
rect 20302 3490 20354 3502
rect 67902 3490 67954 3502
rect 4958 3442 5010 3454
rect 4958 3378 5010 3390
rect 7646 3442 7698 3454
rect 7646 3378 7698 3390
rect 7870 3442 7922 3454
rect 7870 3378 7922 3390
rect 8206 3442 8258 3454
rect 8206 3378 8258 3390
rect 11678 3442 11730 3454
rect 11678 3378 11730 3390
rect 11902 3442 11954 3454
rect 11902 3378 11954 3390
rect 12238 3442 12290 3454
rect 12238 3378 12290 3390
rect 15710 3442 15762 3454
rect 15710 3378 15762 3390
rect 15934 3442 15986 3454
rect 15934 3378 15986 3390
rect 16270 3442 16322 3454
rect 16270 3378 16322 3390
rect 20750 3442 20802 3454
rect 20750 3378 20802 3390
rect 24110 3442 24162 3454
rect 24110 3378 24162 3390
rect 27918 3442 27970 3454
rect 27918 3378 27970 3390
rect 28366 3442 28418 3454
rect 28366 3378 28418 3390
rect 28702 3442 28754 3454
rect 28702 3378 28754 3390
rect 31726 3442 31778 3454
rect 31726 3378 31778 3390
rect 32174 3442 32226 3454
rect 32174 3378 32226 3390
rect 32510 3442 32562 3454
rect 32510 3378 32562 3390
rect 35534 3442 35586 3454
rect 35534 3378 35586 3390
rect 36094 3442 36146 3454
rect 36094 3378 36146 3390
rect 36430 3442 36482 3454
rect 36430 3378 36482 3390
rect 39342 3442 39394 3454
rect 39342 3378 39394 3390
rect 40126 3442 40178 3454
rect 40126 3378 40178 3390
rect 40462 3442 40514 3454
rect 40462 3378 40514 3390
rect 43934 3442 43986 3454
rect 43934 3378 43986 3390
rect 44158 3442 44210 3454
rect 44158 3378 44210 3390
rect 44494 3442 44546 3454
rect 44494 3378 44546 3390
rect 47966 3442 48018 3454
rect 47966 3378 48018 3390
rect 48190 3442 48242 3454
rect 48190 3378 48242 3390
rect 48526 3442 48578 3454
rect 48526 3378 48578 3390
rect 51998 3442 52050 3454
rect 51998 3378 52050 3390
rect 52222 3442 52274 3454
rect 52222 3378 52274 3390
rect 52558 3442 52610 3454
rect 52558 3378 52610 3390
rect 56030 3442 56082 3454
rect 56030 3378 56082 3390
rect 56254 3442 56306 3454
rect 56254 3378 56306 3390
rect 56590 3442 56642 3454
rect 56590 3378 56642 3390
rect 60062 3442 60114 3454
rect 60062 3378 60114 3390
rect 60286 3442 60338 3454
rect 60286 3378 60338 3390
rect 60622 3442 60674 3454
rect 60622 3378 60674 3390
rect 64094 3442 64146 3454
rect 64094 3378 64146 3390
rect 64318 3442 64370 3454
rect 64318 3378 64370 3390
rect 72158 3442 72210 3454
rect 75506 3390 75518 3442
rect 75570 3390 75582 3442
rect 72158 3378 72210 3390
rect 24558 3330 24610 3342
rect 24558 3266 24610 3278
rect 72382 3330 72434 3342
rect 72382 3266 72434 3278
rect 1344 3162 78784 3196
rect 1344 3110 20534 3162
rect 20586 3110 20638 3162
rect 20690 3110 20742 3162
rect 20794 3110 39854 3162
rect 39906 3110 39958 3162
rect 40010 3110 40062 3162
rect 40114 3110 59174 3162
rect 59226 3110 59278 3162
rect 59330 3110 59382 3162
rect 59434 3110 78494 3162
rect 78546 3110 78598 3162
rect 78650 3110 78702 3162
rect 78754 3110 78784 3162
rect 1344 3076 78784 3110
<< via1 >>
rect 10874 36822 10926 36874
rect 10978 36822 11030 36874
rect 11082 36822 11134 36874
rect 30194 36822 30246 36874
rect 30298 36822 30350 36874
rect 30402 36822 30454 36874
rect 49514 36822 49566 36874
rect 49618 36822 49670 36874
rect 49722 36822 49774 36874
rect 68834 36822 68886 36874
rect 68938 36822 68990 36874
rect 69042 36822 69094 36874
rect 43934 36654 43986 36706
rect 47630 36654 47682 36706
rect 56030 36654 56082 36706
rect 64094 36654 64146 36706
rect 71822 36654 71874 36706
rect 75070 36654 75122 36706
rect 1934 36542 1986 36594
rect 6526 36542 6578 36594
rect 8878 36542 8930 36594
rect 11454 36542 11506 36594
rect 13918 36542 13970 36594
rect 16382 36542 16434 36594
rect 18846 36542 18898 36594
rect 19630 36542 19682 36594
rect 21310 36542 21362 36594
rect 22094 36542 22146 36594
rect 23662 36542 23714 36594
rect 26350 36542 26402 36594
rect 31166 36542 31218 36594
rect 31614 36542 31666 36594
rect 34862 36542 34914 36594
rect 35534 36542 35586 36594
rect 38446 36542 38498 36594
rect 41022 36542 41074 36594
rect 3950 36430 4002 36482
rect 6750 36430 6802 36482
rect 9326 36430 9378 36482
rect 11678 36430 11730 36482
rect 14142 36430 14194 36482
rect 17054 36430 17106 36482
rect 19070 36430 19122 36482
rect 21534 36430 21586 36482
rect 24558 36430 24610 36482
rect 25118 36430 25170 36482
rect 27358 36430 27410 36482
rect 29150 36430 29202 36482
rect 30718 36430 30770 36482
rect 32846 36430 32898 36482
rect 33854 36430 33906 36482
rect 34414 36430 34466 36482
rect 36542 36430 36594 36482
rect 38670 36430 38722 36482
rect 39230 36430 39282 36482
rect 43038 36430 43090 36482
rect 46286 36430 46338 36482
rect 49870 36430 49922 36482
rect 53678 36430 53730 36482
rect 55022 36430 55074 36482
rect 58942 36430 58994 36482
rect 62638 36430 62690 36482
rect 66558 36430 66610 36482
rect 70814 36430 70866 36482
rect 74062 36430 74114 36482
rect 7310 36318 7362 36370
rect 9886 36318 9938 36370
rect 12238 36318 12290 36370
rect 14478 36318 14530 36370
rect 24110 36318 24162 36370
rect 27022 36318 27074 36370
rect 29822 36318 29874 36370
rect 30382 36318 30434 36370
rect 32510 36318 32562 36370
rect 52110 36318 52162 36370
rect 60622 36318 60674 36370
rect 17278 36206 17330 36258
rect 17726 36206 17778 36258
rect 25902 36206 25954 36258
rect 26686 36206 26738 36258
rect 27694 36206 27746 36258
rect 28702 36206 28754 36258
rect 28926 36206 28978 36258
rect 30494 36206 30546 36258
rect 32174 36206 32226 36258
rect 33182 36206 33234 36258
rect 36318 36206 36370 36258
rect 40014 36206 40066 36258
rect 46846 36206 46898 36258
rect 50430 36206 50482 36258
rect 65886 36206 65938 36258
rect 67454 36206 67506 36258
rect 70478 36206 70530 36258
rect 20534 36038 20586 36090
rect 20638 36038 20690 36090
rect 20742 36038 20794 36090
rect 39854 36038 39906 36090
rect 39958 36038 40010 36090
rect 40062 36038 40114 36090
rect 59174 36038 59226 36090
rect 59278 36038 59330 36090
rect 59382 36038 59434 36090
rect 78494 36038 78546 36090
rect 78598 36038 78650 36090
rect 78702 36038 78754 36090
rect 3278 35870 3330 35922
rect 4622 35870 4674 35922
rect 24782 35870 24834 35922
rect 28254 35870 28306 35922
rect 30382 35870 30434 35922
rect 65438 35870 65490 35922
rect 76638 35870 76690 35922
rect 17726 35758 17778 35810
rect 28814 35758 28866 35810
rect 37214 35758 37266 35810
rect 38222 35758 38274 35810
rect 48190 35758 48242 35810
rect 48974 35758 49026 35810
rect 50654 35758 50706 35810
rect 54574 35758 54626 35810
rect 63870 35758 63922 35810
rect 67342 35758 67394 35810
rect 71262 35758 71314 35810
rect 4286 35646 4338 35698
rect 10334 35646 10386 35698
rect 13806 35646 13858 35698
rect 17614 35646 17666 35698
rect 19294 35646 19346 35698
rect 25342 35646 25394 35698
rect 29038 35646 29090 35698
rect 29486 35646 29538 35698
rect 30158 35646 30210 35698
rect 31278 35646 31330 35698
rect 32398 35646 32450 35698
rect 33294 35646 33346 35698
rect 36878 35646 36930 35698
rect 38782 35646 38834 35698
rect 45054 35646 45106 35698
rect 46286 35646 46338 35698
rect 47630 35646 47682 35698
rect 47966 35646 48018 35698
rect 48862 35646 48914 35698
rect 49086 35646 49138 35698
rect 50430 35646 50482 35698
rect 50990 35646 51042 35698
rect 51326 35646 51378 35698
rect 54910 35646 54962 35698
rect 60958 35646 61010 35698
rect 64430 35646 64482 35698
rect 67678 35646 67730 35698
rect 68350 35646 68402 35698
rect 71598 35646 71650 35698
rect 73166 35646 73218 35698
rect 76078 35646 76130 35698
rect 5182 35534 5234 35586
rect 11006 35534 11058 35586
rect 13246 35534 13298 35586
rect 14478 35534 14530 35586
rect 16606 35534 16658 35586
rect 18286 35534 18338 35586
rect 19070 35534 19122 35586
rect 20078 35534 20130 35586
rect 22318 35534 22370 35586
rect 23662 35534 23714 35586
rect 26014 35534 26066 35586
rect 28702 35534 28754 35586
rect 30830 35534 30882 35586
rect 31950 35534 32002 35586
rect 33070 35534 33122 35586
rect 35422 35534 35474 35586
rect 36542 35534 36594 35586
rect 37774 35534 37826 35586
rect 39118 35534 39170 35586
rect 39902 35534 39954 35586
rect 42142 35534 42194 35586
rect 44270 35534 44322 35586
rect 45614 35534 45666 35586
rect 46958 35534 47010 35586
rect 47742 35534 47794 35586
rect 52110 35534 52162 35586
rect 54238 35534 54290 35586
rect 55358 35534 55410 35586
rect 58046 35534 58098 35586
rect 60286 35534 60338 35586
rect 69358 35534 69410 35586
rect 72494 35534 72546 35586
rect 75070 35534 75122 35586
rect 17726 35422 17778 35474
rect 29710 35422 29762 35474
rect 30494 35422 30546 35474
rect 33518 35422 33570 35474
rect 33966 35422 34018 35474
rect 37886 35422 37938 35474
rect 40014 35422 40066 35474
rect 45502 35422 45554 35474
rect 49534 35422 49586 35474
rect 10874 35254 10926 35306
rect 10978 35254 11030 35306
rect 11082 35254 11134 35306
rect 30194 35254 30246 35306
rect 30298 35254 30350 35306
rect 30402 35254 30454 35306
rect 49514 35254 49566 35306
rect 49618 35254 49670 35306
rect 49722 35254 49774 35306
rect 68834 35254 68886 35306
rect 68938 35254 68990 35306
rect 69042 35254 69094 35306
rect 2942 35086 2994 35138
rect 25454 35086 25506 35138
rect 40574 35086 40626 35138
rect 44382 35086 44434 35138
rect 3502 34974 3554 35026
rect 4398 34974 4450 35026
rect 13582 34974 13634 35026
rect 14254 34974 14306 35026
rect 14702 34974 14754 35026
rect 17726 34974 17778 35026
rect 18398 34974 18450 35026
rect 18958 34974 19010 35026
rect 33518 34974 33570 35026
rect 43038 34974 43090 35026
rect 44942 34974 44994 35026
rect 45390 34974 45442 35026
rect 46398 34974 46450 35026
rect 52110 34974 52162 35026
rect 53902 34974 53954 35026
rect 57262 34974 57314 35026
rect 67678 34974 67730 35026
rect 68574 34974 68626 35026
rect 73054 34974 73106 35026
rect 73726 34974 73778 35026
rect 1822 34862 1874 34914
rect 2382 34862 2434 34914
rect 15374 34862 15426 34914
rect 16270 34862 16322 34914
rect 16494 34862 16546 34914
rect 17054 34862 17106 34914
rect 18062 34862 18114 34914
rect 21534 34862 21586 34914
rect 26574 34862 26626 34914
rect 26798 34862 26850 34914
rect 28366 34862 28418 34914
rect 29486 34862 29538 34914
rect 30046 34862 30098 34914
rect 30830 34862 30882 34914
rect 31166 34862 31218 34914
rect 32846 34862 32898 34914
rect 33854 34862 33906 34914
rect 34526 34862 34578 34914
rect 34750 34862 34802 34914
rect 35870 34862 35922 34914
rect 36206 34862 36258 34914
rect 37326 34862 37378 34914
rect 37774 34862 37826 34914
rect 38446 34862 38498 34914
rect 39342 34862 39394 34914
rect 40350 34862 40402 34914
rect 40574 34862 40626 34914
rect 43710 34862 43762 34914
rect 45614 34862 45666 34914
rect 45950 34862 46002 34914
rect 47630 34862 47682 34914
rect 47966 34862 48018 34914
rect 49198 34862 49250 34914
rect 54350 34862 54402 34914
rect 60622 34862 60674 34914
rect 64766 34862 64818 34914
rect 70142 34862 70194 34914
rect 3054 34750 3106 34802
rect 15710 34750 15762 34802
rect 22206 34750 22258 34802
rect 25342 34750 25394 34802
rect 25902 34750 25954 34802
rect 27358 34750 27410 34802
rect 27470 34750 27522 34802
rect 29710 34750 29762 34802
rect 34302 34750 34354 34802
rect 38558 34750 38610 34802
rect 42590 34750 42642 34802
rect 43486 34750 43538 34802
rect 44046 34750 44098 34802
rect 44270 34750 44322 34802
rect 45726 34750 45778 34802
rect 46958 34750 47010 34802
rect 49982 34750 50034 34802
rect 55134 34750 55186 34802
rect 57598 34750 57650 34802
rect 57934 34750 57986 34802
rect 61294 34750 61346 34802
rect 65550 34750 65602 34802
rect 70926 34750 70978 34802
rect 4734 34638 4786 34690
rect 15598 34638 15650 34690
rect 15934 34638 15986 34690
rect 24446 34638 24498 34690
rect 25006 34638 25058 34690
rect 27134 34638 27186 34690
rect 28030 34638 28082 34690
rect 28590 34638 28642 34690
rect 29598 34638 29650 34690
rect 35758 34638 35810 34690
rect 36430 34638 36482 34690
rect 36542 34638 36594 34690
rect 39342 34638 39394 34690
rect 41134 34638 41186 34690
rect 54014 34638 54066 34690
rect 63534 34638 63586 34690
rect 75406 34638 75458 34690
rect 76302 34638 76354 34690
rect 20534 34470 20586 34522
rect 20638 34470 20690 34522
rect 20742 34470 20794 34522
rect 39854 34470 39906 34522
rect 39958 34470 40010 34522
rect 40062 34470 40114 34522
rect 59174 34470 59226 34522
rect 59278 34470 59330 34522
rect 59382 34470 59434 34522
rect 78494 34470 78546 34522
rect 78598 34470 78650 34522
rect 78702 34470 78754 34522
rect 13918 34302 13970 34354
rect 16942 34302 16994 34354
rect 20414 34302 20466 34354
rect 24222 34302 24274 34354
rect 26350 34302 26402 34354
rect 27134 34302 27186 34354
rect 27694 34302 27746 34354
rect 29374 34302 29426 34354
rect 33070 34302 33122 34354
rect 33294 34302 33346 34354
rect 41246 34302 41298 34354
rect 41918 34302 41970 34354
rect 44158 34302 44210 34354
rect 48078 34302 48130 34354
rect 55582 34302 55634 34354
rect 58158 34302 58210 34354
rect 65326 34302 65378 34354
rect 24446 34190 24498 34242
rect 28814 34190 28866 34242
rect 43486 34190 43538 34242
rect 44718 34190 44770 34242
rect 45838 34190 45890 34242
rect 58830 34190 58882 34242
rect 60062 34190 60114 34242
rect 66446 34190 66498 34242
rect 70030 34190 70082 34242
rect 71038 34190 71090 34242
rect 71374 34190 71426 34242
rect 4286 34078 4338 34130
rect 11006 34078 11058 34130
rect 14814 34078 14866 34130
rect 15374 34078 15426 34130
rect 17838 34078 17890 34130
rect 18286 34078 18338 34130
rect 20526 34078 20578 34130
rect 22990 34078 23042 34130
rect 23438 34078 23490 34130
rect 23886 34078 23938 34130
rect 24110 34078 24162 34130
rect 25902 34078 25954 34130
rect 26798 34078 26850 34130
rect 28926 34078 28978 34130
rect 29486 34078 29538 34130
rect 29822 34078 29874 34130
rect 32062 34078 32114 34130
rect 33182 34078 33234 34130
rect 33742 34078 33794 34130
rect 33966 34078 34018 34130
rect 34302 34078 34354 34130
rect 36542 34078 36594 34130
rect 36990 34078 37042 34130
rect 40126 34078 40178 34130
rect 40798 34078 40850 34130
rect 41470 34078 41522 34130
rect 41694 34078 41746 34130
rect 42030 34078 42082 34130
rect 44382 34078 44434 34130
rect 45166 34078 45218 34130
rect 49422 34078 49474 34130
rect 53678 34078 53730 34130
rect 54126 34078 54178 34130
rect 54462 34078 54514 34130
rect 57262 34078 57314 34130
rect 58046 34078 58098 34130
rect 59054 34078 59106 34130
rect 60398 34078 60450 34130
rect 60734 34078 60786 34130
rect 65102 34078 65154 34130
rect 65662 34078 65714 34130
rect 69694 34078 69746 34130
rect 70478 34078 70530 34130
rect 70814 34078 70866 34130
rect 73166 34078 73218 34130
rect 75630 34078 75682 34130
rect 4846 33966 4898 34018
rect 11678 33966 11730 34018
rect 15934 33966 15986 34018
rect 18510 33966 18562 34018
rect 19518 33966 19570 34018
rect 21870 33966 21922 34018
rect 25342 33966 25394 34018
rect 27918 33966 27970 34018
rect 28030 33966 28082 34018
rect 29710 33966 29762 34018
rect 29934 33966 29986 34018
rect 31950 33966 32002 34018
rect 36094 33966 36146 34018
rect 37438 33966 37490 34018
rect 39678 33966 39730 34018
rect 41358 33966 41410 34018
rect 48750 33966 48802 34018
rect 49198 33966 49250 34018
rect 51326 33966 51378 34018
rect 54014 33966 54066 34018
rect 55358 33966 55410 34018
rect 55470 33966 55522 34018
rect 57150 33966 57202 34018
rect 61518 33966 61570 34018
rect 63646 33966 63698 34018
rect 68574 33966 68626 34018
rect 69358 33966 69410 34018
rect 73950 33966 74002 34018
rect 1934 33854 1986 33906
rect 32398 33854 32450 33906
rect 38894 33854 38946 33906
rect 56926 33854 56978 33906
rect 77982 33854 78034 33906
rect 10874 33686 10926 33738
rect 10978 33686 11030 33738
rect 11082 33686 11134 33738
rect 30194 33686 30246 33738
rect 30298 33686 30350 33738
rect 30402 33686 30454 33738
rect 49514 33686 49566 33738
rect 49618 33686 49670 33738
rect 49722 33686 49774 33738
rect 68834 33686 68886 33738
rect 68938 33686 68990 33738
rect 69042 33686 69094 33738
rect 12574 33518 12626 33570
rect 15150 33518 15202 33570
rect 15710 33518 15762 33570
rect 29262 33518 29314 33570
rect 31502 33518 31554 33570
rect 35870 33518 35922 33570
rect 37102 33518 37154 33570
rect 48862 33518 48914 33570
rect 56030 33518 56082 33570
rect 57150 33518 57202 33570
rect 61966 33518 62018 33570
rect 66446 33518 66498 33570
rect 3278 33406 3330 33458
rect 13470 33406 13522 33458
rect 19742 33406 19794 33458
rect 21422 33406 21474 33458
rect 23662 33406 23714 33458
rect 24782 33406 24834 33458
rect 25454 33406 25506 33458
rect 27246 33406 27298 33458
rect 31390 33406 31442 33458
rect 32398 33406 32450 33458
rect 33966 33406 34018 33458
rect 36206 33406 36258 33458
rect 38334 33406 38386 33458
rect 43486 33406 43538 33458
rect 44830 33406 44882 33458
rect 45390 33406 45442 33458
rect 55358 33406 55410 33458
rect 70814 33406 70866 33458
rect 72942 33406 72994 33458
rect 14478 33294 14530 33346
rect 14814 33294 14866 33346
rect 15150 33294 15202 33346
rect 15710 33294 15762 33346
rect 18958 33294 19010 33346
rect 19294 33294 19346 33346
rect 22094 33294 22146 33346
rect 23550 33294 23602 33346
rect 25342 33294 25394 33346
rect 26686 33294 26738 33346
rect 28254 33294 28306 33346
rect 29374 33294 29426 33346
rect 30382 33294 30434 33346
rect 33854 33294 33906 33346
rect 37214 33294 37266 33346
rect 37774 33294 37826 33346
rect 39454 33294 39506 33346
rect 40798 33294 40850 33346
rect 45054 33294 45106 33346
rect 45838 33294 45890 33346
rect 49198 33294 49250 33346
rect 51662 33294 51714 33346
rect 51998 33294 52050 33346
rect 54910 33294 54962 33346
rect 55806 33294 55858 33346
rect 56366 33294 56418 33346
rect 58046 33294 58098 33346
rect 58158 33294 58210 33346
rect 58382 33294 58434 33346
rect 59054 33294 59106 33346
rect 59278 33294 59330 33346
rect 61070 33294 61122 33346
rect 66782 33294 66834 33346
rect 70030 33294 70082 33346
rect 12686 33182 12738 33234
rect 13582 33182 13634 33234
rect 16046 33182 16098 33234
rect 16270 33182 16322 33234
rect 18622 33182 18674 33234
rect 18734 33182 18786 33234
rect 20638 33182 20690 33234
rect 20750 33182 20802 33234
rect 21534 33182 21586 33234
rect 21646 33182 21698 33234
rect 25230 33182 25282 33234
rect 25566 33182 25618 33234
rect 29262 33182 29314 33234
rect 30046 33182 30098 33234
rect 31166 33182 31218 33234
rect 31838 33182 31890 33234
rect 32062 33182 32114 33234
rect 32286 33182 32338 33234
rect 32846 33182 32898 33234
rect 36430 33182 36482 33234
rect 37998 33182 38050 33234
rect 43038 33182 43090 33234
rect 51774 33182 51826 33234
rect 54462 33182 54514 33234
rect 57150 33182 57202 33234
rect 57262 33182 57314 33234
rect 59950 33182 60002 33234
rect 67006 33182 67058 33234
rect 67342 33182 67394 33234
rect 76302 33182 76354 33234
rect 14142 33070 14194 33122
rect 15822 33070 15874 33122
rect 16718 33070 16770 33122
rect 18510 33070 18562 33122
rect 20302 33070 20354 33122
rect 20414 33070 20466 33122
rect 21310 33070 21362 33122
rect 22878 33070 22930 33122
rect 23326 33070 23378 33122
rect 23774 33070 23826 33122
rect 24334 33070 24386 33122
rect 25790 33070 25842 33122
rect 26350 33070 26402 33122
rect 28590 33070 28642 33122
rect 29822 33070 29874 33122
rect 34750 33070 34802 33122
rect 37102 33070 37154 33122
rect 42702 33070 42754 33122
rect 43934 33070 43986 33122
rect 46286 33070 46338 33122
rect 48974 33070 49026 33122
rect 57598 33070 57650 33122
rect 65998 33070 66050 33122
rect 75406 33070 75458 33122
rect 20534 32902 20586 32954
rect 20638 32902 20690 32954
rect 20742 32902 20794 32954
rect 39854 32902 39906 32954
rect 39958 32902 40010 32954
rect 40062 32902 40114 32954
rect 59174 32902 59226 32954
rect 59278 32902 59330 32954
rect 59382 32902 59434 32954
rect 78494 32902 78546 32954
rect 78598 32902 78650 32954
rect 78702 32902 78754 32954
rect 14254 32734 14306 32786
rect 14366 32734 14418 32786
rect 16382 32734 16434 32786
rect 20974 32734 21026 32786
rect 22990 32734 23042 32786
rect 33294 32734 33346 32786
rect 36990 32734 37042 32786
rect 39006 32734 39058 32786
rect 39342 32734 39394 32786
rect 43038 32734 43090 32786
rect 44270 32734 44322 32786
rect 45614 32734 45666 32786
rect 46286 32734 46338 32786
rect 49870 32734 49922 32786
rect 57374 32734 57426 32786
rect 59838 32734 59890 32786
rect 67790 32734 67842 32786
rect 71598 32734 71650 32786
rect 72382 32734 72434 32786
rect 13918 32622 13970 32674
rect 15374 32622 15426 32674
rect 19518 32622 19570 32674
rect 23662 32622 23714 32674
rect 25230 32622 25282 32674
rect 28254 32622 28306 32674
rect 37214 32622 37266 32674
rect 38894 32622 38946 32674
rect 44830 32622 44882 32674
rect 45166 32622 45218 32674
rect 46622 32622 46674 32674
rect 50766 32622 50818 32674
rect 59950 32622 60002 32674
rect 66894 32622 66946 32674
rect 70702 32622 70754 32674
rect 14142 32510 14194 32562
rect 14590 32510 14642 32562
rect 14926 32510 14978 32562
rect 15150 32510 15202 32562
rect 15486 32510 15538 32562
rect 18958 32510 19010 32562
rect 19294 32510 19346 32562
rect 19966 32510 20018 32562
rect 25454 32510 25506 32562
rect 25790 32510 25842 32562
rect 26126 32510 26178 32562
rect 27358 32510 27410 32562
rect 28142 32510 28194 32562
rect 29934 32510 29986 32562
rect 30830 32510 30882 32562
rect 31838 32510 31890 32562
rect 36654 32510 36706 32562
rect 37438 32510 37490 32562
rect 37886 32510 37938 32562
rect 39678 32510 39730 32562
rect 39902 32510 39954 32562
rect 43374 32510 43426 32562
rect 43710 32510 43762 32562
rect 50654 32510 50706 32562
rect 50990 32510 51042 32562
rect 51550 32510 51602 32562
rect 58158 32510 58210 32562
rect 60734 32510 60786 32562
rect 66670 32510 66722 32562
rect 67454 32510 67506 32562
rect 70478 32510 70530 32562
rect 72718 32510 72770 32562
rect 75630 32510 75682 32562
rect 15934 32398 15986 32450
rect 19182 32398 19234 32450
rect 20414 32398 20466 32450
rect 22542 32398 22594 32450
rect 23662 32398 23714 32450
rect 25342 32398 25394 32450
rect 26574 32398 26626 32450
rect 27918 32398 27970 32450
rect 30718 32398 30770 32450
rect 33854 32398 33906 32450
rect 34302 32398 34354 32450
rect 35758 32398 35810 32450
rect 36318 32398 36370 32450
rect 37550 32398 37602 32450
rect 38446 32398 38498 32450
rect 42030 32398 42082 32450
rect 42702 32398 42754 32450
rect 50430 32398 50482 32450
rect 52334 32398 52386 32450
rect 54462 32398 54514 32450
rect 58494 32398 58546 32450
rect 59390 32398 59442 32450
rect 61518 32398 61570 32450
rect 63646 32398 63698 32450
rect 66222 32398 66274 32450
rect 69246 32398 69298 32450
rect 69806 32398 69858 32450
rect 75070 32398 75122 32450
rect 23886 32286 23938 32338
rect 36542 32286 36594 32338
rect 43934 32286 43986 32338
rect 59726 32286 59778 32338
rect 71262 32286 71314 32338
rect 77982 32286 78034 32338
rect 10874 32118 10926 32170
rect 10978 32118 11030 32170
rect 11082 32118 11134 32170
rect 30194 32118 30246 32170
rect 30298 32118 30350 32170
rect 30402 32118 30454 32170
rect 49514 32118 49566 32170
rect 49618 32118 49670 32170
rect 49722 32118 49774 32170
rect 68834 32118 68886 32170
rect 68938 32118 68990 32170
rect 69042 32118 69094 32170
rect 29822 31950 29874 32002
rect 37102 31950 37154 32002
rect 44830 31950 44882 32002
rect 60958 31950 61010 32002
rect 1934 31838 1986 31890
rect 15262 31838 15314 31890
rect 18398 31838 18450 31890
rect 20414 31838 20466 31890
rect 23326 31838 23378 31890
rect 25454 31838 25506 31890
rect 29486 31838 29538 31890
rect 31390 31838 31442 31890
rect 33182 31838 33234 31890
rect 37326 31838 37378 31890
rect 39230 31838 39282 31890
rect 46174 31838 46226 31890
rect 53454 31838 53506 31890
rect 59726 31838 59778 31890
rect 61630 31838 61682 31890
rect 73390 31838 73442 31890
rect 4286 31726 4338 31778
rect 18846 31726 18898 31778
rect 20302 31726 20354 31778
rect 22430 31726 22482 31778
rect 22766 31726 22818 31778
rect 23550 31726 23602 31778
rect 24222 31726 24274 31778
rect 24670 31726 24722 31778
rect 26238 31726 26290 31778
rect 26462 31726 26514 31778
rect 26686 31726 26738 31778
rect 30158 31726 30210 31778
rect 31278 31726 31330 31778
rect 31502 31726 31554 31778
rect 31838 31726 31890 31778
rect 32174 31726 32226 31778
rect 32398 31726 32450 31778
rect 33518 31726 33570 31778
rect 37550 31726 37602 31778
rect 38334 31726 38386 31778
rect 39006 31726 39058 31778
rect 41246 31726 41298 31778
rect 42590 31726 42642 31778
rect 43150 31726 43202 31778
rect 51662 31726 51714 31778
rect 53566 31726 53618 31778
rect 53902 31726 53954 31778
rect 70478 31726 70530 31778
rect 75406 31726 75458 31778
rect 8990 31614 9042 31666
rect 16158 31614 16210 31666
rect 17838 31614 17890 31666
rect 22878 31614 22930 31666
rect 25006 31614 25058 31666
rect 27358 31614 27410 31666
rect 30382 31614 30434 31666
rect 30942 31614 30994 31666
rect 32062 31614 32114 31666
rect 41022 31614 41074 31666
rect 42254 31614 42306 31666
rect 42366 31614 42418 31666
rect 42926 31614 42978 31666
rect 43486 31614 43538 31666
rect 44942 31614 44994 31666
rect 49646 31614 49698 31666
rect 49870 31614 49922 31666
rect 50206 31614 50258 31666
rect 50654 31614 50706 31666
rect 50766 31614 50818 31666
rect 51438 31614 51490 31666
rect 51998 31614 52050 31666
rect 53342 31614 53394 31666
rect 60622 31614 60674 31666
rect 60846 31614 60898 31666
rect 61294 31614 61346 31666
rect 61518 31614 61570 31666
rect 64878 31614 64930 31666
rect 65214 31614 65266 31666
rect 65886 31614 65938 31666
rect 69134 31614 69186 31666
rect 69806 31614 69858 31666
rect 71262 31614 71314 31666
rect 8654 31502 8706 31554
rect 9438 31502 9490 31554
rect 15934 31502 15986 31554
rect 16046 31502 16098 31554
rect 23886 31502 23938 31554
rect 27134 31502 27186 31554
rect 27694 31502 27746 31554
rect 32846 31502 32898 31554
rect 37438 31502 37490 31554
rect 38110 31502 38162 31554
rect 43150 31502 43202 31554
rect 43934 31502 43986 31554
rect 45390 31502 45442 31554
rect 46734 31502 46786 31554
rect 48638 31502 48690 31554
rect 48974 31502 49026 31554
rect 49982 31502 50034 31554
rect 50990 31502 51042 31554
rect 51886 31502 51938 31554
rect 58718 31502 58770 31554
rect 65550 31502 65602 31554
rect 66334 31502 66386 31554
rect 69470 31502 69522 31554
rect 70142 31502 70194 31554
rect 75630 31502 75682 31554
rect 20534 31334 20586 31386
rect 20638 31334 20690 31386
rect 20742 31334 20794 31386
rect 39854 31334 39906 31386
rect 39958 31334 40010 31386
rect 40062 31334 40114 31386
rect 59174 31334 59226 31386
rect 59278 31334 59330 31386
rect 59382 31334 59434 31386
rect 78494 31334 78546 31386
rect 78598 31334 78650 31386
rect 78702 31334 78754 31386
rect 17950 31166 18002 31218
rect 18510 31166 18562 31218
rect 20414 31166 20466 31218
rect 31502 31166 31554 31218
rect 33406 31166 33458 31218
rect 35646 31166 35698 31218
rect 36990 31166 37042 31218
rect 40014 31166 40066 31218
rect 40238 31166 40290 31218
rect 43710 31166 43762 31218
rect 49422 31166 49474 31218
rect 49646 31166 49698 31218
rect 51102 31166 51154 31218
rect 60062 31166 60114 31218
rect 71038 31166 71090 31218
rect 9550 31054 9602 31106
rect 16382 31054 16434 31106
rect 19630 31054 19682 31106
rect 19854 31054 19906 31106
rect 20078 31054 20130 31106
rect 20190 31054 20242 31106
rect 22878 31054 22930 31106
rect 24110 31054 24162 31106
rect 30158 31054 30210 31106
rect 30830 31054 30882 31106
rect 36094 31054 36146 31106
rect 39342 31054 39394 31106
rect 44606 31054 44658 31106
rect 48974 31054 49026 31106
rect 49310 31054 49362 31106
rect 51774 31054 51826 31106
rect 51998 31054 52050 31106
rect 65438 31054 65490 31106
rect 69806 31054 69858 31106
rect 74174 31054 74226 31106
rect 74510 31054 74562 31106
rect 9774 30942 9826 30994
rect 14478 30942 14530 30994
rect 14814 30942 14866 30994
rect 15486 30942 15538 30994
rect 15822 30942 15874 30994
rect 18398 30942 18450 30994
rect 18622 30942 18674 30994
rect 19518 30942 19570 30994
rect 21422 30942 21474 30994
rect 24670 30942 24722 30994
rect 25902 30942 25954 30994
rect 26238 30942 26290 30994
rect 28254 30942 28306 30994
rect 28590 30942 28642 30994
rect 29934 30942 29986 30994
rect 30494 30942 30546 30994
rect 31614 30942 31666 30994
rect 35982 30942 36034 30994
rect 37214 30942 37266 30994
rect 37438 30942 37490 30994
rect 37774 30942 37826 30994
rect 37998 30942 38050 30994
rect 38110 30942 38162 30994
rect 39454 30942 39506 30994
rect 39790 30942 39842 30994
rect 41022 30942 41074 30994
rect 42142 30942 42194 30994
rect 43598 30942 43650 30994
rect 43822 30942 43874 30994
rect 44270 30942 44322 30994
rect 47518 30942 47570 30994
rect 50990 30942 51042 30994
rect 51326 30942 51378 30994
rect 51550 30942 51602 30994
rect 52222 30942 52274 30994
rect 57822 30942 57874 30994
rect 59054 30942 59106 30994
rect 59390 30942 59442 30994
rect 59950 30942 60002 30994
rect 60398 30942 60450 30994
rect 64766 30942 64818 30994
rect 70142 30942 70194 30994
rect 71374 30942 71426 30994
rect 74846 30942 74898 30994
rect 14926 30830 14978 30882
rect 16270 30830 16322 30882
rect 16830 30830 16882 30882
rect 18062 30830 18114 30882
rect 20750 30830 20802 30882
rect 23438 30830 23490 30882
rect 25342 30830 25394 30882
rect 34638 30830 34690 30882
rect 36654 30830 36706 30882
rect 36990 30830 37042 30882
rect 41806 30830 41858 30882
rect 42590 30830 42642 30882
rect 43150 30830 43202 30882
rect 47966 30830 48018 30882
rect 50654 30830 50706 30882
rect 57598 30830 57650 30882
rect 58606 30830 58658 30882
rect 59726 30830 59778 30882
rect 67566 30830 67618 30882
rect 68126 30830 68178 30882
rect 72494 30830 72546 30882
rect 75630 30830 75682 30882
rect 77758 30830 77810 30882
rect 17726 30718 17778 30770
rect 38558 30718 38610 30770
rect 44382 30718 44434 30770
rect 44718 30718 44770 30770
rect 57374 30718 57426 30770
rect 58270 30718 58322 30770
rect 58494 30718 58546 30770
rect 59502 30718 59554 30770
rect 10874 30550 10926 30602
rect 10978 30550 11030 30602
rect 11082 30550 11134 30602
rect 30194 30550 30246 30602
rect 30298 30550 30350 30602
rect 30402 30550 30454 30602
rect 49514 30550 49566 30602
rect 49618 30550 49670 30602
rect 49722 30550 49774 30602
rect 68834 30550 68886 30602
rect 68938 30550 68990 30602
rect 69042 30550 69094 30602
rect 16494 30382 16546 30434
rect 17950 30382 18002 30434
rect 20078 30382 20130 30434
rect 26014 30382 26066 30434
rect 36094 30382 36146 30434
rect 36430 30382 36482 30434
rect 53790 30382 53842 30434
rect 9214 30270 9266 30322
rect 11342 30270 11394 30322
rect 19070 30270 19122 30322
rect 23326 30270 23378 30322
rect 24894 30270 24946 30322
rect 25790 30270 25842 30322
rect 28366 30270 28418 30322
rect 34526 30270 34578 30322
rect 35870 30270 35922 30322
rect 39454 30270 39506 30322
rect 41918 30270 41970 30322
rect 43710 30270 43762 30322
rect 46846 30270 46898 30322
rect 61294 30270 61346 30322
rect 69806 30270 69858 30322
rect 73390 30270 73442 30322
rect 74734 30270 74786 30322
rect 76638 30270 76690 30322
rect 8542 30158 8594 30210
rect 14366 30158 14418 30210
rect 14702 30158 14754 30210
rect 15598 30158 15650 30210
rect 17278 30158 17330 30210
rect 17838 30158 17890 30210
rect 18622 30158 18674 30210
rect 19518 30158 19570 30210
rect 21758 30158 21810 30210
rect 22094 30158 22146 30210
rect 23774 30158 23826 30210
rect 23998 30158 24050 30210
rect 24782 30158 24834 30210
rect 25678 30158 25730 30210
rect 28254 30158 28306 30210
rect 29598 30158 29650 30210
rect 31726 30158 31778 30210
rect 34078 30158 34130 30210
rect 34302 30158 34354 30210
rect 34862 30158 34914 30210
rect 37662 30158 37714 30210
rect 38110 30158 38162 30210
rect 38670 30158 38722 30210
rect 39118 30158 39170 30210
rect 41470 30158 41522 30210
rect 42590 30158 42642 30210
rect 48078 30158 48130 30210
rect 53566 30158 53618 30210
rect 56702 30158 56754 30210
rect 58158 30158 58210 30210
rect 58942 30158 58994 30210
rect 59502 30158 59554 30210
rect 60510 30158 60562 30210
rect 60958 30158 61010 30210
rect 61182 30158 61234 30210
rect 64654 30158 64706 30210
rect 68574 30158 68626 30210
rect 69134 30158 69186 30210
rect 72830 30158 72882 30210
rect 73726 30158 73778 30210
rect 75518 30158 75570 30210
rect 77982 30158 78034 30210
rect 3726 30046 3778 30098
rect 15262 30046 15314 30098
rect 15934 30046 15986 30098
rect 16382 30046 16434 30098
rect 20526 30046 20578 30098
rect 28366 30046 28418 30098
rect 29710 30046 29762 30098
rect 33294 30046 33346 30098
rect 37326 30046 37378 30098
rect 43598 30046 43650 30098
rect 43822 30046 43874 30098
rect 47406 30046 47458 30098
rect 57822 30046 57874 30098
rect 58830 30046 58882 30098
rect 60734 30046 60786 30098
rect 61406 30046 61458 30098
rect 61742 30046 61794 30098
rect 65326 30046 65378 30098
rect 72718 30046 72770 30098
rect 75294 30046 75346 30098
rect 76302 30046 76354 30098
rect 76974 30046 77026 30098
rect 77422 30046 77474 30098
rect 3390 29934 3442 29986
rect 5854 29934 5906 29986
rect 15822 29934 15874 29986
rect 26686 29934 26738 29986
rect 29262 29934 29314 29986
rect 31166 29934 31218 29986
rect 33854 29934 33906 29986
rect 33966 29934 34018 29986
rect 35198 29934 35250 29986
rect 38110 29934 38162 29986
rect 43150 29934 43202 29986
rect 44046 29934 44098 29986
rect 44942 29934 44994 29986
rect 45278 29934 45330 29986
rect 45726 29934 45778 29986
rect 46846 29934 46898 29986
rect 46958 29934 47010 29986
rect 47182 29934 47234 29986
rect 47742 29934 47794 29986
rect 54126 29934 54178 29986
rect 57150 29934 57202 29986
rect 60062 29934 60114 29986
rect 62078 29934 62130 29986
rect 67566 29934 67618 29986
rect 68350 29934 68402 29986
rect 72046 29934 72098 29986
rect 74398 29934 74450 29986
rect 20534 29766 20586 29818
rect 20638 29766 20690 29818
rect 20742 29766 20794 29818
rect 39854 29766 39906 29818
rect 39958 29766 40010 29818
rect 40062 29766 40114 29818
rect 59174 29766 59226 29818
rect 59278 29766 59330 29818
rect 59382 29766 59434 29818
rect 78494 29766 78546 29818
rect 78598 29766 78650 29818
rect 78702 29766 78754 29818
rect 5742 29598 5794 29650
rect 9662 29598 9714 29650
rect 16270 29598 16322 29650
rect 17390 29598 17442 29650
rect 17502 29598 17554 29650
rect 19182 29598 19234 29650
rect 20750 29598 20802 29650
rect 22766 29598 22818 29650
rect 29934 29598 29986 29650
rect 30158 29598 30210 29650
rect 32286 29598 32338 29650
rect 35646 29598 35698 29650
rect 38222 29598 38274 29650
rect 39006 29598 39058 29650
rect 40014 29598 40066 29650
rect 42030 29598 42082 29650
rect 42478 29598 42530 29650
rect 43038 29598 43090 29650
rect 47742 29598 47794 29650
rect 49086 29598 49138 29650
rect 49198 29598 49250 29650
rect 51774 29598 51826 29650
rect 51886 29598 51938 29650
rect 53454 29598 53506 29650
rect 54686 29598 54738 29650
rect 59726 29598 59778 29650
rect 60398 29598 60450 29650
rect 62638 29598 62690 29650
rect 65102 29598 65154 29650
rect 65438 29598 65490 29650
rect 70142 29598 70194 29650
rect 74510 29598 74562 29650
rect 3166 29486 3218 29538
rect 6750 29486 6802 29538
rect 7982 29486 8034 29538
rect 10222 29486 10274 29538
rect 10558 29486 10610 29538
rect 13134 29486 13186 29538
rect 13246 29486 13298 29538
rect 15150 29486 15202 29538
rect 17838 29486 17890 29538
rect 20302 29486 20354 29538
rect 20414 29486 20466 29538
rect 20638 29486 20690 29538
rect 20974 29486 21026 29538
rect 22094 29486 22146 29538
rect 24222 29486 24274 29538
rect 26126 29486 26178 29538
rect 26462 29486 26514 29538
rect 27134 29486 27186 29538
rect 32062 29486 32114 29538
rect 33182 29486 33234 29538
rect 35422 29486 35474 29538
rect 35534 29486 35586 29538
rect 36430 29486 36482 29538
rect 38446 29486 38498 29538
rect 40238 29486 40290 29538
rect 43934 29486 43986 29538
rect 46174 29486 46226 29538
rect 47854 29486 47906 29538
rect 49646 29486 49698 29538
rect 49758 29486 49810 29538
rect 55358 29486 55410 29538
rect 60846 29486 60898 29538
rect 64766 29486 64818 29538
rect 66894 29486 66946 29538
rect 67230 29486 67282 29538
rect 70702 29486 70754 29538
rect 71038 29486 71090 29538
rect 72270 29486 72322 29538
rect 75630 29486 75682 29538
rect 2494 29374 2546 29426
rect 6526 29374 6578 29426
rect 8318 29374 8370 29426
rect 9998 29374 10050 29426
rect 13694 29374 13746 29426
rect 14254 29374 14306 29426
rect 14926 29374 14978 29426
rect 15598 29374 15650 29426
rect 16494 29374 16546 29426
rect 16718 29374 16770 29426
rect 17614 29374 17666 29426
rect 19070 29374 19122 29426
rect 19294 29374 19346 29426
rect 21086 29374 21138 29426
rect 22430 29374 22482 29426
rect 23438 29374 23490 29426
rect 25566 29374 25618 29426
rect 26574 29374 26626 29426
rect 27582 29374 27634 29426
rect 29598 29374 29650 29426
rect 30830 29374 30882 29426
rect 31054 29374 31106 29426
rect 33070 29374 33122 29426
rect 33966 29374 34018 29426
rect 35870 29374 35922 29426
rect 36206 29374 36258 29426
rect 36878 29374 36930 29426
rect 37662 29374 37714 29426
rect 38558 29374 38610 29426
rect 38894 29374 38946 29426
rect 40126 29374 40178 29426
rect 42366 29374 42418 29426
rect 42702 29374 42754 29426
rect 43374 29374 43426 29426
rect 44158 29374 44210 29426
rect 44718 29374 44770 29426
rect 48638 29374 48690 29426
rect 49310 29374 49362 29426
rect 51662 29374 51714 29426
rect 51998 29374 52050 29426
rect 52222 29374 52274 29426
rect 53118 29374 53170 29426
rect 53678 29374 53730 29426
rect 54126 29374 54178 29426
rect 54238 29374 54290 29426
rect 54910 29374 54962 29426
rect 55582 29374 55634 29426
rect 58046 29374 58098 29426
rect 58270 29374 58322 29426
rect 59390 29374 59442 29426
rect 59950 29374 60002 29426
rect 60958 29374 61010 29426
rect 61182 29374 61234 29426
rect 62190 29374 62242 29426
rect 62414 29374 62466 29426
rect 62750 29374 62802 29426
rect 62974 29374 63026 29426
rect 65774 29374 65826 29426
rect 66222 29374 66274 29426
rect 72494 29374 72546 29426
rect 74286 29374 74338 29426
rect 74846 29374 74898 29426
rect 5294 29262 5346 29314
rect 7422 29262 7474 29314
rect 11342 29262 11394 29314
rect 11790 29262 11842 29314
rect 15374 29262 15426 29314
rect 16606 29262 16658 29314
rect 19742 29262 19794 29314
rect 28030 29262 28082 29314
rect 28590 29262 28642 29314
rect 30046 29262 30098 29314
rect 31502 29262 31554 29314
rect 33182 29262 33234 29314
rect 35758 29262 35810 29314
rect 41246 29262 41298 29314
rect 41694 29262 41746 29314
rect 45950 29262 46002 29314
rect 52894 29262 52946 29314
rect 53902 29262 53954 29314
rect 67902 29262 67954 29314
rect 69694 29262 69746 29314
rect 73838 29262 73890 29314
rect 77758 29262 77810 29314
rect 6078 29150 6130 29202
rect 13246 29150 13298 29202
rect 31614 29150 31666 29202
rect 32398 29150 32450 29202
rect 36542 29150 36594 29202
rect 49758 29150 49810 29202
rect 58270 29150 58322 29202
rect 59614 29150 59666 29202
rect 66558 29150 66610 29202
rect 70478 29150 70530 29202
rect 10874 28982 10926 29034
rect 10978 28982 11030 29034
rect 11082 28982 11134 29034
rect 30194 28982 30246 29034
rect 30298 28982 30350 29034
rect 30402 28982 30454 29034
rect 49514 28982 49566 29034
rect 49618 28982 49670 29034
rect 49722 28982 49774 29034
rect 68834 28982 68886 29034
rect 68938 28982 68990 29034
rect 69042 28982 69094 29034
rect 13694 28814 13746 28866
rect 21982 28814 22034 28866
rect 24670 28814 24722 28866
rect 25454 28814 25506 28866
rect 25790 28814 25842 28866
rect 35198 28814 35250 28866
rect 40350 28814 40402 28866
rect 40686 28814 40738 28866
rect 48302 28814 48354 28866
rect 54574 28814 54626 28866
rect 57486 28814 57538 28866
rect 59614 28814 59666 28866
rect 59950 28814 60002 28866
rect 66334 28814 66386 28866
rect 66670 28814 66722 28866
rect 5070 28702 5122 28754
rect 7870 28702 7922 28754
rect 9998 28702 10050 28754
rect 13806 28702 13858 28754
rect 14702 28702 14754 28754
rect 20190 28702 20242 28754
rect 20750 28702 20802 28754
rect 30270 28702 30322 28754
rect 31278 28702 31330 28754
rect 37662 28702 37714 28754
rect 38558 28702 38610 28754
rect 40910 28702 40962 28754
rect 41582 28702 41634 28754
rect 42366 28702 42418 28754
rect 42814 28702 42866 28754
rect 46062 28702 46114 28754
rect 49982 28702 50034 28754
rect 53006 28702 53058 28754
rect 54798 28702 54850 28754
rect 58046 28702 58098 28754
rect 58942 28702 58994 28754
rect 61518 28702 61570 28754
rect 72718 28702 72770 28754
rect 75406 28702 75458 28754
rect 2270 28590 2322 28642
rect 2942 28590 2994 28642
rect 5854 28590 5906 28642
rect 7086 28590 7138 28642
rect 14254 28590 14306 28642
rect 16158 28590 16210 28642
rect 17054 28590 17106 28642
rect 18286 28590 18338 28642
rect 19070 28590 19122 28642
rect 19630 28590 19682 28642
rect 21310 28590 21362 28642
rect 21646 28590 21698 28642
rect 23886 28590 23938 28642
rect 24894 28590 24946 28642
rect 25790 28590 25842 28642
rect 26238 28590 26290 28642
rect 27918 28590 27970 28642
rect 29822 28590 29874 28642
rect 30046 28590 30098 28642
rect 31166 28590 31218 28642
rect 32398 28590 32450 28642
rect 33966 28590 34018 28642
rect 34526 28590 34578 28642
rect 35310 28590 35362 28642
rect 35870 28590 35922 28642
rect 36094 28590 36146 28642
rect 36990 28590 37042 28642
rect 39342 28590 39394 28642
rect 39790 28590 39842 28642
rect 41694 28590 41746 28642
rect 46622 28590 46674 28642
rect 47294 28590 47346 28642
rect 47854 28590 47906 28642
rect 51438 28590 51490 28642
rect 52670 28590 52722 28642
rect 53230 28590 53282 28642
rect 54014 28590 54066 28642
rect 54350 28590 54402 28642
rect 55918 28590 55970 28642
rect 57934 28590 57986 28642
rect 58270 28590 58322 28642
rect 58494 28590 58546 28642
rect 58718 28590 58770 28642
rect 59950 28590 60002 28642
rect 61630 28590 61682 28642
rect 62078 28590 62130 28642
rect 62302 28590 62354 28642
rect 65886 28590 65938 28642
rect 67118 28590 67170 28642
rect 71934 28590 71986 28642
rect 73054 28590 73106 28642
rect 5630 28478 5682 28530
rect 15710 28478 15762 28530
rect 26462 28478 26514 28530
rect 26574 28478 26626 28530
rect 27134 28478 27186 28530
rect 28142 28478 28194 28530
rect 30942 28478 30994 28530
rect 34862 28478 34914 28530
rect 36430 28478 36482 28530
rect 38670 28478 38722 28530
rect 39006 28478 39058 28530
rect 41582 28478 41634 28530
rect 46398 28478 46450 28530
rect 48190 28478 48242 28530
rect 48302 28478 48354 28530
rect 50318 28478 50370 28530
rect 53790 28478 53842 28530
rect 54910 28478 54962 28530
rect 55022 28478 55074 28530
rect 55694 28478 55746 28530
rect 57598 28478 57650 28530
rect 59054 28478 59106 28530
rect 59278 28478 59330 28530
rect 62638 28478 62690 28530
rect 67230 28478 67282 28530
rect 11230 28366 11282 28418
rect 17166 28366 17218 28418
rect 24334 28366 24386 28418
rect 24558 28366 24610 28418
rect 26798 28366 26850 28418
rect 27022 28366 27074 28418
rect 34750 28366 34802 28418
rect 36318 28366 36370 28418
rect 39566 28366 39618 28418
rect 39902 28366 39954 28418
rect 40126 28366 40178 28418
rect 46062 28366 46114 28418
rect 46174 28366 46226 28418
rect 51998 28366 52050 28418
rect 52894 28366 52946 28418
rect 53118 28366 53170 28418
rect 56254 28366 56306 28418
rect 56702 28366 56754 28418
rect 57038 28366 57090 28418
rect 57486 28366 57538 28418
rect 60734 28366 60786 28418
rect 62526 28366 62578 28418
rect 76302 28366 76354 28418
rect 20534 28198 20586 28250
rect 20638 28198 20690 28250
rect 20742 28198 20794 28250
rect 39854 28198 39906 28250
rect 39958 28198 40010 28250
rect 40062 28198 40114 28250
rect 59174 28198 59226 28250
rect 59278 28198 59330 28250
rect 59382 28198 59434 28250
rect 78494 28198 78546 28250
rect 78598 28198 78650 28250
rect 78702 28198 78754 28250
rect 5854 28030 5906 28082
rect 9662 28030 9714 28082
rect 15038 28030 15090 28082
rect 17726 28030 17778 28082
rect 19294 28030 19346 28082
rect 19854 28030 19906 28082
rect 21758 28030 21810 28082
rect 23326 28030 23378 28082
rect 24558 28030 24610 28082
rect 25454 28030 25506 28082
rect 27806 28030 27858 28082
rect 28030 28030 28082 28082
rect 28702 28030 28754 28082
rect 33294 28030 33346 28082
rect 34414 28030 34466 28082
rect 34638 28030 34690 28082
rect 35422 28030 35474 28082
rect 38782 28030 38834 28082
rect 41134 28030 41186 28082
rect 43262 28030 43314 28082
rect 43934 28030 43986 28082
rect 44158 28030 44210 28082
rect 44382 28030 44434 28082
rect 48862 28030 48914 28082
rect 49758 28030 49810 28082
rect 49982 28030 50034 28082
rect 50318 28030 50370 28082
rect 51438 28030 51490 28082
rect 54574 28030 54626 28082
rect 60510 28030 60562 28082
rect 61294 28030 61346 28082
rect 61406 28030 61458 28082
rect 72382 28030 72434 28082
rect 72606 28030 72658 28082
rect 74174 28030 74226 28082
rect 4958 27918 5010 27970
rect 5294 27918 5346 27970
rect 10222 27918 10274 27970
rect 10558 27918 10610 27970
rect 11342 27918 11394 27970
rect 18734 27918 18786 27970
rect 20078 27918 20130 27970
rect 21870 27918 21922 27970
rect 22878 27918 22930 27970
rect 23102 27918 23154 27970
rect 24446 27918 24498 27970
rect 25902 27918 25954 27970
rect 32286 27918 32338 27970
rect 33630 27918 33682 27970
rect 34862 27918 34914 27970
rect 38446 27918 38498 27970
rect 39790 27918 39842 27970
rect 40238 27918 40290 27970
rect 41358 27918 41410 27970
rect 42702 27918 42754 27970
rect 42814 27918 42866 27970
rect 48078 27918 48130 27970
rect 49198 27918 49250 27970
rect 50654 27918 50706 27970
rect 59614 27918 59666 27970
rect 70142 27918 70194 27970
rect 71374 27918 71426 27970
rect 73278 27918 73330 27970
rect 75070 27918 75122 27970
rect 4286 27806 4338 27858
rect 11678 27806 11730 27858
rect 15374 27806 15426 27858
rect 17838 27806 17890 27858
rect 18174 27806 18226 27858
rect 19630 27806 19682 27858
rect 20190 27806 20242 27858
rect 20750 27806 20802 27858
rect 23438 27806 23490 27858
rect 25230 27806 25282 27858
rect 26350 27806 26402 27858
rect 28142 27806 28194 27858
rect 29038 27806 29090 27858
rect 30382 27806 30434 27858
rect 30494 27806 30546 27858
rect 30718 27806 30770 27858
rect 31502 27806 31554 27858
rect 32174 27806 32226 27858
rect 33742 27806 33794 27858
rect 34190 27806 34242 27858
rect 34974 27806 35026 27858
rect 37998 27806 38050 27858
rect 38334 27806 38386 27858
rect 41470 27806 41522 27858
rect 42478 27806 42530 27858
rect 44494 27806 44546 27858
rect 46958 27806 47010 27858
rect 47742 27806 47794 27858
rect 50878 27806 50930 27858
rect 52110 27806 52162 27858
rect 53678 27806 53730 27858
rect 54910 27806 54962 27858
rect 58718 27806 58770 27858
rect 59054 27806 59106 27858
rect 60174 27806 60226 27858
rect 60734 27806 60786 27858
rect 61182 27806 61234 27858
rect 62078 27806 62130 27858
rect 62526 27806 62578 27858
rect 63422 27806 63474 27858
rect 68574 27806 68626 27858
rect 68686 27806 68738 27858
rect 68910 27806 68962 27858
rect 69134 27806 69186 27858
rect 70366 27806 70418 27858
rect 70702 27806 70754 27858
rect 70926 27806 70978 27858
rect 71150 27806 71202 27858
rect 71262 27806 71314 27858
rect 71598 27806 71650 27858
rect 72830 27806 72882 27858
rect 73166 27806 73218 27858
rect 74734 27806 74786 27858
rect 75630 27806 75682 27858
rect 1934 27694 1986 27746
rect 6414 27694 6466 27746
rect 6862 27694 6914 27746
rect 12126 27694 12178 27746
rect 15598 27694 15650 27746
rect 16270 27694 16322 27746
rect 16830 27694 16882 27746
rect 20526 27694 20578 27746
rect 21086 27694 21138 27746
rect 23998 27694 24050 27746
rect 26798 27694 26850 27746
rect 27358 27694 27410 27746
rect 31726 27694 31778 27746
rect 37102 27694 37154 27746
rect 39342 27694 39394 27746
rect 45054 27694 45106 27746
rect 45390 27694 45442 27746
rect 51886 27694 51938 27746
rect 55022 27694 55074 27746
rect 55246 27694 55298 27746
rect 56702 27694 56754 27746
rect 59278 27694 59330 27746
rect 68798 27694 68850 27746
rect 5518 27582 5570 27634
rect 9998 27582 10050 27634
rect 16494 27582 16546 27634
rect 24670 27582 24722 27634
rect 30830 27582 30882 27634
rect 39118 27582 39170 27634
rect 39678 27582 39730 27634
rect 40126 27582 40178 27634
rect 47294 27582 47346 27634
rect 53566 27582 53618 27634
rect 62302 27582 62354 27634
rect 70030 27582 70082 27634
rect 77982 27582 78034 27634
rect 10874 27414 10926 27466
rect 10978 27414 11030 27466
rect 11082 27414 11134 27466
rect 30194 27414 30246 27466
rect 30298 27414 30350 27466
rect 30402 27414 30454 27466
rect 49514 27414 49566 27466
rect 49618 27414 49670 27466
rect 49722 27414 49774 27466
rect 68834 27414 68886 27466
rect 68938 27414 68990 27466
rect 69042 27414 69094 27466
rect 18286 27246 18338 27298
rect 24782 27246 24834 27298
rect 30382 27246 30434 27298
rect 39006 27246 39058 27298
rect 42366 27246 42418 27298
rect 53454 27246 53506 27298
rect 58830 27246 58882 27298
rect 66222 27246 66274 27298
rect 73726 27246 73778 27298
rect 74398 27246 74450 27298
rect 4510 27134 4562 27186
rect 9550 27134 9602 27186
rect 10782 27134 10834 27186
rect 12910 27134 12962 27186
rect 18510 27134 18562 27186
rect 19070 27134 19122 27186
rect 25118 27134 25170 27186
rect 28366 27134 28418 27186
rect 37550 27134 37602 27186
rect 38222 27134 38274 27186
rect 44942 27134 44994 27186
rect 53566 27134 53618 27186
rect 58942 27134 58994 27186
rect 59390 27134 59442 27186
rect 60622 27134 60674 27186
rect 62078 27134 62130 27186
rect 69358 27134 69410 27186
rect 6750 27022 6802 27074
rect 10110 27022 10162 27074
rect 17390 27022 17442 27074
rect 18622 27022 18674 27074
rect 25790 27022 25842 27074
rect 26350 27022 26402 27074
rect 26686 27022 26738 27074
rect 27022 27022 27074 27074
rect 27582 27022 27634 27074
rect 30830 27022 30882 27074
rect 31726 27022 31778 27074
rect 32510 27022 32562 27074
rect 33966 27022 34018 27074
rect 36094 27022 36146 27074
rect 37886 27022 37938 27074
rect 38558 27022 38610 27074
rect 38782 27022 38834 27074
rect 39342 27022 39394 27074
rect 40238 27022 40290 27074
rect 42702 27022 42754 27074
rect 43486 27022 43538 27074
rect 44270 27022 44322 27074
rect 53454 27022 53506 27074
rect 54350 27022 54402 27074
rect 59278 27022 59330 27074
rect 59726 27022 59778 27074
rect 61630 27022 61682 27074
rect 62750 27022 62802 27074
rect 66334 27022 66386 27074
rect 67006 27022 67058 27074
rect 67566 27022 67618 27074
rect 69246 27022 69298 27074
rect 70366 27022 70418 27074
rect 72158 27022 72210 27074
rect 73726 27022 73778 27074
rect 74734 27022 74786 27074
rect 75518 27022 75570 27074
rect 76414 27022 76466 27074
rect 3166 26910 3218 26962
rect 7422 26910 7474 26962
rect 16494 26910 16546 26962
rect 16830 26910 16882 26962
rect 17166 26910 17218 26962
rect 21534 26910 21586 26962
rect 21646 26910 21698 26962
rect 21758 26910 21810 26962
rect 21870 26910 21922 26962
rect 22094 26910 22146 26962
rect 22206 26910 22258 26962
rect 22654 26910 22706 26962
rect 24558 26910 24610 26962
rect 26462 26910 26514 26962
rect 30382 26910 30434 26962
rect 30494 26910 30546 26962
rect 31278 26910 31330 26962
rect 32286 26910 32338 26962
rect 35534 26910 35586 26962
rect 39678 26910 39730 26962
rect 39902 26910 39954 26962
rect 41358 26910 41410 26962
rect 41694 26910 41746 26962
rect 43374 26910 43426 26962
rect 43934 26910 43986 26962
rect 44830 26910 44882 26962
rect 45502 26910 45554 26962
rect 45838 26910 45890 26962
rect 59614 26910 59666 26962
rect 61294 26910 61346 26962
rect 66558 26910 66610 26962
rect 70030 26910 70082 26962
rect 73166 26910 73218 26962
rect 75294 26910 75346 26962
rect 2830 26798 2882 26850
rect 17726 26798 17778 26850
rect 22766 26798 22818 26850
rect 22990 26798 23042 26850
rect 26910 26798 26962 26850
rect 31838 26798 31890 26850
rect 32734 26798 32786 26850
rect 38110 26798 38162 26850
rect 39342 26798 39394 26850
rect 39790 26798 39842 26850
rect 40798 26798 40850 26850
rect 45054 26798 45106 26850
rect 48414 26798 48466 26850
rect 50430 26798 50482 26850
rect 76190 26798 76242 26850
rect 20534 26630 20586 26682
rect 20638 26630 20690 26682
rect 20742 26630 20794 26682
rect 39854 26630 39906 26682
rect 39958 26630 40010 26682
rect 40062 26630 40114 26682
rect 59174 26630 59226 26682
rect 59278 26630 59330 26682
rect 59382 26630 59434 26682
rect 78494 26630 78546 26682
rect 78598 26630 78650 26682
rect 78702 26630 78754 26682
rect 7310 26462 7362 26514
rect 11006 26462 11058 26514
rect 11342 26462 11394 26514
rect 11790 26462 11842 26514
rect 22094 26462 22146 26514
rect 23662 26462 23714 26514
rect 25902 26462 25954 26514
rect 32398 26462 32450 26514
rect 36654 26462 36706 26514
rect 38782 26462 38834 26514
rect 42702 26462 42754 26514
rect 44606 26462 44658 26514
rect 46286 26462 46338 26514
rect 50542 26462 50594 26514
rect 50766 26462 50818 26514
rect 52782 26462 52834 26514
rect 54126 26462 54178 26514
rect 57038 26462 57090 26514
rect 58606 26462 58658 26514
rect 59614 26462 59666 26514
rect 59950 26462 60002 26514
rect 61630 26462 61682 26514
rect 63086 26462 63138 26514
rect 65326 26462 65378 26514
rect 66110 26462 66162 26514
rect 70030 26462 70082 26514
rect 73166 26462 73218 26514
rect 2494 26350 2546 26402
rect 8430 26350 8482 26402
rect 8878 26350 8930 26402
rect 16494 26350 16546 26402
rect 20638 26350 20690 26402
rect 26126 26350 26178 26402
rect 26238 26350 26290 26402
rect 31166 26350 31218 26402
rect 32174 26350 32226 26402
rect 33742 26350 33794 26402
rect 36766 26350 36818 26402
rect 37886 26350 37938 26402
rect 45166 26350 45218 26402
rect 48974 26350 49026 26402
rect 51102 26350 51154 26402
rect 57262 26350 57314 26402
rect 58942 26350 58994 26402
rect 59166 26350 59218 26402
rect 59502 26350 59554 26402
rect 61966 26350 62018 26402
rect 63310 26350 63362 26402
rect 63422 26350 63474 26402
rect 65438 26350 65490 26402
rect 71038 26350 71090 26402
rect 72494 26350 72546 26402
rect 73614 26350 73666 26402
rect 74958 26350 75010 26402
rect 1822 26238 1874 26290
rect 7086 26238 7138 26290
rect 7758 26238 7810 26290
rect 8094 26238 8146 26290
rect 14926 26238 14978 26290
rect 16830 26238 16882 26290
rect 18062 26238 18114 26290
rect 19406 26238 19458 26290
rect 19854 26238 19906 26290
rect 21198 26238 21250 26290
rect 21758 26238 21810 26290
rect 24334 26238 24386 26290
rect 27134 26238 27186 26290
rect 27470 26238 27522 26290
rect 28926 26238 28978 26290
rect 29374 26238 29426 26290
rect 31054 26238 31106 26290
rect 33070 26238 33122 26290
rect 35310 26238 35362 26290
rect 37998 26238 38050 26290
rect 38446 26238 38498 26290
rect 38670 26238 38722 26290
rect 40126 26238 40178 26290
rect 42478 26238 42530 26290
rect 42702 26238 42754 26290
rect 43038 26238 43090 26290
rect 45054 26238 45106 26290
rect 45278 26238 45330 26290
rect 46062 26238 46114 26290
rect 49086 26238 49138 26290
rect 50206 26238 50258 26290
rect 50654 26238 50706 26290
rect 50878 26238 50930 26290
rect 52558 26238 52610 26290
rect 52670 26238 52722 26290
rect 52894 26238 52946 26290
rect 53118 26238 53170 26290
rect 57374 26238 57426 26290
rect 59726 26238 59778 26290
rect 64878 26238 64930 26290
rect 65214 26238 65266 26290
rect 65886 26238 65938 26290
rect 65998 26238 66050 26290
rect 66222 26238 66274 26290
rect 66446 26238 66498 26290
rect 66782 26238 66834 26290
rect 68126 26238 68178 26290
rect 68574 26238 68626 26290
rect 69582 26238 69634 26290
rect 71486 26238 71538 26290
rect 72830 26238 72882 26290
rect 73166 26238 73218 26290
rect 74286 26238 74338 26290
rect 4622 26126 4674 26178
rect 9662 26126 9714 26178
rect 16046 26126 16098 26178
rect 16606 26126 16658 26178
rect 18398 26126 18450 26178
rect 18734 26126 18786 26178
rect 19182 26126 19234 26178
rect 20974 26126 21026 26178
rect 22654 26126 22706 26178
rect 25678 26126 25730 26178
rect 26686 26126 26738 26178
rect 28030 26126 28082 26178
rect 28590 26126 28642 26178
rect 29822 26126 29874 26178
rect 30718 26126 30770 26178
rect 31278 26126 31330 26178
rect 32510 26126 32562 26178
rect 37438 26126 37490 26178
rect 37550 26126 37602 26178
rect 39678 26126 39730 26178
rect 43486 26126 43538 26178
rect 48190 26126 48242 26178
rect 49534 26126 49586 26178
rect 64542 26126 64594 26178
rect 77086 26126 77138 26178
rect 19070 26014 19122 26066
rect 22430 26014 22482 26066
rect 45726 26014 45778 26066
rect 46398 26014 46450 26066
rect 58830 26014 58882 26066
rect 10874 25846 10926 25898
rect 10978 25846 11030 25898
rect 11082 25846 11134 25898
rect 30194 25846 30246 25898
rect 30298 25846 30350 25898
rect 30402 25846 30454 25898
rect 49514 25846 49566 25898
rect 49618 25846 49670 25898
rect 49722 25846 49774 25898
rect 68834 25846 68886 25898
rect 68938 25846 68990 25898
rect 69042 25846 69094 25898
rect 1934 25678 1986 25730
rect 11678 25678 11730 25730
rect 12014 25678 12066 25730
rect 27806 25678 27858 25730
rect 33966 25678 34018 25730
rect 50094 25678 50146 25730
rect 76302 25678 76354 25730
rect 76638 25678 76690 25730
rect 15486 25566 15538 25618
rect 18510 25566 18562 25618
rect 19854 25566 19906 25618
rect 24110 25566 24162 25618
rect 27918 25566 27970 25618
rect 30270 25566 30322 25618
rect 35198 25566 35250 25618
rect 35758 25566 35810 25618
rect 39006 25566 39058 25618
rect 40238 25566 40290 25618
rect 43822 25566 43874 25618
rect 44270 25566 44322 25618
rect 46398 25566 46450 25618
rect 47294 25566 47346 25618
rect 48750 25566 48802 25618
rect 49758 25566 49810 25618
rect 55582 25566 55634 25618
rect 58942 25566 58994 25618
rect 66222 25566 66274 25618
rect 67454 25566 67506 25618
rect 69694 25566 69746 25618
rect 73726 25566 73778 25618
rect 77982 25566 78034 25618
rect 4286 25454 4338 25506
rect 11118 25454 11170 25506
rect 12798 25454 12850 25506
rect 14926 25454 14978 25506
rect 16046 25454 16098 25506
rect 16718 25454 16770 25506
rect 17950 25454 18002 25506
rect 20078 25454 20130 25506
rect 20750 25454 20802 25506
rect 21646 25454 21698 25506
rect 23550 25454 23602 25506
rect 24222 25454 24274 25506
rect 25006 25454 25058 25506
rect 26350 25454 26402 25506
rect 27470 25454 27522 25506
rect 28142 25454 28194 25506
rect 33406 25454 33458 25506
rect 33630 25454 33682 25506
rect 34862 25454 34914 25506
rect 38446 25454 38498 25506
rect 40126 25454 40178 25506
rect 40350 25454 40402 25506
rect 44830 25454 44882 25506
rect 45166 25454 45218 25506
rect 45390 25454 45442 25506
rect 46846 25454 46898 25506
rect 48078 25454 48130 25506
rect 48302 25454 48354 25506
rect 49422 25454 49474 25506
rect 50430 25454 50482 25506
rect 53230 25454 53282 25506
rect 53678 25454 53730 25506
rect 54574 25454 54626 25506
rect 56254 25454 56306 25506
rect 56926 25454 56978 25506
rect 59614 25454 59666 25506
rect 59838 25454 59890 25506
rect 63422 25454 63474 25506
rect 67118 25454 67170 25506
rect 67342 25454 67394 25506
rect 68350 25454 68402 25506
rect 69246 25454 69298 25506
rect 71598 25454 71650 25506
rect 71934 25454 71986 25506
rect 72270 25454 72322 25506
rect 73502 25454 73554 25506
rect 75182 25454 75234 25506
rect 12574 25342 12626 25394
rect 13694 25342 13746 25394
rect 22318 25342 22370 25394
rect 26014 25342 26066 25394
rect 26910 25342 26962 25394
rect 27134 25342 27186 25394
rect 29262 25342 29314 25394
rect 29374 25342 29426 25394
rect 38894 25342 38946 25394
rect 39118 25342 39170 25394
rect 39678 25342 39730 25394
rect 47742 25342 47794 25394
rect 47854 25342 47906 25394
rect 48638 25342 48690 25394
rect 50766 25342 50818 25394
rect 54126 25342 54178 25394
rect 54798 25342 54850 25394
rect 57150 25342 57202 25394
rect 64094 25342 64146 25394
rect 67790 25342 67842 25394
rect 69358 25342 69410 25394
rect 73950 25342 74002 25394
rect 76862 25342 76914 25394
rect 77422 25342 77474 25394
rect 4846 25230 4898 25282
rect 10222 25230 10274 25282
rect 10782 25230 10834 25282
rect 28590 25230 28642 25282
rect 29038 25230 29090 25282
rect 29934 25230 29986 25282
rect 33070 25230 33122 25282
rect 37214 25230 37266 25282
rect 37550 25230 37602 25282
rect 38222 25230 38274 25282
rect 39902 25230 39954 25282
rect 40910 25230 40962 25282
rect 41806 25230 41858 25282
rect 45054 25230 45106 25282
rect 49870 25230 49922 25282
rect 58382 25230 58434 25282
rect 67566 25230 67618 25282
rect 68574 25230 68626 25282
rect 20534 25062 20586 25114
rect 20638 25062 20690 25114
rect 20742 25062 20794 25114
rect 39854 25062 39906 25114
rect 39958 25062 40010 25114
rect 40062 25062 40114 25114
rect 59174 25062 59226 25114
rect 59278 25062 59330 25114
rect 59382 25062 59434 25114
rect 78494 25062 78546 25114
rect 78598 25062 78650 25114
rect 78702 25062 78754 25114
rect 3726 24894 3778 24946
rect 9886 24894 9938 24946
rect 26014 24894 26066 24946
rect 27246 24894 27298 24946
rect 28926 24894 28978 24946
rect 29710 24894 29762 24946
rect 37102 24894 37154 24946
rect 38782 24894 38834 24946
rect 46622 24894 46674 24946
rect 47518 24894 47570 24946
rect 49534 24894 49586 24946
rect 52670 24894 52722 24946
rect 53006 24894 53058 24946
rect 55134 24894 55186 24946
rect 59278 24894 59330 24946
rect 63870 24894 63922 24946
rect 69134 24894 69186 24946
rect 69806 24894 69858 24946
rect 72158 24894 72210 24946
rect 74622 24894 74674 24946
rect 4734 24782 4786 24834
rect 5518 24782 5570 24834
rect 14590 24782 14642 24834
rect 14814 24782 14866 24834
rect 15486 24782 15538 24834
rect 17502 24782 17554 24834
rect 19630 24782 19682 24834
rect 19742 24782 19794 24834
rect 28142 24782 28194 24834
rect 31838 24782 31890 24834
rect 37550 24782 37602 24834
rect 40014 24782 40066 24834
rect 41358 24782 41410 24834
rect 45390 24782 45442 24834
rect 45838 24782 45890 24834
rect 57934 24782 57986 24834
rect 58382 24782 58434 24834
rect 60062 24782 60114 24834
rect 65438 24782 65490 24834
rect 65998 24782 66050 24834
rect 68686 24782 68738 24834
rect 72270 24782 72322 24834
rect 74286 24782 74338 24834
rect 76078 24782 76130 24834
rect 4062 24670 4114 24722
rect 4846 24670 4898 24722
rect 5854 24670 5906 24722
rect 9550 24670 9602 24722
rect 10558 24670 10610 24722
rect 15822 24670 15874 24722
rect 16718 24670 16770 24722
rect 18734 24670 18786 24722
rect 19182 24670 19234 24722
rect 19406 24670 19458 24722
rect 20302 24670 20354 24722
rect 20526 24670 20578 24722
rect 22318 24670 22370 24722
rect 23550 24670 23602 24722
rect 27918 24670 27970 24722
rect 28478 24670 28530 24722
rect 29038 24670 29090 24722
rect 33182 24670 33234 24722
rect 34078 24670 34130 24722
rect 36318 24670 36370 24722
rect 37662 24670 37714 24722
rect 37886 24670 37938 24722
rect 39230 24670 39282 24722
rect 39678 24670 39730 24722
rect 41470 24670 41522 24722
rect 42478 24670 42530 24722
rect 44718 24670 44770 24722
rect 45278 24670 45330 24722
rect 46174 24670 46226 24722
rect 46622 24670 46674 24722
rect 51102 24670 51154 24722
rect 51662 24670 51714 24722
rect 53902 24670 53954 24722
rect 55470 24670 55522 24722
rect 56590 24670 56642 24722
rect 57822 24670 57874 24722
rect 58158 24670 58210 24722
rect 59726 24670 59778 24722
rect 62190 24670 62242 24722
rect 63646 24670 63698 24722
rect 64878 24670 64930 24722
rect 65214 24670 65266 24722
rect 69022 24670 69074 24722
rect 69470 24670 69522 24722
rect 72606 24670 72658 24722
rect 73390 24670 73442 24722
rect 73726 24670 73778 24722
rect 75294 24670 75346 24722
rect 6302 24558 6354 24610
rect 11342 24558 11394 24610
rect 13470 24558 13522 24610
rect 16158 24558 16210 24610
rect 17726 24558 17778 24610
rect 20190 24558 20242 24610
rect 23886 24558 23938 24610
rect 26798 24558 26850 24610
rect 30158 24558 30210 24610
rect 30718 24558 30770 24610
rect 32174 24558 32226 24610
rect 33630 24558 33682 24610
rect 36766 24558 36818 24610
rect 38334 24558 38386 24610
rect 39790 24558 39842 24610
rect 41806 24558 41858 24610
rect 42702 24558 42754 24610
rect 43262 24558 43314 24610
rect 44046 24558 44098 24610
rect 50766 24558 50818 24610
rect 53566 24558 53618 24610
rect 56030 24558 56082 24610
rect 57150 24558 57202 24610
rect 58830 24558 58882 24610
rect 60398 24558 60450 24610
rect 60958 24558 61010 24610
rect 62750 24558 62802 24610
rect 71710 24558 71762 24610
rect 78206 24558 78258 24610
rect 13918 24446 13970 24498
rect 14254 24446 14306 24498
rect 19070 24446 19122 24498
rect 28926 24446 28978 24498
rect 36094 24446 36146 24498
rect 41358 24446 41410 24498
rect 54686 24446 54738 24498
rect 10874 24278 10926 24330
rect 10978 24278 11030 24330
rect 11082 24278 11134 24330
rect 30194 24278 30246 24330
rect 30298 24278 30350 24330
rect 30402 24278 30454 24330
rect 49514 24278 49566 24330
rect 49618 24278 49670 24330
rect 49722 24278 49774 24330
rect 68834 24278 68886 24330
rect 68938 24278 68990 24330
rect 69042 24278 69094 24330
rect 21422 24110 21474 24162
rect 22094 24110 22146 24162
rect 28366 24110 28418 24162
rect 31502 24110 31554 24162
rect 31838 24110 31890 24162
rect 34302 24110 34354 24162
rect 36318 24110 36370 24162
rect 61406 24110 61458 24162
rect 1934 23998 1986 24050
rect 4846 23998 4898 24050
rect 8654 23998 8706 24050
rect 16270 23998 16322 24050
rect 19854 23998 19906 24050
rect 21870 23998 21922 24050
rect 25230 23998 25282 24050
rect 26014 23998 26066 24050
rect 27470 23998 27522 24050
rect 29822 23998 29874 24050
rect 33854 23998 33906 24050
rect 39790 23998 39842 24050
rect 44158 23998 44210 24050
rect 45390 23998 45442 24050
rect 45950 23998 46002 24050
rect 49422 23998 49474 24050
rect 52222 23998 52274 24050
rect 52894 23998 52946 24050
rect 54126 23998 54178 24050
rect 56254 23998 56306 24050
rect 58718 23998 58770 24050
rect 61854 23998 61906 24050
rect 64766 23998 64818 24050
rect 72270 23998 72322 24050
rect 75406 23998 75458 24050
rect 4286 23886 4338 23938
rect 5742 23886 5794 23938
rect 9438 23886 9490 23938
rect 11678 23886 11730 23938
rect 15262 23886 15314 23938
rect 16718 23886 16770 23938
rect 17502 23886 17554 23938
rect 18510 23886 18562 23938
rect 19070 23886 19122 23938
rect 21310 23886 21362 23938
rect 23438 23886 23490 23938
rect 29710 23886 29762 23938
rect 32622 23886 32674 23938
rect 33406 23886 33458 23938
rect 34078 23886 34130 23938
rect 35534 23886 35586 23938
rect 35982 23886 36034 23938
rect 37662 23886 37714 23938
rect 38110 23886 38162 23938
rect 38222 23886 38274 23938
rect 38446 23886 38498 23938
rect 38782 23886 38834 23938
rect 39454 23886 39506 23938
rect 41694 23886 41746 23938
rect 42702 23886 42754 23938
rect 42926 23886 42978 23938
rect 43710 23886 43762 23938
rect 47854 23886 47906 23938
rect 48750 23886 48802 23938
rect 53230 23886 53282 23938
rect 54462 23886 54514 23938
rect 57598 23886 57650 23938
rect 58830 23886 58882 23938
rect 61630 23886 61682 23938
rect 62526 23886 62578 23938
rect 70030 23886 70082 23938
rect 70814 23886 70866 23938
rect 71038 23886 71090 23938
rect 72158 23886 72210 23938
rect 72718 23886 72770 23938
rect 73054 23886 73106 23938
rect 6526 23774 6578 23826
rect 9662 23774 9714 23826
rect 9998 23774 10050 23826
rect 11342 23774 11394 23826
rect 22766 23774 22818 23826
rect 22990 23774 23042 23826
rect 26350 23774 26402 23826
rect 28254 23774 28306 23826
rect 29486 23774 29538 23826
rect 30606 23774 30658 23826
rect 31054 23774 31106 23826
rect 32398 23774 32450 23826
rect 35310 23774 35362 23826
rect 41470 23774 41522 23826
rect 43262 23774 43314 23826
rect 43598 23774 43650 23826
rect 47518 23774 47570 23826
rect 55022 23774 55074 23826
rect 57374 23774 57426 23826
rect 59054 23774 59106 23826
rect 59390 23774 59442 23826
rect 59502 23774 59554 23826
rect 66446 23774 66498 23826
rect 69582 23774 69634 23826
rect 71598 23774 71650 23826
rect 72270 23774 72322 23826
rect 9102 23662 9154 23714
rect 13582 23662 13634 23714
rect 21422 23662 21474 23714
rect 22430 23662 22482 23714
rect 23102 23662 23154 23714
rect 23774 23662 23826 23714
rect 25790 23662 25842 23714
rect 26686 23662 26738 23714
rect 27022 23662 27074 23714
rect 28030 23662 28082 23714
rect 28366 23662 28418 23714
rect 37102 23662 37154 23714
rect 43038 23662 43090 23714
rect 50766 23662 50818 23714
rect 53566 23662 53618 23714
rect 54574 23662 54626 23714
rect 57710 23662 57762 23714
rect 57822 23662 57874 23714
rect 57934 23662 57986 23714
rect 58494 23662 58546 23714
rect 58606 23662 58658 23714
rect 59726 23662 59778 23714
rect 60622 23662 60674 23714
rect 64206 23662 64258 23714
rect 66782 23662 66834 23714
rect 69246 23662 69298 23714
rect 69918 23662 69970 23714
rect 72494 23662 72546 23714
rect 76526 23662 76578 23714
rect 20534 23494 20586 23546
rect 20638 23494 20690 23546
rect 20742 23494 20794 23546
rect 39854 23494 39906 23546
rect 39958 23494 40010 23546
rect 40062 23494 40114 23546
rect 59174 23494 59226 23546
rect 59278 23494 59330 23546
rect 59382 23494 59434 23546
rect 78494 23494 78546 23546
rect 78598 23494 78650 23546
rect 78702 23494 78754 23546
rect 6862 23326 6914 23378
rect 8654 23326 8706 23378
rect 15710 23326 15762 23378
rect 16270 23326 16322 23378
rect 18174 23326 18226 23378
rect 19630 23326 19682 23378
rect 22206 23326 22258 23378
rect 22430 23326 22482 23378
rect 22878 23326 22930 23378
rect 23438 23326 23490 23378
rect 24558 23326 24610 23378
rect 25342 23326 25394 23378
rect 27246 23326 27298 23378
rect 30494 23326 30546 23378
rect 31614 23326 31666 23378
rect 33518 23326 33570 23378
rect 33742 23326 33794 23378
rect 36094 23326 36146 23378
rect 40238 23326 40290 23378
rect 41470 23326 41522 23378
rect 42814 23326 42866 23378
rect 46174 23326 46226 23378
rect 47182 23326 47234 23378
rect 47518 23326 47570 23378
rect 50094 23326 50146 23378
rect 51326 23326 51378 23378
rect 51662 23326 51714 23378
rect 51998 23326 52050 23378
rect 52782 23326 52834 23378
rect 53118 23326 53170 23378
rect 60398 23326 60450 23378
rect 60622 23326 60674 23378
rect 61742 23326 61794 23378
rect 62974 23326 63026 23378
rect 65102 23326 65154 23378
rect 65662 23326 65714 23378
rect 70366 23326 70418 23378
rect 7198 23214 7250 23266
rect 15486 23214 15538 23266
rect 16046 23214 16098 23266
rect 19070 23214 19122 23266
rect 21982 23214 22034 23266
rect 22766 23214 22818 23266
rect 26238 23214 26290 23266
rect 28366 23214 28418 23266
rect 30382 23214 30434 23266
rect 36654 23214 36706 23266
rect 39678 23214 39730 23266
rect 42366 23214 42418 23266
rect 53006 23214 53058 23266
rect 55470 23214 55522 23266
rect 57150 23214 57202 23266
rect 59726 23214 59778 23266
rect 61182 23214 61234 23266
rect 63198 23214 63250 23266
rect 66782 23214 66834 23266
rect 71374 23214 71426 23266
rect 73166 23214 73218 23266
rect 76974 23214 77026 23266
rect 1822 23102 1874 23154
rect 15374 23102 15426 23154
rect 15934 23102 15986 23154
rect 18062 23102 18114 23154
rect 18734 23102 18786 23154
rect 25678 23102 25730 23154
rect 26686 23102 26738 23154
rect 27470 23102 27522 23154
rect 29598 23102 29650 23154
rect 30718 23102 30770 23154
rect 31054 23102 31106 23154
rect 31278 23102 31330 23154
rect 32062 23102 32114 23154
rect 32510 23102 32562 23154
rect 34190 23102 34242 23154
rect 34638 23102 34690 23154
rect 35534 23102 35586 23154
rect 36542 23102 36594 23154
rect 37214 23102 37266 23154
rect 39790 23102 39842 23154
rect 40126 23102 40178 23154
rect 40910 23102 40962 23154
rect 41246 23102 41298 23154
rect 42702 23102 42754 23154
rect 43038 23102 43090 23154
rect 45950 23102 46002 23154
rect 50654 23102 50706 23154
rect 50990 23102 51042 23154
rect 54238 23102 54290 23154
rect 56030 23102 56082 23154
rect 58158 23102 58210 23154
rect 58382 23102 58434 23154
rect 59502 23102 59554 23154
rect 60734 23102 60786 23154
rect 60958 23102 61010 23154
rect 61294 23102 61346 23154
rect 62638 23102 62690 23154
rect 63310 23102 63362 23154
rect 65998 23102 66050 23154
rect 70590 23102 70642 23154
rect 71150 23102 71202 23154
rect 72830 23102 72882 23154
rect 73614 23102 73666 23154
rect 76862 23102 76914 23154
rect 2494 22990 2546 23042
rect 4622 22990 4674 23042
rect 15038 22990 15090 23042
rect 16606 22990 16658 23042
rect 22094 22990 22146 23042
rect 24110 22990 24162 23042
rect 26014 22990 26066 23042
rect 29150 22990 29202 23042
rect 35310 22990 35362 23042
rect 38222 22990 38274 23042
rect 39006 22990 39058 23042
rect 41358 22990 41410 23042
rect 41918 22990 41970 23042
rect 43374 22990 43426 23042
rect 43822 22990 43874 23042
rect 44606 22990 44658 23042
rect 45054 22990 45106 23042
rect 45502 22990 45554 23042
rect 46734 22990 46786 23042
rect 49422 22990 49474 23042
rect 54126 22990 54178 23042
rect 58494 22990 58546 23042
rect 60174 22990 60226 23042
rect 62190 22990 62242 23042
rect 68910 22990 68962 23042
rect 71486 22990 71538 23042
rect 72494 22990 72546 23042
rect 74286 22990 74338 23042
rect 76414 22990 76466 23042
rect 34414 22878 34466 22930
rect 64878 22878 64930 22930
rect 65102 22878 65154 22930
rect 77646 22878 77698 22930
rect 77982 22878 78034 22930
rect 10874 22710 10926 22762
rect 10978 22710 11030 22762
rect 11082 22710 11134 22762
rect 30194 22710 30246 22762
rect 30298 22710 30350 22762
rect 30402 22710 30454 22762
rect 49514 22710 49566 22762
rect 49618 22710 49670 22762
rect 49722 22710 49774 22762
rect 68834 22710 68886 22762
rect 68938 22710 68990 22762
rect 69042 22710 69094 22762
rect 22206 22542 22258 22594
rect 26350 22542 26402 22594
rect 40462 22542 40514 22594
rect 51326 22542 51378 22594
rect 62302 22542 62354 22594
rect 66446 22542 66498 22594
rect 66782 22542 66834 22594
rect 68350 22542 68402 22594
rect 76638 22542 76690 22594
rect 2046 22430 2098 22482
rect 5742 22430 5794 22482
rect 19406 22430 19458 22482
rect 19854 22430 19906 22482
rect 20302 22430 20354 22482
rect 30830 22430 30882 22482
rect 35758 22430 35810 22482
rect 37214 22430 37266 22482
rect 39790 22430 39842 22482
rect 44942 22430 44994 22482
rect 46622 22430 46674 22482
rect 50206 22430 50258 22482
rect 51102 22430 51154 22482
rect 56142 22430 56194 22482
rect 58046 22430 58098 22482
rect 65774 22430 65826 22482
rect 69358 22430 69410 22482
rect 75630 22430 75682 22482
rect 4174 22318 4226 22370
rect 4958 22318 5010 22370
rect 17278 22318 17330 22370
rect 18174 22318 18226 22370
rect 18286 22318 18338 22370
rect 18510 22318 18562 22370
rect 18734 22318 18786 22370
rect 22094 22318 22146 22370
rect 23998 22318 24050 22370
rect 24446 22318 24498 22370
rect 25006 22318 25058 22370
rect 26462 22318 26514 22370
rect 26574 22318 26626 22370
rect 27470 22318 27522 22370
rect 27918 22318 27970 22370
rect 28254 22318 28306 22370
rect 28702 22318 28754 22370
rect 29150 22318 29202 22370
rect 29598 22318 29650 22370
rect 31390 22318 31442 22370
rect 32174 22318 32226 22370
rect 32734 22318 32786 22370
rect 33630 22318 33682 22370
rect 35422 22318 35474 22370
rect 36206 22318 36258 22370
rect 37102 22318 37154 22370
rect 39342 22318 39394 22370
rect 39902 22318 39954 22370
rect 41022 22318 41074 22370
rect 42142 22318 42194 22370
rect 42478 22318 42530 22370
rect 43262 22318 43314 22370
rect 44270 22318 44322 22370
rect 45054 22318 45106 22370
rect 45278 22318 45330 22370
rect 45502 22318 45554 22370
rect 46174 22318 46226 22370
rect 47070 22318 47122 22370
rect 48190 22318 48242 22370
rect 48974 22318 49026 22370
rect 54350 22318 54402 22370
rect 58270 22318 58322 22370
rect 60510 22318 60562 22370
rect 61854 22318 61906 22370
rect 63086 22318 63138 22370
rect 65102 22318 65154 22370
rect 65326 22318 65378 22370
rect 69022 22318 69074 22370
rect 69694 22318 69746 22370
rect 70366 22318 70418 22370
rect 72270 22318 72322 22370
rect 74846 22318 74898 22370
rect 78094 22318 78146 22370
rect 2830 22206 2882 22258
rect 3166 22206 3218 22258
rect 3838 22206 3890 22258
rect 4734 22206 4786 22258
rect 16270 22206 16322 22258
rect 16606 22206 16658 22258
rect 24558 22206 24610 22258
rect 25678 22206 25730 22258
rect 29934 22206 29986 22258
rect 30606 22206 30658 22258
rect 31166 22206 31218 22258
rect 32286 22206 32338 22258
rect 34638 22206 34690 22258
rect 36430 22206 36482 22258
rect 36990 22206 37042 22258
rect 40350 22206 40402 22258
rect 41694 22206 41746 22258
rect 42814 22206 42866 22258
rect 54910 22206 54962 22258
rect 59278 22206 59330 22258
rect 60846 22206 60898 22258
rect 67006 22206 67058 22258
rect 67454 22206 67506 22258
rect 68462 22206 68514 22258
rect 69358 22206 69410 22258
rect 71598 22262 71650 22314
rect 69918 22206 69970 22258
rect 73390 22206 73442 22258
rect 74174 22206 74226 22258
rect 76862 22206 76914 22258
rect 77198 22206 77250 22258
rect 11902 22094 11954 22146
rect 12238 22094 12290 22146
rect 12686 22094 12738 22146
rect 13470 22094 13522 22146
rect 13806 22094 13858 22146
rect 14254 22094 14306 22146
rect 16830 22094 16882 22146
rect 16942 22094 16994 22146
rect 17054 22094 17106 22146
rect 18398 22094 18450 22146
rect 22206 22094 22258 22146
rect 22878 22094 22930 22146
rect 23550 22094 23602 22146
rect 25790 22094 25842 22146
rect 26014 22094 26066 22146
rect 30718 22094 30770 22146
rect 30942 22094 30994 22146
rect 41134 22094 41186 22146
rect 43710 22094 43762 22146
rect 44942 22094 44994 22146
rect 47182 22094 47234 22146
rect 49758 22094 49810 22146
rect 50878 22094 50930 22146
rect 51662 22094 51714 22146
rect 52222 22094 52274 22146
rect 54462 22094 54514 22146
rect 57486 22094 57538 22146
rect 61070 22094 61122 22146
rect 68686 22094 68738 22146
rect 69470 22094 69522 22146
rect 75070 22094 75122 22146
rect 76302 22094 76354 22146
rect 77870 22094 77922 22146
rect 20534 21926 20586 21978
rect 20638 21926 20690 21978
rect 20742 21926 20794 21978
rect 39854 21926 39906 21978
rect 39958 21926 40010 21978
rect 40062 21926 40114 21978
rect 59174 21926 59226 21978
rect 59278 21926 59330 21978
rect 59382 21926 59434 21978
rect 78494 21926 78546 21978
rect 78598 21926 78650 21978
rect 78702 21926 78754 21978
rect 2158 21758 2210 21810
rect 12686 21758 12738 21810
rect 13470 21758 13522 21810
rect 14142 21758 14194 21810
rect 14478 21758 14530 21810
rect 15150 21758 15202 21810
rect 16606 21758 16658 21810
rect 18510 21758 18562 21810
rect 19966 21758 20018 21810
rect 22990 21758 23042 21810
rect 23998 21758 24050 21810
rect 24110 21758 24162 21810
rect 27806 21758 27858 21810
rect 29598 21758 29650 21810
rect 29934 21758 29986 21810
rect 31054 21758 31106 21810
rect 31950 21758 32002 21810
rect 38782 21758 38834 21810
rect 41022 21758 41074 21810
rect 41918 21758 41970 21810
rect 42366 21758 42418 21810
rect 46622 21758 46674 21810
rect 47966 21758 48018 21810
rect 50318 21758 50370 21810
rect 50878 21758 50930 21810
rect 51214 21758 51266 21810
rect 51998 21758 52050 21810
rect 52334 21758 52386 21810
rect 59726 21758 59778 21810
rect 59838 21758 59890 21810
rect 60062 21758 60114 21810
rect 64542 21758 64594 21810
rect 65326 21758 65378 21810
rect 66894 21758 66946 21810
rect 72606 21758 72658 21810
rect 72718 21758 72770 21810
rect 73502 21758 73554 21810
rect 74062 21758 74114 21810
rect 74398 21758 74450 21810
rect 1710 21646 1762 21698
rect 15598 21646 15650 21698
rect 18734 21646 18786 21698
rect 19518 21646 19570 21698
rect 20302 21646 20354 21698
rect 24334 21646 24386 21698
rect 26686 21646 26738 21698
rect 29822 21646 29874 21698
rect 36990 21646 37042 21698
rect 38446 21646 38498 21698
rect 39230 21646 39282 21698
rect 51774 21646 51826 21698
rect 57598 21646 57650 21698
rect 59502 21646 59554 21698
rect 64878 21646 64930 21698
rect 65550 21646 65602 21698
rect 66222 21646 66274 21698
rect 67118 21646 67170 21698
rect 67678 21646 67730 21698
rect 70478 21646 70530 21698
rect 71710 21646 71762 21698
rect 73726 21646 73778 21698
rect 74734 21646 74786 21698
rect 75854 21646 75906 21698
rect 2382 21534 2434 21586
rect 2830 21534 2882 21586
rect 6190 21534 6242 21586
rect 10334 21534 10386 21586
rect 10558 21534 10610 21586
rect 10670 21534 10722 21586
rect 11118 21534 11170 21586
rect 11566 21534 11618 21586
rect 13694 21534 13746 21586
rect 15710 21534 15762 21586
rect 15934 21534 15986 21586
rect 18286 21534 18338 21586
rect 18398 21534 18450 21586
rect 18622 21534 18674 21586
rect 19294 21534 19346 21586
rect 19406 21534 19458 21586
rect 20638 21534 20690 21586
rect 23438 21534 23490 21586
rect 23774 21534 23826 21586
rect 23886 21534 23938 21586
rect 26126 21534 26178 21586
rect 26462 21534 26514 21586
rect 27470 21534 27522 21586
rect 27918 21534 27970 21586
rect 29038 21534 29090 21586
rect 29262 21534 29314 21586
rect 30382 21534 30434 21586
rect 31390 21534 31442 21586
rect 34750 21534 34802 21586
rect 35982 21534 36034 21586
rect 36430 21534 36482 21586
rect 38670 21534 38722 21586
rect 38894 21534 38946 21586
rect 40126 21534 40178 21586
rect 42814 21534 42866 21586
rect 43374 21534 43426 21586
rect 43598 21534 43650 21586
rect 44718 21534 44770 21586
rect 45166 21534 45218 21586
rect 45614 21534 45666 21586
rect 47518 21534 47570 21586
rect 47742 21534 47794 21586
rect 48078 21534 48130 21586
rect 48862 21534 48914 21586
rect 49310 21534 49362 21586
rect 49870 21534 49922 21586
rect 50990 21534 51042 21586
rect 51326 21534 51378 21586
rect 52222 21534 52274 21586
rect 58158 21534 58210 21586
rect 58382 21534 58434 21586
rect 59950 21534 60002 21586
rect 63870 21534 63922 21586
rect 65326 21534 65378 21586
rect 67230 21534 67282 21586
rect 70814 21534 70866 21586
rect 71262 21534 71314 21586
rect 72270 21534 72322 21586
rect 72494 21534 72546 21586
rect 72942 21534 72994 21586
rect 75182 21534 75234 21586
rect 3614 21422 3666 21474
rect 5742 21422 5794 21474
rect 6862 21422 6914 21474
rect 8990 21422 9042 21474
rect 11342 21422 11394 21474
rect 11454 21422 11506 21474
rect 12350 21422 12402 21474
rect 13246 21422 13298 21474
rect 17838 21422 17890 21474
rect 21086 21422 21138 21474
rect 22094 21422 22146 21474
rect 22430 21422 22482 21474
rect 25566 21422 25618 21474
rect 28590 21422 28642 21474
rect 30270 21422 30322 21474
rect 32286 21422 32338 21474
rect 33182 21422 33234 21474
rect 34302 21422 34354 21474
rect 36878 21422 36930 21474
rect 39678 21422 39730 21474
rect 41470 21422 41522 21474
rect 45502 21422 45554 21474
rect 47182 21422 47234 21474
rect 47854 21422 47906 21474
rect 50878 21422 50930 21474
rect 52334 21422 52386 21474
rect 58494 21422 58546 21474
rect 60622 21422 60674 21474
rect 60958 21422 61010 21474
rect 63086 21422 63138 21474
rect 71374 21422 71426 21474
rect 77982 21422 78034 21474
rect 1822 21310 1874 21362
rect 21870 21310 21922 21362
rect 22542 21310 22594 21362
rect 22990 21310 23042 21362
rect 41470 21310 41522 21362
rect 41694 21310 41746 21362
rect 44158 21310 44210 21362
rect 45950 21310 46002 21362
rect 10874 21142 10926 21194
rect 10978 21142 11030 21194
rect 11082 21142 11134 21194
rect 30194 21142 30246 21194
rect 30298 21142 30350 21194
rect 30402 21142 30454 21194
rect 49514 21142 49566 21194
rect 49618 21142 49670 21194
rect 49722 21142 49774 21194
rect 68834 21142 68886 21194
rect 68938 21142 68990 21194
rect 69042 21142 69094 21194
rect 2718 20974 2770 21026
rect 6190 20974 6242 21026
rect 24446 20974 24498 21026
rect 25118 20974 25170 21026
rect 25342 20974 25394 21026
rect 25566 20974 25618 21026
rect 46622 20974 46674 21026
rect 47182 20974 47234 21026
rect 73614 20974 73666 21026
rect 11678 20862 11730 20914
rect 16382 20862 16434 20914
rect 17278 20862 17330 20914
rect 17838 20862 17890 20914
rect 20750 20862 20802 20914
rect 21422 20862 21474 20914
rect 22990 20862 23042 20914
rect 24222 20862 24274 20914
rect 24670 20862 24722 20914
rect 25118 20862 25170 20914
rect 25678 20862 25730 20914
rect 27134 20862 27186 20914
rect 28254 20862 28306 20914
rect 31166 20862 31218 20914
rect 31614 20862 31666 20914
rect 34750 20862 34802 20914
rect 39006 20862 39058 20914
rect 41022 20862 41074 20914
rect 42702 20862 42754 20914
rect 43598 20862 43650 20914
rect 45166 20862 45218 20914
rect 46846 20862 46898 20914
rect 47182 20862 47234 20914
rect 56814 20862 56866 20914
rect 59054 20862 59106 20914
rect 59390 20862 59442 20914
rect 67230 20862 67282 20914
rect 70030 20862 70082 20914
rect 1822 20750 1874 20802
rect 6974 20750 7026 20802
rect 7982 20750 8034 20802
rect 9998 20750 10050 20802
rect 10446 20750 10498 20802
rect 10782 20750 10834 20802
rect 11230 20750 11282 20802
rect 11454 20750 11506 20802
rect 13582 20750 13634 20802
rect 16942 20750 16994 20802
rect 21310 20750 21362 20802
rect 21534 20750 21586 20802
rect 21870 20750 21922 20802
rect 25902 20750 25954 20802
rect 27470 20750 27522 20802
rect 28366 20750 28418 20802
rect 29486 20750 29538 20802
rect 30830 20750 30882 20802
rect 32398 20750 32450 20802
rect 33742 20750 33794 20802
rect 36094 20750 36146 20802
rect 37326 20750 37378 20802
rect 41806 20750 41858 20802
rect 42366 20750 42418 20802
rect 44942 20750 44994 20802
rect 45278 20750 45330 20802
rect 45390 20750 45442 20802
rect 48750 20750 48802 20802
rect 49870 20750 49922 20802
rect 50766 20750 50818 20802
rect 52670 20750 52722 20802
rect 53678 20750 53730 20802
rect 56590 20750 56642 20802
rect 58046 20750 58098 20802
rect 61406 20750 61458 20802
rect 62078 20750 62130 20802
rect 62414 20750 62466 20802
rect 62862 20750 62914 20802
rect 63758 20750 63810 20802
rect 64430 20750 64482 20802
rect 71374 20750 71426 20802
rect 73726 20750 73778 20802
rect 4622 20638 4674 20690
rect 4958 20638 5010 20690
rect 5854 20638 5906 20690
rect 6862 20638 6914 20690
rect 7758 20638 7810 20690
rect 14254 20638 14306 20690
rect 16718 20638 16770 20690
rect 21758 20638 21810 20690
rect 22430 20638 22482 20690
rect 22542 20638 22594 20690
rect 26238 20638 26290 20690
rect 28142 20638 28194 20690
rect 29822 20638 29874 20690
rect 33294 20638 33346 20690
rect 34638 20638 34690 20690
rect 38222 20638 38274 20690
rect 40126 20638 40178 20690
rect 40238 20638 40290 20690
rect 43038 20638 43090 20690
rect 49086 20638 49138 20690
rect 50206 20638 50258 20690
rect 50318 20638 50370 20690
rect 50878 20638 50930 20690
rect 51774 20638 51826 20690
rect 51886 20638 51938 20690
rect 55582 20638 55634 20690
rect 63198 20638 63250 20690
rect 63982 20638 64034 20690
rect 65102 20638 65154 20690
rect 72830 20638 72882 20690
rect 10110 20526 10162 20578
rect 10670 20526 10722 20578
rect 11678 20526 11730 20578
rect 12238 20526 12290 20578
rect 12574 20526 12626 20578
rect 17166 20526 17218 20578
rect 17278 20526 17330 20578
rect 18286 20526 18338 20578
rect 18958 20526 19010 20578
rect 19294 20526 19346 20578
rect 19742 20526 19794 20578
rect 22206 20526 22258 20578
rect 23550 20526 23602 20578
rect 26574 20526 26626 20578
rect 30270 20526 30322 20578
rect 38670 20526 38722 20578
rect 40462 20526 40514 20578
rect 41470 20526 41522 20578
rect 43934 20526 43986 20578
rect 45054 20526 45106 20578
rect 45950 20526 46002 20578
rect 47630 20526 47682 20578
rect 49310 20526 49362 20578
rect 50542 20526 50594 20578
rect 51102 20526 51154 20578
rect 52110 20526 52162 20578
rect 52782 20526 52834 20578
rect 53006 20526 53058 20578
rect 53454 20526 53506 20578
rect 55134 20526 55186 20578
rect 58270 20526 58322 20578
rect 60958 20526 61010 20578
rect 61630 20526 61682 20578
rect 74174 20526 74226 20578
rect 75294 20526 75346 20578
rect 76302 20526 76354 20578
rect 20534 20358 20586 20410
rect 20638 20358 20690 20410
rect 20742 20358 20794 20410
rect 39854 20358 39906 20410
rect 39958 20358 40010 20410
rect 40062 20358 40114 20410
rect 59174 20358 59226 20410
rect 59278 20358 59330 20410
rect 59382 20358 59434 20410
rect 78494 20358 78546 20410
rect 78598 20358 78650 20410
rect 78702 20358 78754 20410
rect 7758 20190 7810 20242
rect 25790 20190 25842 20242
rect 26350 20190 26402 20242
rect 30158 20190 30210 20242
rect 44494 20190 44546 20242
rect 49086 20190 49138 20242
rect 49870 20190 49922 20242
rect 51886 20190 51938 20242
rect 56702 20190 56754 20242
rect 69022 20190 69074 20242
rect 69470 20190 69522 20242
rect 3166 20078 3218 20130
rect 3502 20078 3554 20130
rect 7310 20078 7362 20130
rect 8766 20078 8818 20130
rect 9998 20078 10050 20130
rect 10446 20078 10498 20130
rect 16270 20078 16322 20130
rect 16718 20078 16770 20130
rect 28366 20078 28418 20130
rect 32174 20078 32226 20130
rect 32510 20078 32562 20130
rect 33518 20078 33570 20130
rect 33742 20078 33794 20130
rect 33966 20078 34018 20130
rect 36318 20078 36370 20130
rect 42478 20078 42530 20130
rect 42702 20078 42754 20130
rect 43262 20078 43314 20130
rect 44830 20078 44882 20130
rect 45278 20078 45330 20130
rect 45838 20078 45890 20130
rect 48750 20078 48802 20130
rect 48862 20078 48914 20130
rect 49422 20078 49474 20130
rect 50990 20078 51042 20130
rect 55022 20078 55074 20130
rect 59166 20078 59218 20130
rect 61182 20078 61234 20130
rect 64542 20078 64594 20130
rect 65102 20078 65154 20130
rect 65550 20078 65602 20130
rect 69694 20078 69746 20130
rect 70590 20078 70642 20130
rect 8094 19966 8146 20018
rect 8878 19966 8930 20018
rect 9662 19966 9714 20018
rect 10110 19966 10162 20018
rect 10894 19966 10946 20018
rect 11678 19966 11730 20018
rect 13022 19966 13074 20018
rect 13470 19966 13522 20018
rect 14478 19966 14530 20018
rect 16046 19966 16098 20018
rect 16382 19966 16434 20018
rect 23102 19966 23154 20018
rect 27134 19966 27186 20018
rect 27806 19966 27858 20018
rect 29598 19966 29650 20018
rect 31054 19966 31106 20018
rect 34526 19966 34578 20018
rect 35422 19966 35474 20018
rect 37550 19966 37602 20018
rect 37774 19966 37826 20018
rect 40238 19966 40290 20018
rect 41918 19966 41970 20018
rect 50878 19966 50930 20018
rect 52894 19966 52946 20018
rect 54350 19966 54402 20018
rect 59950 19966 60002 20018
rect 60846 19966 60898 20018
rect 64878 19966 64930 20018
rect 66110 19966 66162 20018
rect 66670 19966 66722 20018
rect 69582 19966 69634 20018
rect 69806 19966 69858 20018
rect 70030 19966 70082 20018
rect 70814 19966 70866 20018
rect 71262 19966 71314 20018
rect 72718 19966 72770 20018
rect 75742 19966 75794 20018
rect 3950 19854 4002 19906
rect 4398 19854 4450 19906
rect 14814 19854 14866 19906
rect 17502 19854 17554 19906
rect 17950 19854 18002 19906
rect 20190 19854 20242 19906
rect 22318 19854 22370 19906
rect 23550 19854 23602 19906
rect 23998 19854 24050 19906
rect 26686 19854 26738 19906
rect 31502 19854 31554 19906
rect 35534 19854 35586 19906
rect 41358 19854 41410 19906
rect 43710 19854 43762 19906
rect 50318 19854 50370 19906
rect 55470 19854 55522 19906
rect 56030 19854 56082 19906
rect 57038 19854 57090 19906
rect 63870 19854 63922 19906
rect 72494 19854 72546 19906
rect 77982 19854 78034 19906
rect 3838 19742 3890 19794
rect 10558 19742 10610 19794
rect 11006 19742 11058 19794
rect 15038 19742 15090 19794
rect 16830 19742 16882 19794
rect 17390 19742 17442 19794
rect 17838 19742 17890 19794
rect 23438 19742 23490 19794
rect 33182 19742 33234 19794
rect 38782 19742 38834 19794
rect 42814 19742 42866 19794
rect 71598 19742 71650 19794
rect 75070 19742 75122 19794
rect 10874 19574 10926 19626
rect 10978 19574 11030 19626
rect 11082 19574 11134 19626
rect 30194 19574 30246 19626
rect 30298 19574 30350 19626
rect 30402 19574 30454 19626
rect 49514 19574 49566 19626
rect 49618 19574 49670 19626
rect 49722 19574 49774 19626
rect 68834 19574 68886 19626
rect 68938 19574 68990 19626
rect 69042 19574 69094 19626
rect 18174 19406 18226 19458
rect 23102 19406 23154 19458
rect 27470 19406 27522 19458
rect 29934 19406 29986 19458
rect 58270 19406 58322 19458
rect 69246 19406 69298 19458
rect 2718 19294 2770 19346
rect 4846 19294 4898 19346
rect 13806 19294 13858 19346
rect 14702 19294 14754 19346
rect 21758 19294 21810 19346
rect 22318 19294 22370 19346
rect 22654 19294 22706 19346
rect 27022 19294 27074 19346
rect 28590 19294 28642 19346
rect 33742 19294 33794 19346
rect 38894 19294 38946 19346
rect 40574 19294 40626 19346
rect 51438 19294 51490 19346
rect 53454 19294 53506 19346
rect 55582 19294 55634 19346
rect 61070 19294 61122 19346
rect 2046 19182 2098 19234
rect 12126 19182 12178 19234
rect 15262 19182 15314 19234
rect 15710 19182 15762 19234
rect 16494 19182 16546 19234
rect 16942 19182 16994 19234
rect 17278 19182 17330 19234
rect 18622 19182 18674 19234
rect 22206 19182 22258 19234
rect 22878 19182 22930 19234
rect 23326 19182 23378 19234
rect 26126 19182 26178 19234
rect 26574 19182 26626 19234
rect 27358 19182 27410 19234
rect 27806 19182 27858 19234
rect 28142 19182 28194 19234
rect 29038 19182 29090 19234
rect 29374 19182 29426 19234
rect 29710 19182 29762 19234
rect 30270 19182 30322 19234
rect 33182 19182 33234 19234
rect 34078 19182 34130 19234
rect 35422 19182 35474 19234
rect 36430 19182 36482 19234
rect 39118 19182 39170 19234
rect 40686 19182 40738 19234
rect 42142 19182 42194 19234
rect 42590 19182 42642 19234
rect 43486 19182 43538 19234
rect 43934 19182 43986 19234
rect 47070 19182 47122 19234
rect 52782 19182 52834 19234
rect 56702 19182 56754 19234
rect 57262 19182 57314 19234
rect 57822 19182 57874 19234
rect 58606 19182 58658 19234
rect 59278 19182 59330 19234
rect 61854 19182 61906 19234
rect 68910 19182 68962 19234
rect 10894 19070 10946 19122
rect 11342 19070 11394 19122
rect 11790 19070 11842 19122
rect 12350 19070 12402 19122
rect 14814 19070 14866 19122
rect 16270 19070 16322 19122
rect 18286 19070 18338 19122
rect 18958 19070 19010 19122
rect 21646 19070 21698 19122
rect 24894 19070 24946 19122
rect 27918 19070 27970 19122
rect 35646 19070 35698 19122
rect 41470 19070 41522 19122
rect 43038 19070 43090 19122
rect 44942 19070 44994 19122
rect 47518 19070 47570 19122
rect 56814 19070 56866 19122
rect 59390 19070 59442 19122
rect 61406 19070 61458 19122
rect 9214 18958 9266 19010
rect 12686 18958 12738 19010
rect 14366 18958 14418 19010
rect 14590 18958 14642 19010
rect 16046 18958 16098 19010
rect 16382 18958 16434 19010
rect 18846 18958 18898 19010
rect 20750 18958 20802 19010
rect 21870 18958 21922 19010
rect 23774 18958 23826 19010
rect 24222 18958 24274 19010
rect 25230 18958 25282 19010
rect 25678 18958 25730 19010
rect 29598 18958 29650 19010
rect 30046 18958 30098 19010
rect 37326 18958 37378 19010
rect 38110 18958 38162 19010
rect 41582 18958 41634 19010
rect 56142 18958 56194 19010
rect 56926 18958 56978 19010
rect 67902 18958 67954 19010
rect 68350 18958 68402 19010
rect 70254 19294 70306 19346
rect 71150 19294 71202 19346
rect 74958 19294 75010 19346
rect 76638 19294 76690 19346
rect 78094 19294 78146 19346
rect 70366 19182 70418 19234
rect 70590 19182 70642 19234
rect 73950 19182 74002 19234
rect 76190 19182 76242 19234
rect 69582 19070 69634 19122
rect 69694 19070 69746 19122
rect 70814 19070 70866 19122
rect 73278 19070 73330 19122
rect 75630 19070 75682 19122
rect 77646 19070 77698 19122
rect 77982 19070 78034 19122
rect 69358 18958 69410 19010
rect 69918 18958 69970 19010
rect 70254 18958 70306 19010
rect 74398 18958 74450 19010
rect 75294 18958 75346 19010
rect 75518 18958 75570 19010
rect 77198 18958 77250 19010
rect 77422 18958 77474 19010
rect 77534 18958 77586 19010
rect 20534 18790 20586 18842
rect 20638 18790 20690 18842
rect 20742 18790 20794 18842
rect 39854 18790 39906 18842
rect 39958 18790 40010 18842
rect 40062 18790 40114 18842
rect 59174 18790 59226 18842
rect 59278 18790 59330 18842
rect 59382 18790 59434 18842
rect 78494 18790 78546 18842
rect 78598 18790 78650 18842
rect 78702 18790 78754 18842
rect 4734 18622 4786 18674
rect 19966 18622 20018 18674
rect 21870 18622 21922 18674
rect 28702 18622 28754 18674
rect 36430 18622 36482 18674
rect 42478 18622 42530 18674
rect 69582 18622 69634 18674
rect 69694 18622 69746 18674
rect 70590 18622 70642 18674
rect 5854 18510 5906 18562
rect 17726 18510 17778 18562
rect 19070 18510 19122 18562
rect 20750 18510 20802 18562
rect 20862 18510 20914 18562
rect 22542 18510 22594 18562
rect 26014 18510 26066 18562
rect 34974 18510 35026 18562
rect 35534 18510 35586 18562
rect 37438 18510 37490 18562
rect 43486 18510 43538 18562
rect 48974 18510 49026 18562
rect 54910 18510 54962 18562
rect 55582 18510 55634 18562
rect 56814 18510 56866 18562
rect 60734 18510 60786 18562
rect 62190 18510 62242 18562
rect 63086 18510 63138 18562
rect 70478 18510 70530 18562
rect 71374 18510 71426 18562
rect 72830 18510 72882 18562
rect 77422 18510 77474 18562
rect 3838 18398 3890 18450
rect 5742 18398 5794 18450
rect 6414 18398 6466 18450
rect 11902 18398 11954 18450
rect 12910 18398 12962 18450
rect 13134 18398 13186 18450
rect 14590 18398 14642 18450
rect 17390 18398 17442 18450
rect 18062 18398 18114 18450
rect 19630 18398 19682 18450
rect 20190 18398 20242 18450
rect 20414 18398 20466 18450
rect 21086 18398 21138 18450
rect 21422 18398 21474 18450
rect 21646 18398 21698 18450
rect 23438 18398 23490 18450
rect 23886 18398 23938 18450
rect 23998 18398 24050 18450
rect 26350 18398 26402 18450
rect 27694 18398 27746 18450
rect 29038 18398 29090 18450
rect 29934 18398 29986 18450
rect 30494 18398 30546 18450
rect 34302 18398 34354 18450
rect 34638 18398 34690 18450
rect 36542 18398 36594 18450
rect 37998 18398 38050 18450
rect 39230 18398 39282 18450
rect 40014 18398 40066 18450
rect 42030 18398 42082 18450
rect 43598 18398 43650 18450
rect 44270 18398 44322 18450
rect 44718 18398 44770 18450
rect 45390 18398 45442 18450
rect 48750 18398 48802 18450
rect 53790 18398 53842 18450
rect 54126 18398 54178 18450
rect 54686 18398 54738 18450
rect 55358 18398 55410 18450
rect 55694 18398 55746 18450
rect 55806 18398 55858 18450
rect 56030 18398 56082 18450
rect 56478 18398 56530 18450
rect 56702 18398 56754 18450
rect 57262 18398 57314 18450
rect 58046 18398 58098 18450
rect 60510 18398 60562 18450
rect 61966 18398 62018 18450
rect 62862 18398 62914 18450
rect 65326 18398 65378 18450
rect 66670 18398 66722 18450
rect 67566 18398 67618 18450
rect 68126 18398 68178 18450
rect 69358 18398 69410 18450
rect 69470 18398 69522 18450
rect 69918 18398 69970 18450
rect 70814 18398 70866 18450
rect 71150 18398 71202 18450
rect 73054 18398 73106 18450
rect 73950 18398 74002 18450
rect 78094 18398 78146 18450
rect 1934 18286 1986 18338
rect 14702 18286 14754 18338
rect 16158 18286 16210 18338
rect 16830 18286 16882 18338
rect 20302 18286 20354 18338
rect 24670 18286 24722 18338
rect 26910 18286 26962 18338
rect 27358 18286 27410 18338
rect 28030 18286 28082 18338
rect 29486 18286 29538 18338
rect 40350 18286 40402 18338
rect 41022 18286 41074 18338
rect 42926 18286 42978 18338
rect 46062 18286 46114 18338
rect 48190 18286 48242 18338
rect 49422 18286 49474 18338
rect 53454 18286 53506 18338
rect 60062 18286 60114 18338
rect 61182 18286 61234 18338
rect 63534 18286 63586 18338
rect 64990 18286 65042 18338
rect 65662 18286 65714 18338
rect 67118 18286 67170 18338
rect 68574 18286 68626 18338
rect 72718 18286 72770 18338
rect 75294 18286 75346 18338
rect 5070 18174 5122 18226
rect 15038 18174 15090 18226
rect 18622 18174 18674 18226
rect 21982 18174 22034 18226
rect 22654 18174 22706 18226
rect 26574 18174 26626 18226
rect 26910 18174 26962 18226
rect 27358 18174 27410 18226
rect 45054 18174 45106 18226
rect 61518 18174 61570 18226
rect 10874 18006 10926 18058
rect 10978 18006 11030 18058
rect 11082 18006 11134 18058
rect 30194 18006 30246 18058
rect 30298 18006 30350 18058
rect 30402 18006 30454 18058
rect 49514 18006 49566 18058
rect 49618 18006 49670 18058
rect 49722 18006 49774 18058
rect 68834 18006 68886 18058
rect 68938 18006 68990 18058
rect 69042 18006 69094 18058
rect 17390 17838 17442 17890
rect 17502 17838 17554 17890
rect 17726 17838 17778 17890
rect 20078 17838 20130 17890
rect 22542 17838 22594 17890
rect 23326 17838 23378 17890
rect 40686 17838 40738 17890
rect 53118 17838 53170 17890
rect 63870 17838 63922 17890
rect 5070 17726 5122 17778
rect 6078 17726 6130 17778
rect 12574 17726 12626 17778
rect 13582 17726 13634 17778
rect 14702 17726 14754 17778
rect 15374 17726 15426 17778
rect 16718 17726 16770 17778
rect 18846 17726 18898 17778
rect 21534 17726 21586 17778
rect 22878 17726 22930 17778
rect 23102 17726 23154 17778
rect 25006 17726 25058 17778
rect 29710 17726 29762 17778
rect 33406 17726 33458 17778
rect 37550 17726 37602 17778
rect 40574 17726 40626 17778
rect 45502 17726 45554 17778
rect 49310 17726 49362 17778
rect 54462 17726 54514 17778
rect 57150 17726 57202 17778
rect 57822 17726 57874 17778
rect 58830 17726 58882 17778
rect 61294 17726 61346 17778
rect 63422 17726 63474 17778
rect 65998 17726 66050 17778
rect 67006 17726 67058 17778
rect 68798 17726 68850 17778
rect 69582 17726 69634 17778
rect 73054 17726 73106 17778
rect 75518 17726 75570 17778
rect 2158 17614 2210 17666
rect 6750 17614 6802 17666
rect 12462 17614 12514 17666
rect 14254 17614 14306 17666
rect 15710 17614 15762 17666
rect 20302 17614 20354 17666
rect 20750 17614 20802 17666
rect 29262 17614 29314 17666
rect 31614 17614 31666 17666
rect 33294 17614 33346 17666
rect 34302 17614 34354 17666
rect 34638 17614 34690 17666
rect 35198 17614 35250 17666
rect 36206 17614 36258 17666
rect 36990 17614 37042 17666
rect 40238 17614 40290 17666
rect 41022 17614 41074 17666
rect 43262 17614 43314 17666
rect 43710 17614 43762 17666
rect 46398 17614 46450 17666
rect 47966 17614 48018 17666
rect 48750 17614 48802 17666
rect 53678 17614 53730 17666
rect 55918 17614 55970 17666
rect 56926 17614 56978 17666
rect 57934 17614 57986 17666
rect 58718 17614 58770 17666
rect 58942 17614 58994 17666
rect 59390 17614 59442 17666
rect 60622 17614 60674 17666
rect 64206 17614 64258 17666
rect 64654 17614 64706 17666
rect 65550 17614 65602 17666
rect 69806 17614 69858 17666
rect 71150 17614 71202 17666
rect 71486 17614 71538 17666
rect 72270 17614 72322 17666
rect 74622 17614 74674 17666
rect 76414 17614 76466 17666
rect 76750 17614 76802 17666
rect 76974 17614 77026 17666
rect 2942 17502 2994 17554
rect 6638 17502 6690 17554
rect 7646 17502 7698 17554
rect 11678 17502 11730 17554
rect 12014 17502 12066 17554
rect 15934 17502 15986 17554
rect 16158 17502 16210 17554
rect 16494 17502 16546 17554
rect 16718 17502 16770 17554
rect 16942 17502 16994 17554
rect 18286 17502 18338 17554
rect 18622 17502 18674 17554
rect 19070 17502 19122 17554
rect 19742 17502 19794 17554
rect 22766 17502 22818 17554
rect 26798 17502 26850 17554
rect 27918 17502 27970 17554
rect 30718 17502 30770 17554
rect 31278 17502 31330 17554
rect 33630 17502 33682 17554
rect 34190 17502 34242 17554
rect 35422 17502 35474 17554
rect 36094 17502 36146 17554
rect 38670 17502 38722 17554
rect 39342 17502 39394 17554
rect 44270 17502 44322 17554
rect 47182 17502 47234 17554
rect 47630 17502 47682 17554
rect 48638 17502 48690 17554
rect 51326 17502 51378 17554
rect 52782 17502 52834 17554
rect 53902 17502 53954 17554
rect 55470 17502 55522 17554
rect 58382 17502 58434 17554
rect 64990 17502 65042 17554
rect 73726 17502 73778 17554
rect 77198 17502 77250 17554
rect 77310 17502 77362 17554
rect 5742 17390 5794 17442
rect 7310 17390 7362 17442
rect 8094 17390 8146 17442
rect 12910 17390 12962 17442
rect 16270 17390 16322 17442
rect 18846 17390 18898 17442
rect 19966 17390 20018 17442
rect 22094 17390 22146 17442
rect 23774 17390 23826 17442
rect 24110 17390 24162 17442
rect 24558 17390 24610 17442
rect 25566 17390 25618 17442
rect 27134 17390 27186 17442
rect 27694 17390 27746 17442
rect 28254 17390 28306 17442
rect 32174 17390 32226 17442
rect 44046 17390 44098 17442
rect 44382 17390 44434 17442
rect 46846 17390 46898 17442
rect 50990 17390 51042 17442
rect 57822 17390 57874 17442
rect 58158 17390 58210 17442
rect 59166 17390 59218 17442
rect 66558 17390 66610 17442
rect 67902 17390 67954 17442
rect 68350 17390 68402 17442
rect 75182 17390 75234 17442
rect 75630 17390 75682 17442
rect 76190 17390 76242 17442
rect 76302 17390 76354 17442
rect 20534 17222 20586 17274
rect 20638 17222 20690 17274
rect 20742 17222 20794 17274
rect 39854 17222 39906 17274
rect 39958 17222 40010 17274
rect 40062 17222 40114 17274
rect 59174 17222 59226 17274
rect 59278 17222 59330 17274
rect 59382 17222 59434 17274
rect 78494 17222 78546 17274
rect 78598 17222 78650 17274
rect 78702 17222 78754 17274
rect 11678 17054 11730 17106
rect 16830 17054 16882 17106
rect 23102 17054 23154 17106
rect 24334 17054 24386 17106
rect 25342 17054 25394 17106
rect 27246 17054 27298 17106
rect 27582 17054 27634 17106
rect 28814 17054 28866 17106
rect 30382 17054 30434 17106
rect 34526 17054 34578 17106
rect 39342 17054 39394 17106
rect 40238 17054 40290 17106
rect 41470 17054 41522 17106
rect 53342 17054 53394 17106
rect 54686 17054 54738 17106
rect 55470 17054 55522 17106
rect 56926 17054 56978 17106
rect 59950 17054 60002 17106
rect 71374 17054 71426 17106
rect 72606 17054 72658 17106
rect 4846 16942 4898 16994
rect 6862 16942 6914 16994
rect 16270 16942 16322 16994
rect 23326 16942 23378 16994
rect 24446 16942 24498 16994
rect 25790 16942 25842 16994
rect 28478 16942 28530 16994
rect 34750 16942 34802 16994
rect 39678 16942 39730 16994
rect 41022 16942 41074 16994
rect 42030 16942 42082 16994
rect 42478 16942 42530 16994
rect 43038 16942 43090 16994
rect 46062 16942 46114 16994
rect 47966 16942 48018 16994
rect 50766 16942 50818 16994
rect 55806 16942 55858 16994
rect 56814 16942 56866 16994
rect 57598 16942 57650 16994
rect 63086 16942 63138 16994
rect 67566 16942 67618 16994
rect 68910 16942 68962 16994
rect 69806 16942 69858 16994
rect 70478 16942 70530 16994
rect 71486 16942 71538 16994
rect 72270 16942 72322 16994
rect 77086 16942 77138 16994
rect 3950 16830 4002 16882
rect 6190 16830 6242 16882
rect 10334 16830 10386 16882
rect 10558 16830 10610 16882
rect 10894 16830 10946 16882
rect 11118 16830 11170 16882
rect 11342 16830 11394 16882
rect 11566 16830 11618 16882
rect 11902 16830 11954 16882
rect 15262 16830 15314 16882
rect 15598 16830 15650 16882
rect 16158 16830 16210 16882
rect 16382 16830 16434 16882
rect 17614 16830 17666 16882
rect 19182 16830 19234 16882
rect 19854 16830 19906 16882
rect 20414 16830 20466 16882
rect 23662 16830 23714 16882
rect 24110 16830 24162 16882
rect 26686 16830 26738 16882
rect 30606 16830 30658 16882
rect 32510 16830 32562 16882
rect 33070 16830 33122 16882
rect 33518 16830 33570 16882
rect 35646 16830 35698 16882
rect 37214 16830 37266 16882
rect 38558 16830 38610 16882
rect 41806 16830 41858 16882
rect 42366 16830 42418 16882
rect 42926 16830 42978 16882
rect 43598 16830 43650 16882
rect 44158 16830 44210 16882
rect 44942 16830 44994 16882
rect 46958 16830 47010 16882
rect 47406 16830 47458 16882
rect 48974 16830 49026 16882
rect 50094 16830 50146 16882
rect 54350 16830 54402 16882
rect 55134 16830 55186 16882
rect 55470 16830 55522 16882
rect 56590 16830 56642 16882
rect 57486 16830 57538 16882
rect 58494 16830 58546 16882
rect 59726 16830 59778 16882
rect 60174 16830 60226 16882
rect 63870 16830 63922 16882
rect 65550 16830 65602 16882
rect 65886 16830 65938 16882
rect 66446 16830 66498 16882
rect 66782 16830 66834 16882
rect 68350 16830 68402 16882
rect 69246 16830 69298 16882
rect 70702 16830 70754 16882
rect 71710 16830 71762 16882
rect 77870 16830 77922 16882
rect 8990 16718 9042 16770
rect 12350 16718 12402 16770
rect 14478 16718 14530 16770
rect 15710 16718 15762 16770
rect 18062 16718 18114 16770
rect 18846 16718 18898 16770
rect 28030 16718 28082 16770
rect 29934 16718 29986 16770
rect 32062 16718 32114 16770
rect 34414 16718 34466 16770
rect 35534 16718 35586 16770
rect 44382 16718 44434 16770
rect 46510 16718 46562 16770
rect 52894 16718 52946 16770
rect 60958 16718 61010 16770
rect 74958 16718 75010 16770
rect 1934 16606 1986 16658
rect 12014 16606 12066 16658
rect 19294 16606 19346 16658
rect 25566 16606 25618 16658
rect 25790 16606 25842 16658
rect 30830 16606 30882 16658
rect 32286 16606 32338 16658
rect 35422 16606 35474 16658
rect 39230 16606 39282 16658
rect 39678 16606 39730 16658
rect 10874 16438 10926 16490
rect 10978 16438 11030 16490
rect 11082 16438 11134 16490
rect 30194 16438 30246 16490
rect 30298 16438 30350 16490
rect 30402 16438 30454 16490
rect 49514 16438 49566 16490
rect 49618 16438 49670 16490
rect 49722 16438 49774 16490
rect 68834 16438 68886 16490
rect 68938 16438 68990 16490
rect 69042 16438 69094 16490
rect 7758 16270 7810 16322
rect 18734 16270 18786 16322
rect 32734 16270 32786 16322
rect 32958 16270 33010 16322
rect 33406 16270 33458 16322
rect 40238 16270 40290 16322
rect 67566 16270 67618 16322
rect 69134 16270 69186 16322
rect 9438 16158 9490 16210
rect 10334 16158 10386 16210
rect 12686 16158 12738 16210
rect 13582 16158 13634 16210
rect 14590 16158 14642 16210
rect 16158 16158 16210 16210
rect 16830 16158 16882 16210
rect 17502 16158 17554 16210
rect 22094 16158 22146 16210
rect 29374 16158 29426 16210
rect 34302 16158 34354 16210
rect 41134 16158 41186 16210
rect 41806 16158 41858 16210
rect 45838 16158 45890 16210
rect 46846 16158 46898 16210
rect 48190 16158 48242 16210
rect 51550 16158 51602 16210
rect 55918 16158 55970 16210
rect 58382 16158 58434 16210
rect 58942 16158 58994 16210
rect 59390 16158 59442 16210
rect 66222 16158 66274 16210
rect 69582 16158 69634 16210
rect 76414 16158 76466 16210
rect 3726 16046 3778 16098
rect 8094 16046 8146 16098
rect 8542 16046 8594 16098
rect 11118 16046 11170 16098
rect 15710 16046 15762 16098
rect 15934 16046 15986 16098
rect 17054 16046 17106 16098
rect 17838 16046 17890 16098
rect 18958 16046 19010 16098
rect 25006 16046 25058 16098
rect 26462 16046 26514 16098
rect 29934 16046 29986 16098
rect 31054 16046 31106 16098
rect 32510 16046 32562 16098
rect 35870 16046 35922 16098
rect 36990 16046 37042 16098
rect 38222 16046 38274 16098
rect 38894 16046 38946 16098
rect 39118 16046 39170 16098
rect 41246 16046 41298 16098
rect 42478 16046 42530 16098
rect 43038 16046 43090 16098
rect 43486 16046 43538 16098
rect 43822 16046 43874 16098
rect 44830 16046 44882 16098
rect 47630 16046 47682 16098
rect 48862 16046 48914 16098
rect 50990 16046 51042 16098
rect 53678 16046 53730 16098
rect 54014 16046 54066 16098
rect 54350 16046 54402 16098
rect 54686 16046 54738 16098
rect 57262 16046 57314 16098
rect 57934 16046 57986 16098
rect 68462 16046 68514 16098
rect 73838 16046 73890 16098
rect 74398 16046 74450 16098
rect 76974 16046 77026 16098
rect 3390 15934 3442 15986
rect 4398 15934 4450 15986
rect 8878 15934 8930 15986
rect 11342 15934 11394 15986
rect 11566 15934 11618 15986
rect 12238 15934 12290 15986
rect 14478 15934 14530 15986
rect 15262 15934 15314 15986
rect 16158 15934 16210 15986
rect 19854 15934 19906 15986
rect 24222 15934 24274 15986
rect 27022 15934 27074 15986
rect 27470 15934 27522 15986
rect 30270 15934 30322 15986
rect 31390 15934 31442 15986
rect 31726 15934 31778 15986
rect 32286 15934 32338 15986
rect 36430 15934 36482 15986
rect 42142 15934 42194 15986
rect 44046 15934 44098 15986
rect 49310 15934 49362 15986
rect 52222 15934 52274 15986
rect 56142 15934 56194 15986
rect 66558 15934 66610 15986
rect 4062 15822 4114 15874
rect 10446 15822 10498 15874
rect 14254 15822 14306 15874
rect 14702 15822 14754 15874
rect 14926 15822 14978 15874
rect 15150 15822 15202 15874
rect 16270 15822 16322 15874
rect 20190 15822 20242 15874
rect 20638 15822 20690 15874
rect 35982 15822 36034 15874
rect 42814 15822 42866 15874
rect 44158 15822 44210 15874
rect 46398 15822 46450 15874
rect 64990 15822 65042 15874
rect 65438 15822 65490 15874
rect 65662 15822 65714 15874
rect 74174 15822 74226 15874
rect 76750 15822 76802 15874
rect 20534 15654 20586 15706
rect 20638 15654 20690 15706
rect 20742 15654 20794 15706
rect 39854 15654 39906 15706
rect 39958 15654 40010 15706
rect 40062 15654 40114 15706
rect 59174 15654 59226 15706
rect 59278 15654 59330 15706
rect 59382 15654 59434 15706
rect 78494 15654 78546 15706
rect 78598 15654 78650 15706
rect 78702 15654 78754 15706
rect 5294 15486 5346 15538
rect 7646 15486 7698 15538
rect 21758 15486 21810 15538
rect 22206 15486 22258 15538
rect 23438 15486 23490 15538
rect 26686 15486 26738 15538
rect 30830 15486 30882 15538
rect 31278 15486 31330 15538
rect 32286 15486 32338 15538
rect 32958 15486 33010 15538
rect 33854 15486 33906 15538
rect 34526 15486 34578 15538
rect 34862 15486 34914 15538
rect 35198 15486 35250 15538
rect 39230 15486 39282 15538
rect 43486 15486 43538 15538
rect 43598 15486 43650 15538
rect 44158 15486 44210 15538
rect 44382 15486 44434 15538
rect 46062 15486 46114 15538
rect 48862 15486 48914 15538
rect 49086 15486 49138 15538
rect 50990 15486 51042 15538
rect 52558 15486 52610 15538
rect 54798 15486 54850 15538
rect 55134 15486 55186 15538
rect 56590 15486 56642 15538
rect 56926 15486 56978 15538
rect 57262 15486 57314 15538
rect 58046 15486 58098 15538
rect 63870 15486 63922 15538
rect 67566 15486 67618 15538
rect 68238 15486 68290 15538
rect 68686 15486 68738 15538
rect 69134 15486 69186 15538
rect 2718 15374 2770 15426
rect 5966 15374 6018 15426
rect 6414 15374 6466 15426
rect 6862 15374 6914 15426
rect 16158 15374 16210 15426
rect 17390 15374 17442 15426
rect 24446 15374 24498 15426
rect 29710 15374 29762 15426
rect 32062 15374 32114 15426
rect 32510 15374 32562 15426
rect 33182 15374 33234 15426
rect 33630 15374 33682 15426
rect 34078 15374 34130 15426
rect 36766 15374 36818 15426
rect 42702 15374 42754 15426
rect 50094 15374 50146 15426
rect 55470 15374 55522 15426
rect 57598 15374 57650 15426
rect 59278 15374 59330 15426
rect 64654 15374 64706 15426
rect 65214 15374 65266 15426
rect 65550 15374 65602 15426
rect 66782 15374 66834 15426
rect 70030 15374 70082 15426
rect 74510 15374 74562 15426
rect 2046 15262 2098 15314
rect 5630 15262 5682 15314
rect 7198 15262 7250 15314
rect 11566 15262 11618 15314
rect 12798 15262 12850 15314
rect 13134 15262 13186 15314
rect 14590 15262 14642 15314
rect 17614 15262 17666 15314
rect 17950 15262 18002 15314
rect 18286 15262 18338 15314
rect 18622 15262 18674 15314
rect 21534 15262 21586 15314
rect 23662 15262 23714 15314
rect 24110 15262 24162 15314
rect 24558 15262 24610 15314
rect 25342 15262 25394 15314
rect 25566 15262 25618 15314
rect 25790 15262 25842 15314
rect 26350 15262 26402 15314
rect 26462 15262 26514 15314
rect 28142 15262 28194 15314
rect 29598 15262 29650 15314
rect 31726 15262 31778 15314
rect 33294 15262 33346 15314
rect 35758 15262 35810 15314
rect 36654 15262 36706 15314
rect 37438 15262 37490 15314
rect 40014 15262 40066 15314
rect 40238 15262 40290 15314
rect 40910 15262 40962 15314
rect 41134 15262 41186 15314
rect 43710 15262 43762 15314
rect 44046 15262 44098 15314
rect 44718 15262 44770 15314
rect 47742 15262 47794 15314
rect 48750 15262 48802 15314
rect 49646 15262 49698 15314
rect 51438 15262 51490 15314
rect 56030 15262 56082 15314
rect 59726 15262 59778 15314
rect 60286 15262 60338 15314
rect 64766 15262 64818 15314
rect 66334 15262 66386 15314
rect 67230 15262 67282 15314
rect 69806 15262 69858 15314
rect 73950 15262 74002 15314
rect 74398 15262 74450 15314
rect 76078 15262 76130 15314
rect 4846 15150 4898 15202
rect 14702 15150 14754 15202
rect 16606 15150 16658 15202
rect 18398 15150 18450 15202
rect 19182 15150 19234 15202
rect 23550 15150 23602 15202
rect 27134 15150 27186 15202
rect 27582 15150 27634 15202
rect 35534 15150 35586 15202
rect 36766 15150 36818 15202
rect 38222 15150 38274 15202
rect 40350 15150 40402 15202
rect 45166 15150 45218 15202
rect 45614 15150 45666 15202
rect 48190 15150 48242 15202
rect 51774 15150 51826 15202
rect 53006 15150 53058 15202
rect 59614 15150 59666 15202
rect 66894 15150 66946 15202
rect 73166 15150 73218 15202
rect 77982 15150 78034 15202
rect 15038 15038 15090 15090
rect 15934 15038 15986 15090
rect 16494 15038 16546 15090
rect 17726 15038 17778 15090
rect 26014 15038 26066 15090
rect 28590 15038 28642 15090
rect 32174 15038 32226 15090
rect 33742 15038 33794 15090
rect 36094 15038 36146 15090
rect 73614 15038 73666 15090
rect 10874 14870 10926 14922
rect 10978 14870 11030 14922
rect 11082 14870 11134 14922
rect 30194 14870 30246 14922
rect 30298 14870 30350 14922
rect 30402 14870 30454 14922
rect 49514 14870 49566 14922
rect 49618 14870 49670 14922
rect 49722 14870 49774 14922
rect 68834 14870 68886 14922
rect 68938 14870 68990 14922
rect 69042 14870 69094 14922
rect 26910 14702 26962 14754
rect 27358 14702 27410 14754
rect 38558 14702 38610 14754
rect 57262 14702 57314 14754
rect 1934 14590 1986 14642
rect 13918 14590 13970 14642
rect 17166 14590 17218 14642
rect 18286 14590 18338 14642
rect 22094 14590 22146 14642
rect 26910 14590 26962 14642
rect 32734 14590 32786 14642
rect 37662 14590 37714 14642
rect 37998 14590 38050 14642
rect 40910 14590 40962 14642
rect 42030 14590 42082 14642
rect 49198 14590 49250 14642
rect 51662 14590 51714 14642
rect 54350 14590 54402 14642
rect 56142 14590 56194 14642
rect 59278 14590 59330 14642
rect 64430 14590 64482 14642
rect 65998 14590 66050 14642
rect 68910 14590 68962 14642
rect 71038 14590 71090 14642
rect 4286 14478 4338 14530
rect 6078 14478 6130 14530
rect 6862 14478 6914 14530
rect 14702 14478 14754 14530
rect 16718 14478 16770 14530
rect 17390 14478 17442 14530
rect 18398 14478 18450 14530
rect 18622 14478 18674 14530
rect 18958 14478 19010 14530
rect 21534 14478 21586 14530
rect 27918 14478 27970 14530
rect 28590 14478 28642 14530
rect 29150 14478 29202 14530
rect 29710 14478 29762 14530
rect 30270 14478 30322 14530
rect 31278 14478 31330 14530
rect 32398 14478 32450 14530
rect 33630 14478 33682 14530
rect 34638 14478 34690 14530
rect 35646 14478 35698 14530
rect 36206 14478 36258 14530
rect 37438 14478 37490 14530
rect 38334 14478 38386 14530
rect 39678 14478 39730 14530
rect 39902 14478 39954 14530
rect 41022 14478 41074 14530
rect 46958 14478 47010 14530
rect 48302 14478 48354 14530
rect 50318 14478 50370 14530
rect 51102 14478 51154 14530
rect 52110 14478 52162 14530
rect 52894 14478 52946 14530
rect 54686 14478 54738 14530
rect 55246 14478 55298 14530
rect 56590 14478 56642 14530
rect 56702 14478 56754 14530
rect 57038 14478 57090 14530
rect 57374 14478 57426 14530
rect 57934 14478 57986 14530
rect 58830 14478 58882 14530
rect 59614 14478 59666 14530
rect 63982 14478 64034 14530
rect 64094 14478 64146 14530
rect 64542 14478 64594 14530
rect 66110 14478 66162 14530
rect 66894 14478 66946 14530
rect 71822 14478 71874 14530
rect 75630 14478 75682 14530
rect 76190 14478 76242 14530
rect 6750 14366 6802 14418
rect 7870 14366 7922 14418
rect 18846 14366 18898 14418
rect 41582 14366 41634 14418
rect 47518 14366 47570 14418
rect 50766 14366 50818 14418
rect 53790 14366 53842 14418
rect 56926 14366 56978 14418
rect 57598 14366 57650 14418
rect 59838 14366 59890 14418
rect 65886 14366 65938 14418
rect 76862 14366 76914 14418
rect 77198 14366 77250 14418
rect 77646 14366 77698 14418
rect 4846 14254 4898 14306
rect 5742 14254 5794 14306
rect 7534 14254 7586 14306
rect 12350 14254 12402 14306
rect 15150 14254 15202 14306
rect 16942 14254 16994 14306
rect 17166 14254 17218 14306
rect 17950 14254 18002 14306
rect 18174 14254 18226 14306
rect 21310 14254 21362 14306
rect 27582 14254 27634 14306
rect 38894 14254 38946 14306
rect 39790 14254 39842 14306
rect 42590 14254 42642 14306
rect 55582 14254 55634 14306
rect 59278 14254 59330 14306
rect 59390 14254 59442 14306
rect 63534 14254 63586 14306
rect 64318 14254 64370 14306
rect 72270 14254 72322 14306
rect 74622 14254 74674 14306
rect 76526 14254 76578 14306
rect 20534 14086 20586 14138
rect 20638 14086 20690 14138
rect 20742 14086 20794 14138
rect 39854 14086 39906 14138
rect 39958 14086 40010 14138
rect 40062 14086 40114 14138
rect 59174 14086 59226 14138
rect 59278 14086 59330 14138
rect 59382 14086 59434 14138
rect 78494 14086 78546 14138
rect 78598 14086 78650 14138
rect 78702 14086 78754 14138
rect 11902 13918 11954 13970
rect 13022 13918 13074 13970
rect 16494 13918 16546 13970
rect 17838 13918 17890 13970
rect 24334 13918 24386 13970
rect 25454 13918 25506 13970
rect 30046 13918 30098 13970
rect 33406 13918 33458 13970
rect 34190 13918 34242 13970
rect 34862 13918 34914 13970
rect 37550 13918 37602 13970
rect 39230 13918 39282 13970
rect 43038 13918 43090 13970
rect 46398 13918 46450 13970
rect 47854 13918 47906 13970
rect 47966 13918 48018 13970
rect 52894 13918 52946 13970
rect 55582 13918 55634 13970
rect 56142 13918 56194 13970
rect 59726 13918 59778 13970
rect 63310 13918 63362 13970
rect 63534 13918 63586 13970
rect 63646 13918 63698 13970
rect 66110 13918 66162 13970
rect 70030 13918 70082 13970
rect 8430 13806 8482 13858
rect 10334 13806 10386 13858
rect 10558 13806 10610 13858
rect 13918 13806 13970 13858
rect 14030 13806 14082 13858
rect 15934 13806 15986 13858
rect 23102 13806 23154 13858
rect 23998 13806 24050 13858
rect 28366 13806 28418 13858
rect 30494 13806 30546 13858
rect 31838 13806 31890 13858
rect 33070 13806 33122 13858
rect 33966 13806 34018 13858
rect 34414 13806 34466 13858
rect 35646 13806 35698 13858
rect 37886 13806 37938 13858
rect 40910 13806 40962 13858
rect 41246 13806 41298 13858
rect 41694 13806 41746 13858
rect 43262 13806 43314 13858
rect 43598 13806 43650 13858
rect 45166 13806 45218 13858
rect 46734 13806 46786 13858
rect 50430 13806 50482 13858
rect 54462 13806 54514 13858
rect 60734 13806 60786 13858
rect 61966 13806 62018 13858
rect 62862 13806 62914 13858
rect 63870 13806 63922 13858
rect 65438 13806 65490 13858
rect 66222 13806 66274 13858
rect 70590 13806 70642 13858
rect 71150 13806 71202 13858
rect 73278 13806 73330 13858
rect 74062 13806 74114 13858
rect 74398 13806 74450 13858
rect 76862 13806 76914 13858
rect 2158 13694 2210 13746
rect 8766 13694 8818 13746
rect 9662 13694 9714 13746
rect 9998 13694 10050 13746
rect 11678 13694 11730 13746
rect 12126 13694 12178 13746
rect 12350 13694 12402 13746
rect 12686 13694 12738 13746
rect 15822 13694 15874 13746
rect 16046 13694 16098 13746
rect 17390 13694 17442 13746
rect 17614 13694 17666 13746
rect 17726 13694 17778 13746
rect 17950 13694 18002 13746
rect 22766 13694 22818 13746
rect 22990 13694 23042 13746
rect 27134 13694 27186 13746
rect 28254 13694 28306 13746
rect 28478 13694 28530 13746
rect 29038 13694 29090 13746
rect 31502 13694 31554 13746
rect 32062 13694 32114 13746
rect 33294 13694 33346 13746
rect 33630 13694 33682 13746
rect 38110 13694 38162 13746
rect 42590 13694 42642 13746
rect 42814 13694 42866 13746
rect 42926 13694 42978 13746
rect 43822 13694 43874 13746
rect 44046 13694 44098 13746
rect 45390 13694 45442 13746
rect 47294 13694 47346 13746
rect 47630 13694 47682 13746
rect 49086 13694 49138 13746
rect 50206 13694 50258 13746
rect 51662 13694 51714 13746
rect 53342 13694 53394 13746
rect 54910 13694 54962 13746
rect 55246 13694 55298 13746
rect 56702 13694 56754 13746
rect 58046 13694 58098 13746
rect 58382 13694 58434 13746
rect 58830 13694 58882 13746
rect 61294 13694 61346 13746
rect 62190 13694 62242 13746
rect 63422 13694 63474 13746
rect 64430 13694 64482 13746
rect 66894 13694 66946 13746
rect 67902 13694 67954 13746
rect 68238 13694 68290 13746
rect 70366 13694 70418 13746
rect 71710 13694 71762 13746
rect 72718 13694 72770 13746
rect 73390 13694 73442 13746
rect 77646 13694 77698 13746
rect 2942 13582 2994 13634
rect 5070 13582 5122 13634
rect 7198 13582 7250 13634
rect 11342 13582 11394 13634
rect 12910 13582 12962 13634
rect 21086 13582 21138 13634
rect 25342 13582 25394 13634
rect 26014 13582 26066 13634
rect 26686 13582 26738 13634
rect 27806 13582 27858 13634
rect 29486 13582 29538 13634
rect 34078 13582 34130 13634
rect 36094 13582 36146 13634
rect 36654 13582 36706 13634
rect 37102 13582 37154 13634
rect 38446 13582 38498 13634
rect 40014 13582 40066 13634
rect 42142 13582 42194 13634
rect 43934 13582 43986 13634
rect 45950 13582 46002 13634
rect 49870 13582 49922 13634
rect 74734 13582 74786 13634
rect 13918 13470 13970 13522
rect 23550 13470 23602 13522
rect 26910 13470 26962 13522
rect 27582 13470 27634 13522
rect 30718 13470 30770 13522
rect 40126 13470 40178 13522
rect 52446 13470 52498 13522
rect 72382 13470 72434 13522
rect 10874 13302 10926 13354
rect 10978 13302 11030 13354
rect 11082 13302 11134 13354
rect 30194 13302 30246 13354
rect 30298 13302 30350 13354
rect 30402 13302 30454 13354
rect 49514 13302 49566 13354
rect 49618 13302 49670 13354
rect 49722 13302 49774 13354
rect 68834 13302 68886 13354
rect 68938 13302 68990 13354
rect 69042 13302 69094 13354
rect 18622 13134 18674 13186
rect 31278 13134 31330 13186
rect 31838 13134 31890 13186
rect 33070 13134 33122 13186
rect 45390 13134 45442 13186
rect 45726 13134 45778 13186
rect 55470 13134 55522 13186
rect 56254 13134 56306 13186
rect 74510 13134 74562 13186
rect 8094 13022 8146 13074
rect 10222 13022 10274 13074
rect 16942 13022 16994 13074
rect 20078 13022 20130 13074
rect 20414 13022 20466 13074
rect 24222 13022 24274 13074
rect 25118 13022 25170 13074
rect 27582 13022 27634 13074
rect 29262 13022 29314 13074
rect 32734 13022 32786 13074
rect 37214 13022 37266 13074
rect 39118 13022 39170 13074
rect 41918 13022 41970 13074
rect 42254 13022 42306 13074
rect 44270 13022 44322 13074
rect 44942 13022 44994 13074
rect 50206 13022 50258 13074
rect 55806 13022 55858 13074
rect 56254 13022 56306 13074
rect 57038 13022 57090 13074
rect 58494 13022 58546 13074
rect 59726 13022 59778 13074
rect 61630 13022 61682 13074
rect 63758 13022 63810 13074
rect 64206 13022 64258 13074
rect 65326 13022 65378 13074
rect 72606 13022 72658 13074
rect 2718 12910 2770 12962
rect 3614 12910 3666 12962
rect 7422 12910 7474 12962
rect 14590 12910 14642 12962
rect 15934 12910 15986 12962
rect 16270 12910 16322 12962
rect 16382 12910 16434 12962
rect 17502 12910 17554 12962
rect 18286 12910 18338 12962
rect 19518 12910 19570 12962
rect 20526 12910 20578 12962
rect 20862 12910 20914 12962
rect 21534 12910 21586 12962
rect 22990 12910 23042 12962
rect 24446 12910 24498 12962
rect 24894 12910 24946 12962
rect 25230 12910 25282 12962
rect 26126 12910 26178 12962
rect 26462 12910 26514 12962
rect 26686 12910 26738 12962
rect 27918 12910 27970 12962
rect 28702 12910 28754 12962
rect 32286 12910 32338 12962
rect 32846 12910 32898 12962
rect 33294 12910 33346 12962
rect 33742 12910 33794 12962
rect 34638 12910 34690 12962
rect 34974 12910 35026 12962
rect 35198 12910 35250 12962
rect 35310 12910 35362 12962
rect 35422 12910 35474 12962
rect 37662 12910 37714 12962
rect 39678 12910 39730 12962
rect 40350 12910 40402 12962
rect 41470 12910 41522 12962
rect 42366 12910 42418 12962
rect 46398 12910 46450 12962
rect 47070 12910 47122 12962
rect 48302 12910 48354 12962
rect 48638 12910 48690 12962
rect 48974 12910 49026 12962
rect 51550 12910 51602 12962
rect 55358 12910 55410 12962
rect 56702 12910 56754 12962
rect 56814 12910 56866 12962
rect 57150 12910 57202 12962
rect 57822 12910 57874 12962
rect 59278 12910 59330 12962
rect 60846 12910 60898 12962
rect 65550 12910 65602 12962
rect 66222 12910 66274 12962
rect 66670 12910 66722 12962
rect 69694 12910 69746 12962
rect 73166 12910 73218 12962
rect 73950 12910 74002 12962
rect 2382 12798 2434 12850
rect 3278 12798 3330 12850
rect 6526 12798 6578 12850
rect 11790 12798 11842 12850
rect 12798 12798 12850 12850
rect 13806 12798 13858 12850
rect 14030 12798 14082 12850
rect 17278 12798 17330 12850
rect 17726 12798 17778 12850
rect 17838 12798 17890 12850
rect 18062 12798 18114 12850
rect 18846 12798 18898 12850
rect 18958 12798 19010 12850
rect 20302 12798 20354 12850
rect 21758 12798 21810 12850
rect 24222 12798 24274 12850
rect 24670 12798 24722 12850
rect 27246 12798 27298 12850
rect 31390 12798 31442 12850
rect 31726 12798 31778 12850
rect 34526 12798 34578 12850
rect 46286 12798 46338 12850
rect 50878 12798 50930 12850
rect 57038 12798 57090 12850
rect 57934 12798 57986 12850
rect 64878 12798 64930 12850
rect 66894 12798 66946 12850
rect 70366 12798 70418 12850
rect 72942 12798 72994 12850
rect 73726 12798 73778 12850
rect 74846 12798 74898 12850
rect 75294 12798 75346 12850
rect 6190 12686 6242 12738
rect 11902 12686 11954 12738
rect 12910 12686 12962 12738
rect 14254 12686 14306 12738
rect 15038 12686 15090 12738
rect 15486 12686 15538 12738
rect 16046 12686 16098 12738
rect 16158 12686 16210 12738
rect 18510 12686 18562 12738
rect 19182 12686 19234 12738
rect 21198 12686 21250 12738
rect 21310 12686 21362 12738
rect 23774 12686 23826 12738
rect 24110 12686 24162 12738
rect 25454 12686 25506 12738
rect 26910 12686 26962 12738
rect 27022 12686 27074 12738
rect 32398 12686 32450 12738
rect 32622 12686 32674 12738
rect 35534 12686 35586 12738
rect 36094 12686 36146 12738
rect 36430 12686 36482 12738
rect 37438 12686 37490 12738
rect 59054 12686 59106 12738
rect 64654 12686 64706 12738
rect 73278 12686 73330 12738
rect 75630 12686 75682 12738
rect 20534 12518 20586 12570
rect 20638 12518 20690 12570
rect 20742 12518 20794 12570
rect 39854 12518 39906 12570
rect 39958 12518 40010 12570
rect 40062 12518 40114 12570
rect 59174 12518 59226 12570
rect 59278 12518 59330 12570
rect 59382 12518 59434 12570
rect 78494 12518 78546 12570
rect 78598 12518 78650 12570
rect 78702 12518 78754 12570
rect 23214 12350 23266 12402
rect 25230 12350 25282 12402
rect 32062 12350 32114 12402
rect 33518 12350 33570 12402
rect 33630 12350 33682 12402
rect 33854 12350 33906 12402
rect 34526 12350 34578 12402
rect 38670 12350 38722 12402
rect 39454 12350 39506 12402
rect 41470 12350 41522 12402
rect 41694 12350 41746 12402
rect 42366 12350 42418 12402
rect 43598 12350 43650 12402
rect 47854 12350 47906 12402
rect 53566 12350 53618 12402
rect 55806 12350 55858 12402
rect 56814 12350 56866 12402
rect 57374 12350 57426 12402
rect 58158 12350 58210 12402
rect 58382 12350 58434 12402
rect 60174 12350 60226 12402
rect 60398 12350 60450 12402
rect 61070 12350 61122 12402
rect 61742 12350 61794 12402
rect 64542 12350 64594 12402
rect 65102 12350 65154 12402
rect 65662 12350 65714 12402
rect 65886 12350 65938 12402
rect 69806 12350 69858 12402
rect 70478 12350 70530 12402
rect 2830 12238 2882 12290
rect 6302 12238 6354 12290
rect 17614 12238 17666 12290
rect 18958 12238 19010 12290
rect 20638 12238 20690 12290
rect 20974 12238 21026 12290
rect 22430 12238 22482 12290
rect 23998 12238 24050 12290
rect 26798 12238 26850 12290
rect 28142 12238 28194 12290
rect 28702 12238 28754 12290
rect 33294 12238 33346 12290
rect 39006 12238 39058 12290
rect 40126 12238 40178 12290
rect 41246 12238 41298 12290
rect 41806 12238 41858 12290
rect 45166 12238 45218 12290
rect 53454 12238 53506 12290
rect 54238 12238 54290 12290
rect 59390 12238 59442 12290
rect 62414 12238 62466 12290
rect 62862 12238 62914 12290
rect 66558 12238 66610 12290
rect 70814 12238 70866 12290
rect 77086 12238 77138 12290
rect 3166 12126 3218 12178
rect 5518 12126 5570 12178
rect 12350 12126 12402 12178
rect 12686 12126 12738 12178
rect 14254 12126 14306 12178
rect 15710 12126 15762 12178
rect 18622 12126 18674 12178
rect 18846 12126 18898 12178
rect 19406 12126 19458 12178
rect 19854 12126 19906 12178
rect 20414 12126 20466 12178
rect 22878 12126 22930 12178
rect 24222 12126 24274 12178
rect 24334 12126 24386 12178
rect 24446 12126 24498 12178
rect 24670 12126 24722 12178
rect 25678 12126 25730 12178
rect 25790 12126 25842 12178
rect 26014 12126 26066 12178
rect 27022 12126 27074 12178
rect 27918 12126 27970 12178
rect 28926 12126 28978 12178
rect 33742 12126 33794 12178
rect 36206 12126 36258 12178
rect 38110 12126 38162 12178
rect 39902 12126 39954 12178
rect 42478 12126 42530 12178
rect 42814 12126 42866 12178
rect 43038 12126 43090 12178
rect 43486 12126 43538 12178
rect 44494 12126 44546 12178
rect 50654 12126 50706 12178
rect 51774 12126 51826 12178
rect 52334 12126 52386 12178
rect 54910 12126 54962 12178
rect 57934 12126 57986 12178
rect 58046 12126 58098 12178
rect 58270 12126 58322 12178
rect 59054 12126 59106 12178
rect 60398 12126 60450 12178
rect 62078 12126 62130 12178
rect 63422 12126 63474 12178
rect 63870 12126 63922 12178
rect 65550 12126 65602 12178
rect 66894 12126 66946 12178
rect 70142 12126 70194 12178
rect 77758 12126 77810 12178
rect 8430 12014 8482 12066
rect 12126 12014 12178 12066
rect 15822 12014 15874 12066
rect 21310 12014 21362 12066
rect 22206 12014 22258 12066
rect 23662 12014 23714 12066
rect 27694 12014 27746 12066
rect 32510 12014 32562 12066
rect 35422 12014 35474 12066
rect 36990 12014 37042 12066
rect 39342 12014 39394 12066
rect 41806 12014 41858 12066
rect 43150 12014 43202 12066
rect 43934 12014 43986 12066
rect 47294 12014 47346 12066
rect 50094 12014 50146 12066
rect 74958 12014 75010 12066
rect 16270 11902 16322 11954
rect 20078 11902 20130 11954
rect 20526 11902 20578 11954
rect 29262 11902 29314 11954
rect 31950 11902 32002 11954
rect 32622 11902 32674 11954
rect 10874 11734 10926 11786
rect 10978 11734 11030 11786
rect 11082 11734 11134 11786
rect 30194 11734 30246 11786
rect 30298 11734 30350 11786
rect 30402 11734 30454 11786
rect 49514 11734 49566 11786
rect 49618 11734 49670 11786
rect 49722 11734 49774 11786
rect 68834 11734 68886 11786
rect 68938 11734 68990 11786
rect 69042 11734 69094 11786
rect 6638 11566 6690 11618
rect 18398 11566 18450 11618
rect 19182 11566 19234 11618
rect 19294 11566 19346 11618
rect 19518 11566 19570 11618
rect 21758 11566 21810 11618
rect 48190 11566 48242 11618
rect 2494 11454 2546 11506
rect 4622 11454 4674 11506
rect 5070 11454 5122 11506
rect 6974 11454 7026 11506
rect 8318 11454 8370 11506
rect 16494 11454 16546 11506
rect 17278 11454 17330 11506
rect 18286 11454 18338 11506
rect 21310 11454 21362 11506
rect 22206 11454 22258 11506
rect 26798 11454 26850 11506
rect 27246 11454 27298 11506
rect 27470 11454 27522 11506
rect 31950 11454 32002 11506
rect 34190 11454 34242 11506
rect 35982 11454 36034 11506
rect 39006 11454 39058 11506
rect 40014 11454 40066 11506
rect 40350 11454 40402 11506
rect 40798 11454 40850 11506
rect 42142 11454 42194 11506
rect 42366 11454 42418 11506
rect 43598 11454 43650 11506
rect 46734 11454 46786 11506
rect 50206 11454 50258 11506
rect 56030 11454 56082 11506
rect 57374 11454 57426 11506
rect 60734 11454 60786 11506
rect 61518 11454 61570 11506
rect 67790 11454 67842 11506
rect 1822 11342 1874 11394
rect 7758 11342 7810 11394
rect 14590 11342 14642 11394
rect 15262 11342 15314 11394
rect 15934 11342 15986 11394
rect 16718 11342 16770 11394
rect 16830 11342 16882 11394
rect 21534 11342 21586 11394
rect 22766 11342 22818 11394
rect 23214 11342 23266 11394
rect 23550 11342 23602 11394
rect 23774 11342 23826 11394
rect 24446 11342 24498 11394
rect 25342 11342 25394 11394
rect 25566 11342 25618 11394
rect 25678 11342 25730 11394
rect 27134 11342 27186 11394
rect 27694 11342 27746 11394
rect 28030 11342 28082 11394
rect 28142 11342 28194 11394
rect 28366 11342 28418 11394
rect 29262 11342 29314 11394
rect 30718 11342 30770 11394
rect 31166 11342 31218 11394
rect 31838 11342 31890 11394
rect 38222 11342 38274 11394
rect 41694 11342 41746 11394
rect 43374 11342 43426 11394
rect 43822 11342 43874 11394
rect 44046 11342 44098 11394
rect 44942 11342 44994 11394
rect 49758 11342 49810 11394
rect 53118 11342 53170 11394
rect 53902 11342 53954 11394
rect 55022 11342 55074 11394
rect 57710 11342 57762 11394
rect 58382 11342 58434 11394
rect 58718 11342 58770 11394
rect 59390 11342 59442 11394
rect 64990 11342 65042 11394
rect 75630 11342 75682 11394
rect 7534 11230 7586 11282
rect 12014 11230 12066 11282
rect 12798 11230 12850 11282
rect 13806 11230 13858 11282
rect 14030 11230 14082 11282
rect 15486 11230 15538 11282
rect 16158 11230 16210 11282
rect 18622 11230 18674 11282
rect 22542 11230 22594 11282
rect 24110 11230 24162 11282
rect 24558 11230 24610 11282
rect 25118 11230 25170 11282
rect 37998 11230 38050 11282
rect 41806 11230 41858 11282
rect 48526 11230 48578 11282
rect 48862 11230 48914 11282
rect 52110 11230 52162 11282
rect 52782 11230 52834 11282
rect 53790 11230 53842 11282
rect 59502 11230 59554 11282
rect 65662 11230 65714 11282
rect 72494 11230 72546 11282
rect 72606 11230 72658 11282
rect 76750 11230 76802 11282
rect 77086 11230 77138 11282
rect 8766 11118 8818 11170
rect 11230 11118 11282 11170
rect 11790 11118 11842 11170
rect 12126 11118 12178 11170
rect 12910 11118 12962 11170
rect 14254 11118 14306 11170
rect 15374 11118 15426 11170
rect 16382 11118 16434 11170
rect 19966 11118 20018 11170
rect 22878 11118 22930 11170
rect 22990 11118 23042 11170
rect 23998 11118 24050 11170
rect 24670 11118 24722 11170
rect 25454 11118 25506 11170
rect 26350 11118 26402 11170
rect 29710 11118 29762 11170
rect 30158 11118 30210 11170
rect 30494 11118 30546 11170
rect 30606 11118 30658 11170
rect 33182 11118 33234 11170
rect 36430 11118 36482 11170
rect 36990 11118 37042 11170
rect 37326 11118 37378 11170
rect 39454 11118 39506 11170
rect 41246 11118 41298 11170
rect 41358 11118 41410 11170
rect 41918 11118 41970 11170
rect 42814 11118 42866 11170
rect 43598 11118 43650 11170
rect 47854 11118 47906 11170
rect 49422 11118 49474 11170
rect 51774 11118 51826 11170
rect 54462 11118 54514 11170
rect 54798 11118 54850 11170
rect 56814 11118 56866 11170
rect 57934 11118 57986 11170
rect 61070 11118 61122 11170
rect 72270 11118 72322 11170
rect 72830 11118 72882 11170
rect 74622 11118 74674 11170
rect 76414 11118 76466 11170
rect 20534 10950 20586 11002
rect 20638 10950 20690 11002
rect 20742 10950 20794 11002
rect 39854 10950 39906 11002
rect 39958 10950 40010 11002
rect 40062 10950 40114 11002
rect 59174 10950 59226 11002
rect 59278 10950 59330 11002
rect 59382 10950 59434 11002
rect 78494 10950 78546 11002
rect 78598 10950 78650 11002
rect 78702 10950 78754 11002
rect 4734 10782 4786 10834
rect 17278 10782 17330 10834
rect 18062 10782 18114 10834
rect 20190 10782 20242 10834
rect 20974 10782 21026 10834
rect 21198 10782 21250 10834
rect 23214 10782 23266 10834
rect 24670 10782 24722 10834
rect 25454 10782 25506 10834
rect 26126 10782 26178 10834
rect 27806 10782 27858 10834
rect 37886 10782 37938 10834
rect 38222 10782 38274 10834
rect 41694 10782 41746 10834
rect 42702 10782 42754 10834
rect 46398 10782 46450 10834
rect 54350 10782 54402 10834
rect 54798 10782 54850 10834
rect 56702 10782 56754 10834
rect 66446 10782 66498 10834
rect 67230 10782 67282 10834
rect 68126 10782 68178 10834
rect 76526 10782 76578 10834
rect 5854 10670 5906 10722
rect 8878 10670 8930 10722
rect 9550 10670 9602 10722
rect 17502 10670 17554 10722
rect 19966 10670 20018 10722
rect 20414 10670 20466 10722
rect 22654 10670 22706 10722
rect 30382 10670 30434 10722
rect 33966 10670 34018 10722
rect 39678 10670 39730 10722
rect 40014 10670 40066 10722
rect 41918 10670 41970 10722
rect 4286 10558 4338 10610
rect 5630 10558 5682 10610
rect 8654 10558 8706 10610
rect 10110 10558 10162 10610
rect 12350 10558 12402 10610
rect 12574 10558 12626 10610
rect 14254 10558 14306 10610
rect 15486 10558 15538 10610
rect 17614 10558 17666 10610
rect 20526 10558 20578 10610
rect 20862 10558 20914 10610
rect 22206 10558 22258 10610
rect 23886 10558 23938 10610
rect 24110 10558 24162 10610
rect 24222 10614 24274 10666
rect 47854 10670 47906 10722
rect 48190 10670 48242 10722
rect 51662 10670 51714 10722
rect 55918 10670 55970 10722
rect 61742 10670 61794 10722
rect 64990 10670 65042 10722
rect 65438 10670 65490 10722
rect 69358 10670 69410 10722
rect 69582 10670 69634 10722
rect 76750 10670 76802 10722
rect 77422 10670 77474 10722
rect 28590 10558 28642 10610
rect 29710 10558 29762 10610
rect 34302 10558 34354 10610
rect 42254 10558 42306 10610
rect 43150 10558 43202 10610
rect 43374 10558 43426 10610
rect 43598 10558 43650 10610
rect 43822 10558 43874 10610
rect 50878 10558 50930 10610
rect 55806 10558 55858 10610
rect 57934 10558 57986 10610
rect 61966 10558 62018 10610
rect 65998 10558 66050 10610
rect 66782 10558 66834 10610
rect 69134 10558 69186 10610
rect 72606 10558 72658 10610
rect 76974 10558 77026 10610
rect 77646 10558 77698 10610
rect 1934 10446 1986 10498
rect 6414 10446 6466 10498
rect 6974 10446 7026 10498
rect 10558 10446 10610 10498
rect 15710 10446 15762 10498
rect 18510 10446 18562 10498
rect 21758 10446 21810 10498
rect 23662 10446 23714 10498
rect 27694 10446 27746 10498
rect 32510 10446 32562 10498
rect 38670 10446 38722 10498
rect 41134 10446 41186 10498
rect 43486 10446 43538 10498
rect 44270 10446 44322 10498
rect 53790 10446 53842 10498
rect 58606 10446 58658 10498
rect 60734 10446 60786 10498
rect 63870 10446 63922 10498
rect 65662 10446 65714 10498
rect 68574 10446 68626 10498
rect 69246 10446 69298 10498
rect 73390 10446 73442 10498
rect 75518 10446 75570 10498
rect 76078 10446 76130 10498
rect 5070 10334 5122 10386
rect 16046 10334 16098 10386
rect 39118 10334 39170 10386
rect 39454 10334 39506 10386
rect 41134 10334 41186 10386
rect 41470 10334 41522 10386
rect 41582 10334 41634 10386
rect 55134 10334 55186 10386
rect 75742 10334 75794 10386
rect 76526 10334 76578 10386
rect 10874 10166 10926 10218
rect 10978 10166 11030 10218
rect 11082 10166 11134 10218
rect 30194 10166 30246 10218
rect 30298 10166 30350 10218
rect 30402 10166 30454 10218
rect 49514 10166 49566 10218
rect 49618 10166 49670 10218
rect 49722 10166 49774 10218
rect 68834 10166 68886 10218
rect 68938 10166 68990 10218
rect 69042 10166 69094 10218
rect 16830 9998 16882 10050
rect 17390 9998 17442 10050
rect 17950 9998 18002 10050
rect 21310 9998 21362 10050
rect 45278 9998 45330 10050
rect 51662 9998 51714 10050
rect 6190 9886 6242 9938
rect 7422 9886 7474 9938
rect 9550 9886 9602 9938
rect 12798 9886 12850 9938
rect 14254 9886 14306 9938
rect 16382 9886 16434 9938
rect 16718 9886 16770 9938
rect 17390 9886 17442 9938
rect 21422 9886 21474 9938
rect 21870 9886 21922 9938
rect 22766 9886 22818 9938
rect 24894 9886 24946 9938
rect 25342 9886 25394 9938
rect 25790 9886 25842 9938
rect 31950 9886 32002 9938
rect 33742 9886 33794 9938
rect 35870 9886 35922 9938
rect 37214 9886 37266 9938
rect 41246 9886 41298 9938
rect 42590 9886 42642 9938
rect 43150 9886 43202 9938
rect 48302 9886 48354 9938
rect 50430 9886 50482 9938
rect 53454 9886 53506 9938
rect 54798 9886 54850 9938
rect 56926 9886 56978 9938
rect 61854 9886 61906 9938
rect 63982 9886 64034 9938
rect 65438 9886 65490 9938
rect 69246 9886 69298 9938
rect 71374 9886 71426 9938
rect 4174 9774 4226 9826
rect 4734 9774 4786 9826
rect 5742 9774 5794 9826
rect 10334 9774 10386 9826
rect 12462 9774 12514 9826
rect 13582 9774 13634 9826
rect 19854 9774 19906 9826
rect 20190 9774 20242 9826
rect 20414 9774 20466 9826
rect 20750 9774 20802 9826
rect 31166 9774 31218 9826
rect 32958 9774 33010 9826
rect 37550 9774 37602 9826
rect 38334 9774 38386 9826
rect 46062 9774 46114 9826
rect 46734 9774 46786 9826
rect 47518 9774 47570 9826
rect 52894 9774 52946 9826
rect 54014 9774 54066 9826
rect 61070 9774 61122 9826
rect 68574 9774 68626 9826
rect 71710 9774 71762 9826
rect 72830 9774 72882 9826
rect 73502 9774 73554 9826
rect 74286 9774 74338 9826
rect 76414 9774 76466 9826
rect 3166 9662 3218 9714
rect 3838 9662 3890 9714
rect 4958 9662 5010 9714
rect 17838 9662 17890 9714
rect 19294 9662 19346 9714
rect 19630 9662 19682 9714
rect 26574 9662 26626 9714
rect 31390 9662 31442 9714
rect 31502 9662 31554 9714
rect 32398 9662 32450 9714
rect 39118 9662 39170 9714
rect 45950 9662 46002 9714
rect 47070 9662 47122 9714
rect 51102 9662 51154 9714
rect 51326 9662 51378 9714
rect 57822 9662 57874 9714
rect 64990 9662 65042 9714
rect 65886 9662 65938 9714
rect 66558 9662 66610 9714
rect 72046 9662 72098 9714
rect 73838 9662 73890 9714
rect 77086 9662 77138 9714
rect 2830 9550 2882 9602
rect 12126 9550 12178 9602
rect 19742 9550 19794 9602
rect 20638 9550 20690 9602
rect 26910 9550 26962 9602
rect 41694 9550 41746 9602
rect 43598 9550 43650 9602
rect 44942 9550 44994 9602
rect 51998 9550 52050 9602
rect 52670 9550 52722 9602
rect 57486 9550 57538 9602
rect 66222 9550 66274 9602
rect 73278 9550 73330 9602
rect 73390 9550 73442 9602
rect 76750 9550 76802 9602
rect 20534 9382 20586 9434
rect 20638 9382 20690 9434
rect 20742 9382 20794 9434
rect 39854 9382 39906 9434
rect 39958 9382 40010 9434
rect 40062 9382 40114 9434
rect 59174 9382 59226 9434
rect 59278 9382 59330 9434
rect 59382 9382 59434 9434
rect 78494 9382 78546 9434
rect 78598 9382 78650 9434
rect 78702 9382 78754 9434
rect 6638 9214 6690 9266
rect 7086 9214 7138 9266
rect 7534 9214 7586 9266
rect 7870 9214 7922 9266
rect 9662 9214 9714 9266
rect 13246 9214 13298 9266
rect 14926 9214 14978 9266
rect 34526 9214 34578 9266
rect 39118 9214 39170 9266
rect 49646 9214 49698 9266
rect 56030 9214 56082 9266
rect 61294 9214 61346 9266
rect 61966 9214 62018 9266
rect 68574 9214 68626 9266
rect 68798 9214 68850 9266
rect 69582 9214 69634 9266
rect 69806 9214 69858 9266
rect 71374 9214 71426 9266
rect 72382 9214 72434 9266
rect 73614 9214 73666 9266
rect 73950 9214 74002 9266
rect 5182 9102 5234 9154
rect 5518 9102 5570 9154
rect 8430 9102 8482 9154
rect 10782 9102 10834 9154
rect 11454 9102 11506 9154
rect 12350 9102 12402 9154
rect 12686 9102 12738 9154
rect 13470 9102 13522 9154
rect 13582 9102 13634 9154
rect 14030 9102 14082 9154
rect 19518 9102 19570 9154
rect 22990 9102 23042 9154
rect 26910 9102 26962 9154
rect 30494 9102 30546 9154
rect 35422 9102 35474 9154
rect 38446 9102 38498 9154
rect 47182 9102 47234 9154
rect 47518 9102 47570 9154
rect 48750 9102 48802 9154
rect 52558 9102 52610 9154
rect 57598 9102 57650 9154
rect 62526 9102 62578 9154
rect 63086 9102 63138 9154
rect 63534 9102 63586 9154
rect 65774 9102 65826 9154
rect 4286 8990 4338 9042
rect 5742 8990 5794 9042
rect 8990 8990 9042 9042
rect 10670 8990 10722 9042
rect 18846 8990 18898 9042
rect 23326 8990 23378 9042
rect 26126 8990 26178 9042
rect 30830 8990 30882 9042
rect 34862 8990 34914 9042
rect 35646 8990 35698 9042
rect 36206 8990 36258 9042
rect 38670 8990 38722 9042
rect 39342 8990 39394 9042
rect 46174 8990 46226 9042
rect 47742 8990 47794 9042
rect 48078 8990 48130 9042
rect 48974 8990 49026 9042
rect 53230 8990 53282 9042
rect 56814 8990 56866 9042
rect 62302 8990 62354 9042
rect 63758 8990 63810 9042
rect 65102 8990 65154 9042
rect 69918 8990 69970 9042
rect 70366 8990 70418 9042
rect 72270 8990 72322 9042
rect 72606 8990 72658 9042
rect 76078 8990 76130 9042
rect 21646 8878 21698 8930
rect 29038 8878 29090 8930
rect 34078 8878 34130 8930
rect 37998 8878 38050 8930
rect 43262 8878 43314 8930
rect 45390 8878 45442 8930
rect 50430 8851 50482 8903
rect 59726 8878 59778 8930
rect 60846 8878 60898 8930
rect 67902 8878 67954 8930
rect 69246 8878 69298 8930
rect 72942 8878 72994 8930
rect 1934 8766 1986 8818
rect 6078 8766 6130 8818
rect 9998 8766 10050 8818
rect 11790 8766 11842 8818
rect 12126 8766 12178 8818
rect 77982 8766 78034 8818
rect 10874 8598 10926 8650
rect 10978 8598 11030 8650
rect 11082 8598 11134 8650
rect 30194 8598 30246 8650
rect 30298 8598 30350 8650
rect 30402 8598 30454 8650
rect 49514 8598 49566 8650
rect 49618 8598 49670 8650
rect 49722 8598 49774 8650
rect 68834 8598 68886 8650
rect 68938 8598 68990 8650
rect 69042 8598 69094 8650
rect 26462 8430 26514 8482
rect 57822 8430 57874 8482
rect 2494 8318 2546 8370
rect 4622 8318 4674 8370
rect 5182 8318 5234 8370
rect 32510 8374 32562 8426
rect 66558 8430 66610 8482
rect 9214 8318 9266 8370
rect 12686 8318 12738 8370
rect 14030 8318 14082 8370
rect 17502 8318 17554 8370
rect 18286 8318 18338 8370
rect 19854 8318 19906 8370
rect 21422 8318 21474 8370
rect 22766 8318 22818 8370
rect 24894 8318 24946 8370
rect 30382 8318 30434 8370
rect 34414 8318 34466 8370
rect 40574 8318 40626 8370
rect 47294 8318 47346 8370
rect 49422 8318 49474 8370
rect 58158 8318 58210 8370
rect 63310 8318 63362 8370
rect 66222 8318 66274 8370
rect 67118 8318 67170 8370
rect 73614 8318 73666 8370
rect 1822 8206 1874 8258
rect 5966 8206 6018 8258
rect 9886 8206 9938 8258
rect 14590 8206 14642 8258
rect 19070 8206 19122 8258
rect 20078 8206 20130 8258
rect 20750 8206 20802 8258
rect 21982 8206 22034 8258
rect 26798 8206 26850 8258
rect 27470 8206 27522 8258
rect 28142 8206 28194 8258
rect 29710 8206 29762 8258
rect 34974 8206 35026 8258
rect 35646 8206 35698 8258
rect 37438 8206 37490 8258
rect 38222 8206 38274 8258
rect 44942 8206 44994 8258
rect 46510 8206 46562 8258
rect 56702 8206 56754 8258
rect 65662 8206 65714 8258
rect 70702 8206 70754 8258
rect 10558 8094 10610 8146
rect 15374 8094 15426 8146
rect 18846 8094 18898 8146
rect 20190 8094 20242 8146
rect 20414 8094 20466 8146
rect 27358 8094 27410 8146
rect 37102 8094 37154 8146
rect 38110 8094 38162 8146
rect 39566 8094 39618 8146
rect 45166 8094 45218 8146
rect 57150 8094 57202 8146
rect 58382 8094 58434 8146
rect 58718 8094 58770 8146
rect 65550 8094 65602 8146
rect 71486 8094 71538 8146
rect 5630 7982 5682 8034
rect 13582 7982 13634 8034
rect 17950 7982 18002 8034
rect 20638 7982 20690 8034
rect 26014 7982 26066 8034
rect 34750 7982 34802 8034
rect 35870 7982 35922 8034
rect 38782 7982 38834 8034
rect 39902 7982 39954 8034
rect 55246 7982 55298 8034
rect 69806 7982 69858 8034
rect 70366 7982 70418 8034
rect 20534 7814 20586 7866
rect 20638 7814 20690 7866
rect 20742 7814 20794 7866
rect 39854 7814 39906 7866
rect 39958 7814 40010 7866
rect 40062 7814 40114 7866
rect 59174 7814 59226 7866
rect 59278 7814 59330 7866
rect 59382 7814 59434 7866
rect 78494 7814 78546 7866
rect 78598 7814 78650 7866
rect 78702 7814 78754 7866
rect 9662 7646 9714 7698
rect 10782 7646 10834 7698
rect 15598 7646 15650 7698
rect 17502 7646 17554 7698
rect 19518 7646 19570 7698
rect 20526 7646 20578 7698
rect 23438 7646 23490 7698
rect 25342 7646 25394 7698
rect 31054 7646 31106 7698
rect 33182 7646 33234 7698
rect 41022 7646 41074 7698
rect 41470 7646 41522 7698
rect 44606 7646 44658 7698
rect 72382 7646 72434 7698
rect 72494 7646 72546 7698
rect 72718 7646 72770 7698
rect 2382 7534 2434 7586
rect 2718 7534 2770 7586
rect 3838 7534 3890 7586
rect 8654 7534 8706 7586
rect 11118 7534 11170 7586
rect 15934 7534 15986 7586
rect 23998 7534 24050 7586
rect 24334 7534 24386 7586
rect 25902 7534 25954 7586
rect 31726 7534 31778 7586
rect 32174 7534 32226 7586
rect 36542 7534 36594 7586
rect 40126 7534 40178 7586
rect 42590 7534 42642 7586
rect 43934 7534 43986 7586
rect 55582 7534 55634 7586
rect 62974 7534 63026 7586
rect 69694 7534 69746 7586
rect 70366 7534 70418 7586
rect 76750 7534 76802 7586
rect 3054 7422 3106 7474
rect 8094 7422 8146 7474
rect 8878 7422 8930 7474
rect 23774 7422 23826 7474
rect 31390 7422 31442 7474
rect 37326 7422 37378 7474
rect 39454 7422 39506 7474
rect 40238 7422 40290 7474
rect 44046 7422 44098 7474
rect 52446 7422 52498 7474
rect 55806 7422 55858 7474
rect 62638 7422 62690 7474
rect 69918 7422 69970 7474
rect 70702 7422 70754 7474
rect 71150 7422 71202 7474
rect 72270 7422 72322 7474
rect 76974 7422 77026 7474
rect 5966 7310 6018 7362
rect 7422 7310 7474 7362
rect 34414 7310 34466 7362
rect 53118 7310 53170 7362
rect 55246 7310 55298 7362
rect 68910 7310 68962 7362
rect 69246 7310 69298 7362
rect 71486 7310 71538 7362
rect 73278 7310 73330 7362
rect 76526 7310 76578 7362
rect 7758 7198 7810 7250
rect 39118 7198 39170 7250
rect 42926 7198 42978 7250
rect 43262 7198 43314 7250
rect 10874 7030 10926 7082
rect 10978 7030 11030 7082
rect 11082 7030 11134 7082
rect 30194 7030 30246 7082
rect 30298 7030 30350 7082
rect 30402 7030 30454 7082
rect 49514 7030 49566 7082
rect 49618 7030 49670 7082
rect 49722 7030 49774 7082
rect 68834 7030 68886 7082
rect 68938 7030 68990 7082
rect 69042 7030 69094 7082
rect 48974 6862 49026 6914
rect 54686 6862 54738 6914
rect 58830 6862 58882 6914
rect 59502 6862 59554 6914
rect 60062 6862 60114 6914
rect 14254 6750 14306 6802
rect 25006 6750 25058 6802
rect 28142 6750 28194 6802
rect 39678 6750 39730 6802
rect 41918 6750 41970 6802
rect 61966 6750 62018 6802
rect 4286 6638 4338 6690
rect 4846 6638 4898 6690
rect 11342 6638 11394 6690
rect 13694 6638 13746 6690
rect 25566 6638 25618 6690
rect 32622 6638 32674 6690
rect 39006 6638 39058 6690
rect 42926 6638 42978 6690
rect 43262 6638 43314 6690
rect 55470 6638 55522 6690
rect 56030 6638 56082 6690
rect 57262 6638 57314 6690
rect 58270 6638 58322 6690
rect 59166 6638 59218 6690
rect 64094 6638 64146 6690
rect 64878 6638 64930 6690
rect 65326 6638 65378 6690
rect 66222 6638 66274 6690
rect 69694 6638 69746 6690
rect 70702 6638 70754 6690
rect 71710 6638 71762 6690
rect 2494 6526 2546 6578
rect 11006 6526 11058 6578
rect 20078 6526 20130 6578
rect 20414 6526 20466 6578
rect 21646 6526 21698 6578
rect 26574 6526 26626 6578
rect 26910 6526 26962 6578
rect 27470 6526 27522 6578
rect 27918 6526 27970 6578
rect 35758 6526 35810 6578
rect 36094 6526 36146 6578
rect 49198 6526 49250 6578
rect 49758 6526 49810 6578
rect 50430 6526 50482 6578
rect 53342 6526 53394 6578
rect 53678 6526 53730 6578
rect 54350 6526 54402 6578
rect 55246 6526 55298 6578
rect 58046 6526 58098 6578
rect 65662 6526 65714 6578
rect 68686 6526 68738 6578
rect 69022 6526 69074 6578
rect 70926 6526 70978 6578
rect 71262 6526 71314 6578
rect 13470 6414 13522 6466
rect 21310 6414 21362 6466
rect 25342 6414 25394 6466
rect 28478 6414 28530 6466
rect 29374 6414 29426 6466
rect 35422 6414 35474 6466
rect 43598 6414 43650 6466
rect 48638 6414 48690 6466
rect 57598 6414 57650 6466
rect 59726 6414 59778 6466
rect 60622 6414 60674 6466
rect 61742 6414 61794 6466
rect 67342 6414 67394 6466
rect 69358 6414 69410 6466
rect 70030 6414 70082 6466
rect 70142 6414 70194 6466
rect 70254 6414 70306 6466
rect 72270 6414 72322 6466
rect 72606 6414 72658 6466
rect 20534 6246 20586 6298
rect 20638 6246 20690 6298
rect 20742 6246 20794 6298
rect 39854 6246 39906 6298
rect 39958 6246 40010 6298
rect 40062 6246 40114 6298
rect 59174 6246 59226 6298
rect 59278 6246 59330 6298
rect 59382 6246 59434 6298
rect 78494 6246 78546 6298
rect 78598 6246 78650 6298
rect 78702 6246 78754 6298
rect 10110 6078 10162 6130
rect 10782 6078 10834 6130
rect 13134 6078 13186 6130
rect 14254 6078 14306 6130
rect 19742 6078 19794 6130
rect 21310 6078 21362 6130
rect 26014 6078 26066 6130
rect 36206 6078 36258 6130
rect 37102 6078 37154 6130
rect 37998 6078 38050 6130
rect 42702 6078 42754 6130
rect 51774 6078 51826 6130
rect 55358 6078 55410 6130
rect 55694 6078 55746 6130
rect 56590 6078 56642 6130
rect 62638 6078 62690 6130
rect 67118 6078 67170 6130
rect 71374 6078 71426 6130
rect 72158 6078 72210 6130
rect 72382 6078 72434 6130
rect 72942 6078 72994 6130
rect 73390 6078 73442 6130
rect 11118 5966 11170 6018
rect 12462 5966 12514 6018
rect 15822 5966 15874 6018
rect 16158 5966 16210 6018
rect 16830 5966 16882 6018
rect 18510 5966 18562 6018
rect 20414 5966 20466 6018
rect 21982 5966 22034 6018
rect 23438 5966 23490 6018
rect 32174 5966 32226 6018
rect 32510 5966 32562 6018
rect 33294 5966 33346 6018
rect 35198 5966 35250 6018
rect 37438 5966 37490 6018
rect 42366 5966 42418 6018
rect 43822 5966 43874 6018
rect 48190 5966 48242 6018
rect 49534 5966 49586 6018
rect 56030 5966 56082 6018
rect 58158 5966 58210 6018
rect 61742 5966 61794 6018
rect 63198 5966 63250 6018
rect 63534 5966 63586 6018
rect 65662 5966 65714 6018
rect 66334 5966 66386 6018
rect 8990 5854 9042 5906
rect 10334 5854 10386 5906
rect 12686 5854 12738 5906
rect 14590 5854 14642 5906
rect 16606 5854 16658 5906
rect 17838 5854 17890 5906
rect 18398 5854 18450 5906
rect 19966 5854 20018 5906
rect 20638 5854 20690 5906
rect 21758 5854 21810 5906
rect 23550 5854 23602 5906
rect 26350 5854 26402 5906
rect 29486 5854 29538 5906
rect 33630 5854 33682 5906
rect 34302 5854 34354 5906
rect 34638 5854 34690 5906
rect 35310 5854 35362 5906
rect 43038 5854 43090 5906
rect 47966 5854 48018 5906
rect 48862 5854 48914 5906
rect 56926 5854 56978 5906
rect 57486 5854 57538 5906
rect 60846 5854 60898 5906
rect 62078 5854 62130 5906
rect 62974 5854 63026 5906
rect 65438 5854 65490 5906
rect 65886 5854 65938 5906
rect 66670 5854 66722 5906
rect 70030 5854 70082 5906
rect 70590 5854 70642 5906
rect 71598 5854 71650 5906
rect 72494 5854 72546 5906
rect 76078 5854 76130 5906
rect 6078 5742 6130 5794
rect 8206 5742 8258 5794
rect 13582 5742 13634 5794
rect 15038 5742 15090 5794
rect 19294 5742 19346 5794
rect 24222 5742 24274 5794
rect 26686 5742 26738 5794
rect 28814 5742 28866 5794
rect 36654 5742 36706 5794
rect 38670 5742 38722 5794
rect 45950 5742 46002 5794
rect 55022 5742 55074 5794
rect 60286 5742 60338 5794
rect 61406 5742 61458 5794
rect 69358 5742 69410 5794
rect 70926 5742 70978 5794
rect 77982 5742 78034 5794
rect 11566 5630 11618 5682
rect 11902 5630 11954 5682
rect 17502 5630 17554 5682
rect 22430 5630 22482 5682
rect 22766 5630 22818 5682
rect 55022 5630 55074 5682
rect 55358 5630 55410 5682
rect 10874 5462 10926 5514
rect 10978 5462 11030 5514
rect 11082 5462 11134 5514
rect 30194 5462 30246 5514
rect 30298 5462 30350 5514
rect 30402 5462 30454 5514
rect 49514 5462 49566 5514
rect 49618 5462 49670 5514
rect 49722 5462 49774 5514
rect 68834 5462 68886 5514
rect 68938 5462 68990 5514
rect 69042 5462 69094 5514
rect 45278 5294 45330 5346
rect 54574 5294 54626 5346
rect 62190 5294 62242 5346
rect 62526 5294 62578 5346
rect 66670 5294 66722 5346
rect 12910 5182 12962 5234
rect 13918 5182 13970 5234
rect 17054 5182 17106 5234
rect 19182 5182 19234 5234
rect 22206 5182 22258 5234
rect 24334 5182 24386 5234
rect 28478 5182 28530 5234
rect 32734 5182 32786 5234
rect 34862 5182 34914 5234
rect 37438 5182 37490 5234
rect 41806 5182 41858 5234
rect 46622 5182 46674 5234
rect 47070 5182 47122 5234
rect 50654 5182 50706 5234
rect 59390 5182 59442 5234
rect 59950 5182 60002 5234
rect 68462 5182 68514 5234
rect 70254 5182 70306 5234
rect 72494 5182 72546 5234
rect 76974 5182 77026 5234
rect 7534 5070 7586 5122
rect 8990 5070 9042 5122
rect 9998 5070 10050 5122
rect 14702 5070 14754 5122
rect 15710 5070 15762 5122
rect 16270 5070 16322 5122
rect 20750 5070 20802 5122
rect 21534 5070 21586 5122
rect 25678 5070 25730 5122
rect 29486 5070 29538 5122
rect 31950 5070 32002 5122
rect 35422 5070 35474 5122
rect 36206 5070 36258 5122
rect 37102 5070 37154 5122
rect 38222 5070 38274 5122
rect 39006 5070 39058 5122
rect 42702 5070 42754 5122
rect 44270 5070 44322 5122
rect 44942 5070 44994 5122
rect 45726 5070 45778 5122
rect 47854 5070 47906 5122
rect 53006 5070 53058 5122
rect 53566 5070 53618 5122
rect 54238 5070 54290 5122
rect 55358 5070 55410 5122
rect 55918 5070 55970 5122
rect 57150 5070 57202 5122
rect 57822 5070 57874 5122
rect 58158 5070 58210 5122
rect 58830 5070 58882 5122
rect 60734 5070 60786 5122
rect 61182 5070 61234 5122
rect 61630 5070 61682 5122
rect 62974 5070 63026 5122
rect 63870 5070 63922 5122
rect 65102 5070 65154 5122
rect 65774 5070 65826 5122
rect 66334 5070 66386 5122
rect 67230 5070 67282 5122
rect 67566 5070 67618 5122
rect 67902 5070 67954 5122
rect 68350 5070 68402 5122
rect 69022 5070 69074 5122
rect 69582 5070 69634 5122
rect 75742 5070 75794 5122
rect 76414 5070 76466 5122
rect 7758 4958 7810 5010
rect 10782 4958 10834 5010
rect 14478 4958 14530 5010
rect 26350 4958 26402 5010
rect 29150 4958 29202 5010
rect 31614 4958 31666 5010
rect 35982 4958 36034 5010
rect 38110 4958 38162 5010
rect 39678 4958 39730 5010
rect 43262 4958 43314 5010
rect 43598 4958 43650 5010
rect 43934 4958 43986 5010
rect 46062 4958 46114 5010
rect 48526 4958 48578 5010
rect 52670 4958 52722 5010
rect 55246 4958 55298 5010
rect 56254 4958 56306 5010
rect 57262 4958 57314 5010
rect 60510 4958 60562 5010
rect 63310 4958 63362 5010
rect 64766 4958 64818 5010
rect 65550 4958 65602 5010
rect 67678 4958 67730 5010
rect 68574 4958 68626 5010
rect 9214 4846 9266 4898
rect 13582 4846 13634 4898
rect 15374 4846 15426 4898
rect 20414 4846 20466 4898
rect 31278 4846 31330 4898
rect 35646 4846 35698 4898
rect 42926 4846 42978 4898
rect 53342 4846 53394 4898
rect 58606 4846 58658 4898
rect 20534 4678 20586 4730
rect 20638 4678 20690 4730
rect 20742 4678 20794 4730
rect 39854 4678 39906 4730
rect 39958 4678 40010 4730
rect 40062 4678 40114 4730
rect 59174 4678 59226 4730
rect 59278 4678 59330 4730
rect 59382 4678 59434 4730
rect 78494 4678 78546 4730
rect 78598 4678 78650 4730
rect 78702 4678 78754 4730
rect 12798 4510 12850 4562
rect 17614 4510 17666 4562
rect 23326 4510 23378 4562
rect 26126 4510 26178 4562
rect 33294 4510 33346 4562
rect 35086 4510 35138 4562
rect 40014 4510 40066 4562
rect 42814 4510 42866 4562
rect 48190 4510 48242 4562
rect 50654 4510 50706 4562
rect 10334 4398 10386 4450
rect 13134 4398 13186 4450
rect 14702 4398 14754 4450
rect 18510 4398 18562 4450
rect 20638 4398 20690 4450
rect 23886 4398 23938 4450
rect 24446 4398 24498 4450
rect 25790 4398 25842 4450
rect 27806 4398 27858 4450
rect 30382 4398 30434 4450
rect 34190 4398 34242 4450
rect 37662 4398 37714 4450
rect 42142 4398 42194 4450
rect 44382 4398 44434 4450
rect 49422 4398 49474 4450
rect 49870 4398 49922 4450
rect 53006 4398 53058 4450
rect 56030 4398 56082 4450
rect 57374 4398 57426 4450
rect 61406 4398 61458 4450
rect 65998 4398 66050 4450
rect 4286 4286 4338 4338
rect 9662 4286 9714 4338
rect 14030 4286 14082 4338
rect 17950 4286 18002 4338
rect 18734 4286 18786 4338
rect 19406 4286 19458 4338
rect 19854 4286 19906 4338
rect 23662 4286 23714 4338
rect 25454 4286 25506 4338
rect 26462 4286 26514 4338
rect 26910 4286 26962 4338
rect 27246 4286 27298 4338
rect 28030 4286 28082 4338
rect 29710 4286 29762 4338
rect 33630 4286 33682 4338
rect 34414 4286 34466 4338
rect 38446 4286 38498 4338
rect 40350 4286 40402 4338
rect 41022 4286 41074 4338
rect 41358 4286 41410 4338
rect 42030 4286 42082 4338
rect 43710 4286 43762 4338
rect 47966 4286 48018 4338
rect 48862 4286 48914 4338
rect 49198 4286 49250 4338
rect 52334 4286 52386 4338
rect 55806 4286 55858 4338
rect 56590 4286 56642 4338
rect 60622 4286 60674 4338
rect 65214 4286 65266 4338
rect 68686 4286 68738 4338
rect 75630 4286 75682 4338
rect 4734 4174 4786 4226
rect 5182 4174 5234 4226
rect 12462 4174 12514 4226
rect 16830 4174 16882 4226
rect 22766 4174 22818 4226
rect 32510 4174 32562 4226
rect 35534 4174 35586 4226
rect 46510 4174 46562 4226
rect 55134 4174 55186 4226
rect 59502 4174 59554 4226
rect 63534 4174 63586 4226
rect 68126 4174 68178 4226
rect 1934 4062 1986 4114
rect 69470 4062 69522 4114
rect 77982 4062 78034 4114
rect 10874 3894 10926 3946
rect 10978 3894 11030 3946
rect 11082 3894 11134 3946
rect 30194 3894 30246 3946
rect 30298 3894 30350 3946
rect 30402 3894 30454 3946
rect 49514 3894 49566 3946
rect 49618 3894 49670 3946
rect 49722 3894 49774 3946
rect 68834 3894 68886 3946
rect 68938 3894 68990 3946
rect 69042 3894 69094 3946
rect 1934 3614 1986 3666
rect 5742 3614 5794 3666
rect 36878 3614 36930 3666
rect 57038 3614 57090 3666
rect 64766 3614 64818 3666
rect 67118 3614 67170 3666
rect 68350 3614 68402 3666
rect 68686 3614 68738 3666
rect 4286 3502 4338 3554
rect 4734 3502 4786 3554
rect 20302 3502 20354 3554
rect 20974 3502 21026 3554
rect 24782 3502 24834 3554
rect 67902 3502 67954 3554
rect 72606 3502 72658 3554
rect 77198 3502 77250 3554
rect 4958 3390 5010 3442
rect 7646 3390 7698 3442
rect 7870 3390 7922 3442
rect 8206 3390 8258 3442
rect 11678 3390 11730 3442
rect 11902 3390 11954 3442
rect 12238 3390 12290 3442
rect 15710 3390 15762 3442
rect 15934 3390 15986 3442
rect 16270 3390 16322 3442
rect 20750 3390 20802 3442
rect 24110 3390 24162 3442
rect 27918 3390 27970 3442
rect 28366 3390 28418 3442
rect 28702 3390 28754 3442
rect 31726 3390 31778 3442
rect 32174 3390 32226 3442
rect 32510 3390 32562 3442
rect 35534 3390 35586 3442
rect 36094 3390 36146 3442
rect 36430 3390 36482 3442
rect 39342 3390 39394 3442
rect 40126 3390 40178 3442
rect 40462 3390 40514 3442
rect 43934 3390 43986 3442
rect 44158 3390 44210 3442
rect 44494 3390 44546 3442
rect 47966 3390 48018 3442
rect 48190 3390 48242 3442
rect 48526 3390 48578 3442
rect 51998 3390 52050 3442
rect 52222 3390 52274 3442
rect 52558 3390 52610 3442
rect 56030 3390 56082 3442
rect 56254 3390 56306 3442
rect 56590 3390 56642 3442
rect 60062 3390 60114 3442
rect 60286 3390 60338 3442
rect 60622 3390 60674 3442
rect 64094 3390 64146 3442
rect 64318 3390 64370 3442
rect 72158 3390 72210 3442
rect 75518 3390 75570 3442
rect 24558 3278 24610 3330
rect 72382 3278 72434 3330
rect 20534 3110 20586 3162
rect 20638 3110 20690 3162
rect 20742 3110 20794 3162
rect 39854 3110 39906 3162
rect 39958 3110 40010 3162
rect 40062 3110 40114 3162
rect 59174 3110 59226 3162
rect 59278 3110 59330 3162
rect 59382 3110 59434 3162
rect 78494 3110 78546 3162
rect 78598 3110 78650 3162
rect 78702 3110 78754 3162
<< metal2 >>
rect 1568 39200 1680 40000
rect 4032 39200 4144 40000
rect 6496 39200 6608 40000
rect 8960 39200 9072 40000
rect 11424 39200 11536 40000
rect 13888 39200 14000 40000
rect 16352 39200 16464 40000
rect 18816 39200 18928 40000
rect 21280 39200 21392 40000
rect 23744 39200 23856 40000
rect 26208 39200 26320 40000
rect 28672 39200 28784 40000
rect 31136 39200 31248 40000
rect 33600 39200 33712 40000
rect 35532 39228 35924 39284
rect 1596 35252 1652 39200
rect 3388 38388 3444 38398
rect 1932 36594 1988 36606
rect 1932 36542 1934 36594
rect 1986 36542 1988 36594
rect 1932 35924 1988 36542
rect 1932 35858 1988 35868
rect 3276 35924 3332 35934
rect 3388 35924 3444 38332
rect 3276 35922 3444 35924
rect 3276 35870 3278 35922
rect 3330 35870 3444 35922
rect 3276 35868 3444 35870
rect 3948 36482 4004 36494
rect 3948 36430 3950 36482
rect 4002 36430 4004 36482
rect 3276 35858 3332 35868
rect 1596 35196 1876 35252
rect 1820 35028 1876 35196
rect 2940 35140 2996 35150
rect 2940 35046 2996 35084
rect 3948 35140 4004 36430
rect 4060 35924 4116 39200
rect 6524 36596 6580 39200
rect 8876 36596 8932 36606
rect 8988 36596 9044 39200
rect 10872 36876 11136 36886
rect 10928 36820 10976 36876
rect 11032 36820 11080 36876
rect 10872 36810 11136 36820
rect 11452 36596 11508 39200
rect 13916 36596 13972 39200
rect 14476 37604 14532 37614
rect 6524 36594 6804 36596
rect 6524 36542 6526 36594
rect 6578 36542 6804 36594
rect 6524 36540 6804 36542
rect 6524 36530 6580 36540
rect 6748 36482 6804 36540
rect 8876 36594 9380 36596
rect 8876 36542 8878 36594
rect 8930 36542 9380 36594
rect 8876 36540 9380 36542
rect 8876 36530 8932 36540
rect 6748 36430 6750 36482
rect 6802 36430 6804 36482
rect 6748 36418 6804 36430
rect 9324 36482 9380 36540
rect 11452 36594 11732 36596
rect 11452 36542 11454 36594
rect 11506 36542 11732 36594
rect 11452 36540 11732 36542
rect 11452 36530 11508 36540
rect 9324 36430 9326 36482
rect 9378 36430 9380 36482
rect 9324 36418 9380 36430
rect 11676 36482 11732 36540
rect 13916 36594 14196 36596
rect 13916 36542 13918 36594
rect 13970 36542 14196 36594
rect 13916 36540 14196 36542
rect 13916 36530 13972 36540
rect 11676 36430 11678 36482
rect 11730 36430 11732 36482
rect 11676 36418 11732 36430
rect 14140 36482 14196 36540
rect 14140 36430 14142 36482
rect 14194 36430 14196 36482
rect 14140 36418 14196 36430
rect 7308 36372 7364 36382
rect 7308 36278 7364 36316
rect 9884 36370 9940 36382
rect 9884 36318 9886 36370
rect 9938 36318 9940 36370
rect 4620 35924 4676 35934
rect 4060 35922 4676 35924
rect 4060 35870 4622 35922
rect 4674 35870 4676 35922
rect 4060 35868 4676 35870
rect 3948 35074 4004 35084
rect 4284 35698 4340 35710
rect 4284 35646 4286 35698
rect 4338 35646 4340 35698
rect 1820 34914 1876 34972
rect 3500 35028 3556 35038
rect 3500 34934 3556 34972
rect 1820 34862 1822 34914
rect 1874 34862 1876 34914
rect 1820 34850 1876 34862
rect 2380 34914 2436 34926
rect 2380 34862 2382 34914
rect 2434 34862 2436 34914
rect 1932 33906 1988 33918
rect 1932 33854 1934 33906
rect 1986 33854 1988 33906
rect 1932 33460 1988 33854
rect 1932 33394 1988 33404
rect 1932 31890 1988 31902
rect 1932 31838 1934 31890
rect 1986 31838 1988 31890
rect 1932 30996 1988 31838
rect 1932 30930 1988 30940
rect 2268 28756 2324 28766
rect 2268 28642 2324 28700
rect 2268 28590 2270 28642
rect 2322 28590 2324 28642
rect 1932 28532 1988 28542
rect 1932 27746 1988 28476
rect 1932 27694 1934 27746
rect 1986 27694 1988 27746
rect 1932 27682 1988 27694
rect 1820 26740 1876 26750
rect 1708 26684 1820 26740
rect 1708 22932 1764 26684
rect 1820 26674 1876 26684
rect 1820 26290 1876 26302
rect 1820 26238 1822 26290
rect 1874 26238 1876 26290
rect 1820 23940 1876 26238
rect 1932 26068 1988 26078
rect 1932 25730 1988 26012
rect 1932 25678 1934 25730
rect 1986 25678 1988 25730
rect 1932 25666 1988 25678
rect 1820 23156 1876 23884
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 1820 23154 1988 23156
rect 1820 23102 1822 23154
rect 1874 23102 1988 23154
rect 1820 23100 1988 23102
rect 1820 23090 1876 23100
rect 1932 23044 1988 23100
rect 1932 22988 2212 23044
rect 1708 22876 2100 22932
rect 2044 22482 2100 22876
rect 2044 22430 2046 22482
rect 2098 22430 2100 22482
rect 2044 22260 2100 22430
rect 1708 22204 2100 22260
rect 1708 21698 1764 22204
rect 1708 21646 1710 21698
rect 1762 21646 1764 21698
rect 1708 21634 1764 21646
rect 2156 21810 2212 22988
rect 2156 21758 2158 21810
rect 2210 21758 2212 21810
rect 1820 21362 1876 21374
rect 1820 21310 1822 21362
rect 1874 21310 1876 21362
rect 1820 20802 1876 21310
rect 2156 21364 2212 21758
rect 2268 21588 2324 28590
rect 2380 23380 2436 34862
rect 3052 34802 3108 34814
rect 3052 34750 3054 34802
rect 3106 34750 3108 34802
rect 3052 34356 3108 34750
rect 4284 34692 4340 35646
rect 4396 35026 4452 35868
rect 4620 35858 4676 35868
rect 4396 34974 4398 35026
rect 4450 34974 4452 35026
rect 4396 34962 4452 34974
rect 5180 35586 5236 35598
rect 5180 35534 5182 35586
rect 5234 35534 5236 35586
rect 4732 34692 4788 34702
rect 4284 34690 4788 34692
rect 4284 34638 4734 34690
rect 4786 34638 4788 34690
rect 4284 34636 4788 34638
rect 3108 34300 3332 34356
rect 3052 34290 3108 34300
rect 3276 33458 3332 34300
rect 4284 34130 4340 34142
rect 4284 34078 4286 34130
rect 4338 34078 4340 34130
rect 4284 34020 4340 34078
rect 4284 33954 4340 33964
rect 3276 33406 3278 33458
rect 3330 33406 3332 33458
rect 3276 33394 3332 33406
rect 4732 33348 4788 34636
rect 4844 34020 4900 34030
rect 4844 33926 4900 33964
rect 4732 33282 4788 33292
rect 4284 31780 4340 31790
rect 4284 31686 4340 31724
rect 4060 31220 4116 31230
rect 3948 31164 4060 31220
rect 3724 30100 3780 30110
rect 3724 30006 3780 30044
rect 3388 29988 3444 29998
rect 3164 29986 3444 29988
rect 3164 29934 3390 29986
rect 3442 29934 3444 29986
rect 3164 29932 3444 29934
rect 3164 29538 3220 29932
rect 3388 29922 3444 29932
rect 3164 29486 3166 29538
rect 3218 29486 3220 29538
rect 3164 29474 3220 29486
rect 2492 29428 2548 29438
rect 2492 29334 2548 29372
rect 2940 28644 2996 28654
rect 2940 28550 2996 28588
rect 3164 26964 3220 26974
rect 3164 26962 3332 26964
rect 3164 26910 3166 26962
rect 3218 26910 3332 26962
rect 3164 26908 3332 26910
rect 3164 26898 3220 26908
rect 2828 26852 2884 26862
rect 2492 26850 2884 26852
rect 2492 26798 2830 26850
rect 2882 26798 2884 26850
rect 2492 26796 2884 26798
rect 2492 26402 2548 26796
rect 2828 26786 2884 26796
rect 2492 26350 2494 26402
rect 2546 26350 2548 26402
rect 2492 26338 2548 26350
rect 3276 25844 3332 26908
rect 3276 25788 3780 25844
rect 3724 24946 3780 25788
rect 3724 24894 3726 24946
rect 3778 24894 3780 24946
rect 3724 24882 3780 24894
rect 2380 23314 2436 23324
rect 2492 23044 2548 23054
rect 2492 23042 2884 23044
rect 2492 22990 2494 23042
rect 2546 22990 2884 23042
rect 2492 22988 2884 22990
rect 2492 22978 2548 22988
rect 2828 22258 2884 22988
rect 2828 22206 2830 22258
rect 2882 22206 2884 22258
rect 2828 22194 2884 22206
rect 3164 22260 3220 22270
rect 3164 22166 3220 22204
rect 3836 22260 3892 22270
rect 3836 22166 3892 22204
rect 3948 21700 4004 31164
rect 4060 31154 4116 31164
rect 5180 31108 5236 35534
rect 9884 35028 9940 36318
rect 12236 36370 12292 36382
rect 12236 36318 12238 36370
rect 12290 36318 12292 36370
rect 9884 34962 9940 34972
rect 10332 35698 10388 35710
rect 10332 35646 10334 35698
rect 10386 35646 10388 35698
rect 10332 34132 10388 35646
rect 11004 35588 11060 35598
rect 11004 35586 11284 35588
rect 11004 35534 11006 35586
rect 11058 35534 11284 35586
rect 11004 35532 11284 35534
rect 11004 35522 11060 35532
rect 10872 35308 11136 35318
rect 10928 35252 10976 35308
rect 11032 35252 11080 35308
rect 10872 35242 11136 35252
rect 10332 34066 10388 34076
rect 11004 34132 11060 34142
rect 11004 34038 11060 34076
rect 10872 33740 11136 33750
rect 10928 33684 10976 33740
rect 11032 33684 11080 33740
rect 10872 33674 11136 33684
rect 11228 33460 11284 35532
rect 12236 35364 12292 36318
rect 14476 36370 14532 37548
rect 16380 36594 16436 39200
rect 16380 36542 16382 36594
rect 16434 36542 16436 36594
rect 16380 36484 16436 36542
rect 18844 36596 18900 39200
rect 20860 37380 20916 37390
rect 19628 36708 19684 36718
rect 18844 36594 19124 36596
rect 18844 36542 18846 36594
rect 18898 36542 19124 36594
rect 18844 36540 19124 36542
rect 18844 36530 18900 36540
rect 16380 36418 16436 36428
rect 17052 36484 17108 36494
rect 17052 36390 17108 36428
rect 19068 36482 19124 36540
rect 19628 36594 19684 36652
rect 19628 36542 19630 36594
rect 19682 36542 19684 36594
rect 19628 36530 19684 36542
rect 19068 36430 19070 36482
rect 19122 36430 19124 36482
rect 19068 36418 19124 36430
rect 14476 36318 14478 36370
rect 14530 36318 14532 36370
rect 14476 36306 14532 36318
rect 13804 36260 13860 36270
rect 13804 35700 13860 36204
rect 17276 36258 17332 36270
rect 17276 36206 17278 36258
rect 17330 36206 17332 36258
rect 17276 35924 17332 36206
rect 17724 36260 17780 36270
rect 17724 36166 17780 36204
rect 20532 36092 20796 36102
rect 20588 36036 20636 36092
rect 20692 36036 20740 36092
rect 20532 36026 20796 36036
rect 17276 35858 17332 35868
rect 14700 35812 14756 35822
rect 13580 35698 14308 35700
rect 13580 35646 13806 35698
rect 13858 35646 14308 35698
rect 13580 35644 14308 35646
rect 13244 35588 13300 35598
rect 13244 35494 13300 35532
rect 12236 35298 12292 35308
rect 13580 35026 13636 35644
rect 13580 34974 13582 35026
rect 13634 34974 13636 35026
rect 13580 34962 13636 34974
rect 13804 34132 13860 35644
rect 14252 35026 14308 35644
rect 14252 34974 14254 35026
rect 14306 34974 14308 35026
rect 14252 34962 14308 34974
rect 14476 35586 14532 35598
rect 14476 35534 14478 35586
rect 14530 35534 14532 35586
rect 14476 34468 14532 35534
rect 14700 35028 14756 35756
rect 17724 35812 17780 35822
rect 17724 35810 17892 35812
rect 17724 35758 17726 35810
rect 17778 35758 17892 35810
rect 17724 35756 17892 35758
rect 17724 35746 17780 35756
rect 17612 35700 17668 35710
rect 17500 35698 17668 35700
rect 17500 35646 17614 35698
rect 17666 35646 17668 35698
rect 17500 35644 17668 35646
rect 15372 35588 15428 35598
rect 14700 35026 14868 35028
rect 14700 34974 14702 35026
rect 14754 34974 14868 35026
rect 14700 34972 14868 34974
rect 14700 34962 14756 34972
rect 14476 34402 14532 34412
rect 13916 34354 13972 34366
rect 13916 34302 13918 34354
rect 13970 34302 13972 34354
rect 13916 34244 13972 34302
rect 14812 34244 14868 34972
rect 15372 34916 15428 35532
rect 16604 35586 16660 35598
rect 16604 35534 16606 35586
rect 16658 35534 16660 35586
rect 16604 35476 16660 35534
rect 16604 35410 16660 35420
rect 17052 35476 17108 35486
rect 16268 34916 16324 34926
rect 15372 34822 15428 34860
rect 15708 34860 16100 34916
rect 15708 34802 15764 34860
rect 15708 34750 15710 34802
rect 15762 34750 15764 34802
rect 15708 34738 15764 34750
rect 15596 34692 15652 34702
rect 13916 34188 14868 34244
rect 11676 34018 11732 34030
rect 11676 33966 11678 34018
rect 11730 33966 11732 34018
rect 11676 33572 11732 33966
rect 11676 33506 11732 33516
rect 12572 33572 12628 33582
rect 12572 33478 12628 33516
rect 11228 33394 11284 33404
rect 13468 33460 13524 33470
rect 13468 33366 13524 33404
rect 12684 33234 12740 33246
rect 12684 33182 12686 33234
rect 12738 33182 12740 33234
rect 12684 32788 12740 33182
rect 13580 33236 13636 33246
rect 13580 33142 13636 33180
rect 13804 33012 13860 34076
rect 14812 34130 14868 34188
rect 15484 34690 15652 34692
rect 15484 34638 15598 34690
rect 15650 34638 15652 34690
rect 15484 34636 15652 34638
rect 14812 34078 14814 34130
rect 14866 34078 14868 34130
rect 14812 34066 14868 34078
rect 15372 34132 15428 34142
rect 15484 34132 15540 34636
rect 15596 34626 15652 34636
rect 15932 34692 15988 34702
rect 15932 34598 15988 34636
rect 16044 34580 16100 34860
rect 16268 34822 16324 34860
rect 16492 34914 16548 34926
rect 16492 34862 16494 34914
rect 16546 34862 16548 34914
rect 16492 34580 16548 34862
rect 16044 34524 16548 34580
rect 16940 34916 16996 34926
rect 15372 34130 15540 34132
rect 15372 34078 15374 34130
rect 15426 34078 15540 34130
rect 15372 34076 15540 34078
rect 15820 34468 15876 34478
rect 15372 34066 15428 34076
rect 15148 33572 15204 33582
rect 15708 33572 15764 33582
rect 15148 33570 15764 33572
rect 15148 33518 15150 33570
rect 15202 33518 15710 33570
rect 15762 33518 15764 33570
rect 15148 33516 15764 33518
rect 15148 33506 15204 33516
rect 15708 33506 15764 33516
rect 14476 33348 14532 33358
rect 14812 33348 14868 33358
rect 14532 33346 14868 33348
rect 14532 33294 14814 33346
rect 14866 33294 14868 33346
rect 14532 33292 14868 33294
rect 14476 33254 14532 33292
rect 14140 33122 14196 33134
rect 14140 33070 14142 33122
rect 14194 33070 14196 33122
rect 14140 33012 14196 33070
rect 13804 32956 14084 33012
rect 14140 32956 14420 33012
rect 12684 32722 12740 32732
rect 13916 32676 13972 32686
rect 10872 32172 11136 32182
rect 10928 32116 10976 32172
rect 11032 32116 11080 32172
rect 10872 32106 11136 32116
rect 13916 31948 13972 32620
rect 13692 31892 13972 31948
rect 8988 31666 9044 31678
rect 8988 31614 8990 31666
rect 9042 31614 9044 31666
rect 8652 31556 8708 31566
rect 5180 31042 5236 31052
rect 8540 31554 8708 31556
rect 8540 31502 8654 31554
rect 8706 31502 8708 31554
rect 8540 31500 8708 31502
rect 8988 31556 9044 31614
rect 9436 31556 9492 31566
rect 8988 31554 9492 31556
rect 8988 31502 9438 31554
rect 9490 31502 9492 31554
rect 8988 31500 9492 31502
rect 8540 30210 8596 31500
rect 8652 31490 8708 31500
rect 9436 31444 9492 31500
rect 9548 31444 9604 31454
rect 9996 31444 10052 31454
rect 9436 31388 9548 31444
rect 9548 31378 9604 31388
rect 9884 31388 9996 31444
rect 9548 31108 9604 31118
rect 9212 31106 9604 31108
rect 9212 31054 9550 31106
rect 9602 31054 9604 31106
rect 9212 31052 9604 31054
rect 9212 30322 9268 31052
rect 9548 31042 9604 31052
rect 9772 30996 9828 31006
rect 9212 30270 9214 30322
rect 9266 30270 9268 30322
rect 9212 30258 9268 30270
rect 9660 30994 9828 30996
rect 9660 30942 9774 30994
rect 9826 30942 9828 30994
rect 9660 30940 9828 30942
rect 8540 30158 8542 30210
rect 8594 30158 8596 30210
rect 5740 30100 5796 30110
rect 5740 29650 5796 30044
rect 5740 29598 5742 29650
rect 5794 29598 5796 29650
rect 5740 29586 5796 29598
rect 5852 29986 5908 29998
rect 5852 29934 5854 29986
rect 5906 29934 5908 29986
rect 4956 29540 5012 29550
rect 4284 27972 4340 27982
rect 4284 27860 4340 27916
rect 4956 27970 5012 29484
rect 5292 29314 5348 29326
rect 5292 29262 5294 29314
rect 5346 29262 5348 29314
rect 5292 29204 5348 29262
rect 5852 29204 5908 29934
rect 6748 29540 6804 29550
rect 6748 29446 6804 29484
rect 7980 29538 8036 29550
rect 7980 29486 7982 29538
rect 8034 29486 8036 29538
rect 6524 29426 6580 29438
rect 6524 29374 6526 29426
rect 6578 29374 6580 29426
rect 6524 29316 6580 29374
rect 6076 29204 6132 29214
rect 5852 29148 6076 29204
rect 5292 29138 5348 29148
rect 6076 29110 6132 29148
rect 4956 27918 4958 27970
rect 5010 27918 5012 27970
rect 4284 27858 4564 27860
rect 4284 27806 4286 27858
rect 4338 27806 4564 27858
rect 4284 27804 4564 27806
rect 4284 27794 4340 27804
rect 4508 27186 4564 27804
rect 4508 27134 4510 27186
rect 4562 27134 4564 27186
rect 4508 27122 4564 27134
rect 4956 26908 5012 27918
rect 5068 28754 5124 28766
rect 5068 28702 5070 28754
rect 5122 28702 5124 28754
rect 5068 27636 5124 28702
rect 5628 28644 5684 28654
rect 5628 28530 5684 28588
rect 5628 28478 5630 28530
rect 5682 28478 5684 28530
rect 5628 28466 5684 28478
rect 5852 28642 5908 28654
rect 5852 28590 5854 28642
rect 5906 28590 5908 28642
rect 5852 28082 5908 28590
rect 5852 28030 5854 28082
rect 5906 28030 5908 28082
rect 5852 28018 5908 28030
rect 5292 27970 5348 27982
rect 5292 27918 5294 27970
rect 5346 27918 5348 27970
rect 5292 27860 5348 27918
rect 5292 27794 5348 27804
rect 6412 27746 6468 27758
rect 6412 27694 6414 27746
rect 6466 27694 6468 27746
rect 5516 27636 5572 27646
rect 6412 27636 6468 27694
rect 5068 27634 6468 27636
rect 5068 27582 5518 27634
rect 5570 27582 6468 27634
rect 5068 27580 6468 27582
rect 5516 27570 5572 27580
rect 4732 26852 5012 26908
rect 4620 26180 4676 26190
rect 4060 26178 4676 26180
rect 4060 26126 4622 26178
rect 4674 26126 4676 26178
rect 4060 26124 4676 26126
rect 4060 24722 4116 26124
rect 4620 26114 4676 26124
rect 4284 25506 4340 25518
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 4284 25284 4340 25454
rect 4284 25218 4340 25228
rect 4060 24670 4062 24722
rect 4114 24670 4116 24722
rect 4060 21812 4116 24670
rect 4732 24836 4788 26852
rect 6076 25396 6132 25406
rect 4844 25284 4900 25294
rect 4844 25190 4900 25228
rect 4284 24164 4340 24174
rect 4284 23938 4340 24108
rect 4284 23886 4286 23938
rect 4338 23886 4340 23938
rect 4284 23874 4340 23886
rect 4620 23044 4676 23054
rect 4060 21746 4116 21756
rect 4172 23042 4676 23044
rect 4172 22990 4622 23042
rect 4674 22990 4676 23042
rect 4172 22988 4676 22990
rect 4172 22370 4228 22988
rect 4620 22978 4676 22988
rect 4172 22318 4174 22370
rect 4226 22318 4228 22370
rect 3388 21644 4004 21700
rect 4172 21700 4228 22318
rect 4732 22258 4788 24780
rect 5516 24836 5572 24846
rect 5516 24742 5572 24780
rect 4844 24722 4900 24734
rect 4844 24670 4846 24722
rect 4898 24670 4900 24722
rect 4844 24612 4900 24670
rect 5852 24724 5908 24734
rect 6076 24724 6132 25340
rect 5852 24722 6132 24724
rect 5852 24670 5854 24722
rect 5906 24670 6132 24722
rect 5852 24668 6132 24670
rect 5852 24658 5908 24668
rect 4844 24546 4900 24556
rect 4844 24164 4900 24174
rect 4844 24050 4900 24108
rect 4844 23998 4846 24050
rect 4898 23998 4900 24050
rect 4844 23986 4900 23998
rect 5740 23940 5796 23950
rect 5740 23846 5796 23884
rect 5740 23380 5796 23390
rect 5740 22482 5796 23324
rect 5740 22430 5742 22482
rect 5794 22430 5796 22482
rect 4956 22372 5012 22382
rect 4956 22278 5012 22316
rect 5740 22372 5796 22430
rect 5796 22316 6020 22372
rect 5740 22306 5796 22316
rect 4732 22206 4734 22258
rect 4786 22206 4788 22258
rect 4732 22194 4788 22206
rect 2380 21588 2436 21598
rect 2268 21586 2436 21588
rect 2268 21534 2382 21586
rect 2434 21534 2436 21586
rect 2268 21532 2436 21534
rect 2380 21522 2436 21532
rect 2828 21586 2884 21598
rect 2828 21534 2830 21586
rect 2882 21534 2884 21586
rect 2828 21364 2884 21534
rect 2156 21308 2884 21364
rect 2716 21028 2772 21038
rect 2716 20934 2772 20972
rect 1820 20750 1822 20802
rect 1874 20750 1876 20802
rect 1820 20738 1876 20750
rect 3164 20132 3220 20142
rect 2716 20130 3220 20132
rect 2716 20078 3166 20130
rect 3218 20078 3220 20130
rect 2716 20076 3220 20078
rect 2716 19346 2772 20076
rect 3164 20066 3220 20076
rect 2716 19294 2718 19346
rect 2770 19294 2772 19346
rect 2716 19282 2772 19294
rect 2044 19236 2100 19246
rect 2044 19234 2212 19236
rect 2044 19182 2046 19234
rect 2098 19182 2212 19234
rect 2044 19180 2212 19182
rect 2044 19170 2100 19180
rect 1932 18676 1988 18686
rect 1932 18338 1988 18620
rect 1932 18286 1934 18338
rect 1986 18286 1988 18338
rect 1932 18274 1988 18286
rect 2156 17668 2212 19180
rect 3388 18452 3444 21644
rect 4172 21634 4228 21644
rect 4956 21812 5012 21822
rect 3612 21476 3668 21486
rect 3612 21474 4676 21476
rect 3612 21422 3614 21474
rect 3666 21422 4676 21474
rect 3612 21420 4676 21422
rect 3612 21410 3668 21420
rect 4620 20690 4676 21420
rect 4956 20916 5012 21756
rect 4956 20850 5012 20860
rect 5740 21474 5796 21486
rect 5740 21422 5742 21474
rect 5794 21422 5796 21474
rect 5740 20804 5796 21422
rect 5740 20738 5796 20748
rect 4620 20638 4622 20690
rect 4674 20638 4676 20690
rect 4620 20626 4676 20638
rect 4956 20692 5012 20702
rect 4956 20598 5012 20636
rect 5852 20692 5908 20702
rect 5852 20598 5908 20636
rect 3500 20132 3556 20142
rect 3500 20130 4788 20132
rect 3500 20078 3502 20130
rect 3554 20078 4788 20130
rect 3500 20076 4788 20078
rect 3500 20066 3556 20076
rect 3948 19908 4004 19918
rect 4396 19908 4452 19918
rect 3948 19906 4452 19908
rect 3948 19854 3950 19906
rect 4002 19854 4398 19906
rect 4450 19854 4452 19906
rect 3948 19852 4452 19854
rect 3948 19842 4004 19852
rect 3836 19794 3892 19806
rect 3836 19742 3838 19794
rect 3890 19742 3892 19794
rect 3836 18676 3892 19742
rect 4396 19796 4452 19852
rect 4396 19730 4452 19740
rect 3836 18620 4004 18676
rect 3836 18452 3892 18462
rect 3388 18450 3892 18452
rect 3388 18398 3838 18450
rect 3890 18398 3892 18450
rect 3388 18396 3892 18398
rect 2044 17666 2212 17668
rect 2044 17614 2158 17666
rect 2210 17614 2212 17666
rect 2044 17612 2212 17614
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 1932 16146 1988 16156
rect 2044 15316 2100 17612
rect 2156 17602 2212 17612
rect 2940 17556 2996 17566
rect 2940 17554 3332 17556
rect 2940 17502 2942 17554
rect 2994 17502 3332 17554
rect 2940 17500 3332 17502
rect 2940 17490 2996 17500
rect 3276 15988 3332 17500
rect 3836 17108 3892 18396
rect 3836 17042 3892 17052
rect 3948 16882 4004 18620
rect 4732 18674 4788 20076
rect 4732 18622 4734 18674
rect 4786 18622 4788 18674
rect 4732 18610 4788 18622
rect 4844 19346 4900 19358
rect 4844 19294 4846 19346
rect 4898 19294 4900 19346
rect 4844 18228 4900 19294
rect 5404 19348 5460 19358
rect 5068 18228 5124 18238
rect 4844 18226 5236 18228
rect 4844 18174 5070 18226
rect 5122 18174 5236 18226
rect 4844 18172 5236 18174
rect 5068 18162 5124 18172
rect 5068 17780 5124 17790
rect 5068 17686 5124 17724
rect 5180 17668 5236 18172
rect 5292 17668 5348 17678
rect 5180 17612 5292 17668
rect 5292 17602 5348 17612
rect 4732 17108 4788 17118
rect 4788 17052 4900 17108
rect 4732 17042 4788 17052
rect 4844 16994 4900 17052
rect 4844 16942 4846 16994
rect 4898 16942 4900 16994
rect 4844 16930 4900 16942
rect 3948 16830 3950 16882
rect 4002 16830 4004 16882
rect 3948 16818 4004 16830
rect 3724 16100 3780 16110
rect 3724 16006 3780 16044
rect 3388 15988 3444 15998
rect 3276 15986 3444 15988
rect 3276 15934 3390 15986
rect 3442 15934 3444 15986
rect 3276 15932 3444 15934
rect 3388 15922 3444 15932
rect 4396 15988 4452 15998
rect 4396 15894 4452 15932
rect 5292 15988 5348 15998
rect 2716 15876 2772 15886
rect 2716 15426 2772 15820
rect 4060 15876 4116 15886
rect 4060 15782 4116 15820
rect 5292 15538 5348 15932
rect 5292 15486 5294 15538
rect 5346 15486 5348 15538
rect 5292 15474 5348 15486
rect 2716 15374 2718 15426
rect 2770 15374 2772 15426
rect 2716 15362 2772 15374
rect 4844 15316 4900 15326
rect 2044 15314 2212 15316
rect 2044 15262 2046 15314
rect 2098 15262 2212 15314
rect 2044 15260 2212 15262
rect 2044 15250 2100 15260
rect 1932 14642 1988 14654
rect 1932 14590 1934 14642
rect 1986 14590 1988 14642
rect 1932 13748 1988 14590
rect 1932 13682 1988 13692
rect 2156 13748 2212 15260
rect 4844 15202 4900 15260
rect 4844 15150 4846 15202
rect 4898 15150 4900 15202
rect 4844 15138 4900 15150
rect 5404 15148 5460 19292
rect 5852 18562 5908 18574
rect 5852 18510 5854 18562
rect 5906 18510 5908 18562
rect 5740 18452 5796 18462
rect 5740 18358 5796 18396
rect 5852 17556 5908 18510
rect 5852 17490 5908 17500
rect 5740 17442 5796 17454
rect 5740 17390 5742 17442
rect 5794 17390 5796 17442
rect 5628 16212 5684 16222
rect 5628 15316 5684 16156
rect 5740 16100 5796 17390
rect 5740 16034 5796 16044
rect 5964 15540 6020 22316
rect 6076 21028 6132 24668
rect 6188 24612 6244 24622
rect 6300 24612 6356 24622
rect 6244 24610 6356 24612
rect 6244 24558 6302 24610
rect 6354 24558 6356 24610
rect 6244 24556 6356 24558
rect 6188 22036 6244 24556
rect 6300 24546 6356 24556
rect 6412 24388 6468 27580
rect 6300 24332 6468 24388
rect 6300 22260 6356 24332
rect 6524 24052 6580 29260
rect 7420 29316 7476 29326
rect 7420 29222 7476 29260
rect 6748 29204 6804 29214
rect 6748 27860 6804 29148
rect 7084 28756 7140 28766
rect 7084 28642 7140 28700
rect 7868 28756 7924 28766
rect 7980 28756 8036 29486
rect 7868 28754 8036 28756
rect 7868 28702 7870 28754
rect 7922 28702 8036 28754
rect 7868 28700 8036 28702
rect 8316 29426 8372 29438
rect 8316 29374 8318 29426
rect 8370 29374 8372 29426
rect 7868 28690 7924 28700
rect 7084 28590 7086 28642
rect 7138 28590 7140 28642
rect 7084 28578 7140 28590
rect 8316 28084 8372 29374
rect 8540 29428 8596 30158
rect 9660 29650 9716 30940
rect 9772 30930 9828 30940
rect 9660 29598 9662 29650
rect 9714 29598 9716 29650
rect 9660 29586 9716 29598
rect 8540 29362 8596 29372
rect 8316 28018 8372 28028
rect 9660 28084 9716 28094
rect 9660 27990 9716 28028
rect 6748 27794 6804 27804
rect 6860 27748 6916 27758
rect 6916 27692 7028 27748
rect 6860 27654 6916 27692
rect 6748 27076 6804 27086
rect 6748 26982 6804 27020
rect 6300 22194 6356 22204
rect 6412 23996 6580 24052
rect 6188 21980 6356 22036
rect 6188 21812 6244 21822
rect 6188 21586 6244 21756
rect 6188 21534 6190 21586
rect 6242 21534 6244 21586
rect 6188 21522 6244 21534
rect 6188 21028 6244 21038
rect 6076 21026 6244 21028
rect 6076 20974 6190 21026
rect 6242 20974 6244 21026
rect 6076 20972 6244 20974
rect 6188 20962 6244 20972
rect 6300 18228 6356 21980
rect 6412 18452 6468 23996
rect 6524 23828 6580 23838
rect 6524 23826 6692 23828
rect 6524 23774 6526 23826
rect 6578 23774 6692 23826
rect 6524 23772 6692 23774
rect 6524 23762 6580 23772
rect 6636 23380 6692 23772
rect 6860 23380 6916 23390
rect 6636 23378 6916 23380
rect 6636 23326 6862 23378
rect 6914 23326 6916 23378
rect 6636 23324 6916 23326
rect 6860 23314 6916 23324
rect 6972 21700 7028 27692
rect 9548 27186 9604 27198
rect 9548 27134 9550 27186
rect 9602 27134 9604 27186
rect 7420 26962 7476 26974
rect 7420 26910 7422 26962
rect 7474 26910 7476 26962
rect 7308 26516 7364 26526
rect 7420 26516 7476 26910
rect 7308 26514 7476 26516
rect 7308 26462 7310 26514
rect 7362 26462 7476 26514
rect 7308 26460 7476 26462
rect 7308 26450 7364 26460
rect 8428 26402 8484 26414
rect 8428 26350 8430 26402
rect 8482 26350 8484 26402
rect 7084 26292 7140 26302
rect 7756 26292 7812 26302
rect 7084 26290 7812 26292
rect 7084 26238 7086 26290
rect 7138 26238 7758 26290
rect 7810 26238 7812 26290
rect 7084 26236 7812 26238
rect 7084 26226 7140 26236
rect 7756 26226 7812 26236
rect 8092 26292 8148 26302
rect 8092 26198 8148 26236
rect 8428 25172 8484 26350
rect 8876 26404 8932 26414
rect 8876 26310 8932 26348
rect 9548 26292 9604 27134
rect 9884 26740 9940 31388
rect 9996 31378 10052 31388
rect 10872 30604 11136 30614
rect 10928 30548 10976 30604
rect 11032 30548 11080 30604
rect 10872 30538 11136 30548
rect 11340 30322 11396 30334
rect 11340 30270 11342 30322
rect 11394 30270 11396 30322
rect 10220 29538 10276 29550
rect 10220 29486 10222 29538
rect 10274 29486 10276 29538
rect 9996 29428 10052 29438
rect 9996 29334 10052 29372
rect 10220 29316 10276 29486
rect 10220 29250 10276 29260
rect 10556 29538 10612 29550
rect 10556 29486 10558 29538
rect 10610 29486 10612 29538
rect 9996 28754 10052 28766
rect 9996 28702 9998 28754
rect 10050 28702 10052 28754
rect 9996 27636 10052 28702
rect 10220 27970 10276 27982
rect 10220 27918 10222 27970
rect 10274 27918 10276 27970
rect 10220 27748 10276 27918
rect 10220 27682 10276 27692
rect 10556 27970 10612 29486
rect 11340 29428 11396 30270
rect 13132 30212 13188 30222
rect 13132 29538 13188 30156
rect 13132 29486 13134 29538
rect 13186 29486 13188 29538
rect 13132 29474 13188 29486
rect 13244 29540 13300 29550
rect 13244 29538 13636 29540
rect 13244 29486 13246 29538
rect 13298 29486 13636 29538
rect 13244 29484 13636 29486
rect 13244 29474 13300 29484
rect 11340 29314 11396 29372
rect 11340 29262 11342 29314
rect 11394 29262 11396 29314
rect 10872 29036 11136 29046
rect 10928 28980 10976 29036
rect 11032 28980 11080 29036
rect 10872 28970 11136 28980
rect 10556 27918 10558 27970
rect 10610 27918 10612 27970
rect 9996 27542 10052 27580
rect 9884 26674 9940 26684
rect 10108 27076 10164 27086
rect 9548 26226 9604 26236
rect 9884 26404 9940 26414
rect 8428 24612 8484 25116
rect 9660 26178 9716 26190
rect 9660 26126 9662 26178
rect 9714 26126 9716 26178
rect 9660 25172 9716 26126
rect 9660 25106 9716 25116
rect 8428 24546 8484 24556
rect 9548 24948 9604 24958
rect 9548 24722 9604 24892
rect 9548 24670 9550 24722
rect 9602 24670 9604 24722
rect 8652 24050 8708 24062
rect 8652 23998 8654 24050
rect 8706 23998 8708 24050
rect 8652 23940 8708 23998
rect 9436 23940 9492 23950
rect 8652 23938 9492 23940
rect 8652 23886 9438 23938
rect 9490 23886 9492 23938
rect 8652 23884 9492 23886
rect 9100 23714 9156 23726
rect 9100 23662 9102 23714
rect 9154 23662 9156 23714
rect 8652 23380 8708 23390
rect 8652 23286 8708 23324
rect 7196 23268 7252 23278
rect 7196 23174 7252 23212
rect 9100 23268 9156 23662
rect 9100 23202 9156 23212
rect 6748 21644 7028 21700
rect 8652 23044 8708 23054
rect 6748 21028 6804 21644
rect 6860 21476 6916 21486
rect 6860 21474 7812 21476
rect 6860 21422 6862 21474
rect 6914 21422 7812 21474
rect 6860 21420 7812 21422
rect 6860 21410 6916 21420
rect 6748 20972 7476 21028
rect 6972 20804 7028 20814
rect 6972 20802 7364 20804
rect 6972 20750 6974 20802
rect 7026 20750 7364 20802
rect 6972 20748 7364 20750
rect 6972 20738 7028 20748
rect 6860 20692 6916 20702
rect 6860 20598 6916 20636
rect 7308 20132 7364 20748
rect 7308 20038 7364 20076
rect 6412 18358 6468 18396
rect 6300 18172 6804 18228
rect 6076 17780 6132 17790
rect 6076 17686 6132 17724
rect 6748 17666 6804 18172
rect 6748 17614 6750 17666
rect 6802 17614 6804 17666
rect 6636 17556 6692 17566
rect 6412 17500 6636 17556
rect 6188 16882 6244 16894
rect 6188 16830 6190 16882
rect 6242 16830 6244 16882
rect 6188 15988 6244 16830
rect 6188 15922 6244 15932
rect 5964 15426 6020 15484
rect 5964 15374 5966 15426
rect 6018 15374 6020 15426
rect 5964 15362 6020 15374
rect 6412 15428 6468 17500
rect 6636 17462 6692 17500
rect 6748 17444 6804 17614
rect 7308 17444 7364 17454
rect 6748 17378 6804 17388
rect 6860 17442 7364 17444
rect 6860 17390 7310 17442
rect 7362 17390 7364 17442
rect 6860 17388 7364 17390
rect 6860 16994 6916 17388
rect 7308 17378 7364 17388
rect 6860 16942 6862 16994
rect 6914 16942 6916 16994
rect 6860 16930 6916 16942
rect 6860 15428 6916 15438
rect 6412 15426 6916 15428
rect 6412 15374 6414 15426
rect 6466 15374 6862 15426
rect 6914 15374 6916 15426
rect 6412 15372 6916 15374
rect 6412 15362 6468 15372
rect 5628 15222 5684 15260
rect 5180 15092 5460 15148
rect 4284 14532 4340 14542
rect 4284 14530 4452 14532
rect 4284 14478 4286 14530
rect 4338 14478 4452 14530
rect 4284 14476 4452 14478
rect 4284 14466 4340 14476
rect 4396 14308 4452 14476
rect 4844 14308 4900 14318
rect 4396 14306 4900 14308
rect 4396 14254 4846 14306
rect 4898 14254 4900 14306
rect 4396 14252 4900 14254
rect 2156 13746 2436 13748
rect 2156 13694 2158 13746
rect 2210 13694 2436 13746
rect 2156 13692 2436 13694
rect 2156 13682 2212 13692
rect 2380 12850 2436 13692
rect 2940 13636 2996 13646
rect 2940 13634 3332 13636
rect 2940 13582 2942 13634
rect 2994 13582 3332 13634
rect 2940 13580 3332 13582
rect 2940 13570 2996 13580
rect 2716 13076 2772 13086
rect 2716 12964 2772 13020
rect 2716 12962 2996 12964
rect 2716 12910 2718 12962
rect 2770 12910 2996 12962
rect 2716 12908 2996 12910
rect 2716 12898 2772 12908
rect 2380 12798 2382 12850
rect 2434 12798 2436 12850
rect 2380 12786 2436 12798
rect 2828 12292 2884 12302
rect 2492 12290 2884 12292
rect 2492 12238 2830 12290
rect 2882 12238 2884 12290
rect 2492 12236 2884 12238
rect 1820 12180 1876 12190
rect 1820 11394 1876 12124
rect 2492 11506 2548 12236
rect 2828 12226 2884 12236
rect 2492 11454 2494 11506
rect 2546 11454 2548 11506
rect 2492 11442 2548 11454
rect 1820 11342 1822 11394
rect 1874 11342 1876 11394
rect 1820 8428 1876 11342
rect 1932 11284 1988 11294
rect 1932 10498 1988 11228
rect 1932 10446 1934 10498
rect 1986 10446 1988 10498
rect 1932 10434 1988 10446
rect 2828 9604 2884 9614
rect 2492 9602 2884 9604
rect 2492 9550 2830 9602
rect 2882 9550 2884 9602
rect 2492 9548 2884 9550
rect 1932 8820 1988 8830
rect 1932 8726 1988 8764
rect 1708 8372 1876 8428
rect 1708 8260 1764 8372
rect 2492 8370 2548 9548
rect 2828 9538 2884 9548
rect 2940 8428 2996 12908
rect 3276 12850 3332 13580
rect 3612 12964 3668 12974
rect 3612 12870 3668 12908
rect 3276 12798 3278 12850
rect 3330 12798 3332 12850
rect 3276 12786 3332 12798
rect 3164 12178 3220 12190
rect 3164 12126 3166 12178
rect 3218 12126 3220 12178
rect 3164 10836 3220 12126
rect 3164 10770 3220 10780
rect 4284 11508 4340 11518
rect 4284 10610 4340 11452
rect 4284 10558 4286 10610
rect 4338 10558 4340 10610
rect 4284 10546 4340 10558
rect 4172 9828 4228 9838
rect 4172 9734 4228 9772
rect 3164 9716 3220 9726
rect 3164 9622 3220 9660
rect 3836 9716 3892 9726
rect 3836 9622 3892 9660
rect 4284 9268 4340 9278
rect 4284 9042 4340 9212
rect 4284 8990 4286 9042
rect 4338 8990 4340 9042
rect 4284 8978 4340 8990
rect 2492 8318 2494 8370
rect 2546 8318 2548 8370
rect 2492 8306 2548 8318
rect 2716 8372 2996 8428
rect 1820 8260 1876 8270
rect 1708 8258 1876 8260
rect 1708 8206 1822 8258
rect 1874 8206 1876 8258
rect 1708 8204 1876 8206
rect 1820 7588 1876 8204
rect 2716 7700 2772 8372
rect 2380 7588 2436 7598
rect 1820 7586 2436 7588
rect 1820 7534 2382 7586
rect 2434 7534 2436 7586
rect 1820 7532 2436 7534
rect 2380 7364 2436 7532
rect 2716 7586 2772 7644
rect 2716 7534 2718 7586
rect 2770 7534 2772 7586
rect 2716 7522 2772 7534
rect 3836 8036 3892 8046
rect 3836 7586 3892 7980
rect 3836 7534 3838 7586
rect 3890 7534 3892 7586
rect 3836 7522 3892 7534
rect 3052 7476 3108 7486
rect 2940 7474 3108 7476
rect 2940 7422 3054 7474
rect 3106 7422 3108 7474
rect 2940 7420 3108 7422
rect 2940 7364 2996 7420
rect 3052 7410 3108 7420
rect 2380 7308 2996 7364
rect 4284 6692 4340 6702
rect 4284 6598 4340 6636
rect 2492 6580 2548 6590
rect 2492 6486 2548 6524
rect 4396 5012 4452 14252
rect 4844 14242 4900 14252
rect 5068 14308 5124 14318
rect 4844 13972 4900 13982
rect 4620 11506 4676 11518
rect 4620 11454 4622 11506
rect 4674 11454 4676 11506
rect 4620 10388 4676 11454
rect 4732 10836 4788 10846
rect 4732 10742 4788 10780
rect 4620 10322 4676 10332
rect 4732 9940 4788 9950
rect 4620 9828 4676 9838
rect 4620 8370 4676 9772
rect 4732 9826 4788 9884
rect 4732 9774 4734 9826
rect 4786 9774 4788 9826
rect 4732 9762 4788 9774
rect 4844 9492 4900 13916
rect 5068 13634 5124 14252
rect 5068 13582 5070 13634
rect 5122 13582 5124 13634
rect 5068 13570 5124 13582
rect 5068 11508 5124 11518
rect 5180 11508 5236 15092
rect 6076 14530 6132 14542
rect 6076 14478 6078 14530
rect 6130 14478 6132 14530
rect 5740 14306 5796 14318
rect 5740 14254 5742 14306
rect 5794 14254 5796 14306
rect 5740 12964 5796 14254
rect 6076 14308 6132 14478
rect 6748 14418 6804 15372
rect 6860 15362 6916 15372
rect 7196 15314 7252 15326
rect 7196 15262 7198 15314
rect 7250 15262 7252 15314
rect 7196 15092 7252 15262
rect 7196 15026 7252 15036
rect 6860 14532 6916 14542
rect 7420 14532 7476 20972
rect 7756 20690 7812 21420
rect 7980 20804 8036 20814
rect 7756 20638 7758 20690
rect 7810 20638 7812 20690
rect 7756 20626 7812 20638
rect 7868 20802 8036 20804
rect 7868 20750 7982 20802
rect 8034 20750 8036 20802
rect 7868 20748 8036 20750
rect 7756 20244 7812 20254
rect 7868 20244 7924 20748
rect 7980 20738 8036 20748
rect 7756 20242 7924 20244
rect 7756 20190 7758 20242
rect 7810 20190 7924 20242
rect 7756 20188 7924 20190
rect 7756 20178 7812 20188
rect 8540 20132 8596 20142
rect 8092 20020 8148 20030
rect 8092 19926 8148 19964
rect 7532 18452 7588 18462
rect 7532 16212 7588 18396
rect 7644 17556 7700 17566
rect 7644 17554 7812 17556
rect 7644 17502 7646 17554
rect 7698 17502 7812 17554
rect 7644 17500 7812 17502
rect 7644 17490 7700 17500
rect 7756 16322 7812 17500
rect 7756 16270 7758 16322
rect 7810 16270 7812 16322
rect 7756 16258 7812 16270
rect 7980 17444 8036 17454
rect 8092 17444 8148 17454
rect 8036 17442 8148 17444
rect 8036 17390 8094 17442
rect 8146 17390 8148 17442
rect 8036 17388 8148 17390
rect 7532 16156 7700 16212
rect 7644 16100 7700 16156
rect 7644 16044 7812 16100
rect 6860 14530 7476 14532
rect 6860 14478 6862 14530
rect 6914 14478 7476 14530
rect 6860 14476 7476 14478
rect 7532 15988 7588 15998
rect 6860 14466 6916 14476
rect 6748 14366 6750 14418
rect 6802 14366 6804 14418
rect 6748 14354 6804 14366
rect 6076 14242 6132 14252
rect 5740 12898 5796 12908
rect 7084 13636 7140 14476
rect 7532 14308 7588 15932
rect 7420 14306 7588 14308
rect 7420 14254 7534 14306
rect 7586 14254 7588 14306
rect 7420 14252 7588 14254
rect 7196 13636 7252 13646
rect 7084 13634 7252 13636
rect 7084 13582 7198 13634
rect 7250 13582 7252 13634
rect 7084 13580 7252 13582
rect 6524 12850 6580 12862
rect 6524 12798 6526 12850
rect 6578 12798 6580 12850
rect 6188 12740 6244 12750
rect 6188 12738 6356 12740
rect 6188 12686 6190 12738
rect 6242 12686 6356 12738
rect 6188 12684 6356 12686
rect 6188 12674 6244 12684
rect 6300 12290 6356 12684
rect 6300 12238 6302 12290
rect 6354 12238 6356 12290
rect 6300 12226 6356 12238
rect 5516 12180 5572 12190
rect 5516 12086 5572 12124
rect 6524 11620 6580 12798
rect 6636 11620 6692 11630
rect 6524 11618 6692 11620
rect 6524 11566 6638 11618
rect 6690 11566 6692 11618
rect 6524 11564 6692 11566
rect 6636 11554 6692 11564
rect 5124 11452 5236 11508
rect 6972 11508 7028 11518
rect 5068 11414 5124 11452
rect 6972 11414 7028 11452
rect 6188 10836 6244 10846
rect 5180 10724 5236 10734
rect 5068 10388 5124 10398
rect 5068 10052 5124 10332
rect 5068 9986 5124 9996
rect 4956 9716 5012 9726
rect 5180 9716 5236 10668
rect 5852 10724 5908 10734
rect 5852 10630 5908 10668
rect 5628 10612 5684 10622
rect 5628 10518 5684 10556
rect 6188 9940 6244 10780
rect 6972 10612 7028 10622
rect 7084 10612 7140 13580
rect 7196 13570 7252 13580
rect 7420 12962 7476 14252
rect 7532 14242 7588 14252
rect 7644 15540 7700 15550
rect 7420 12910 7422 12962
rect 7474 12910 7476 12962
rect 7420 12898 7476 12910
rect 7644 11508 7700 15484
rect 7028 10556 7140 10612
rect 7308 11452 7700 11508
rect 6412 10498 6468 10510
rect 6412 10446 6414 10498
rect 6466 10446 6468 10498
rect 6412 10052 6468 10446
rect 6412 9986 6468 9996
rect 6636 10500 6692 10510
rect 6188 9846 6244 9884
rect 5740 9828 5796 9838
rect 5740 9734 5796 9772
rect 4956 9714 5236 9716
rect 4956 9662 4958 9714
rect 5010 9662 5236 9714
rect 4956 9660 5236 9662
rect 4956 9650 5012 9660
rect 4844 9436 5012 9492
rect 4620 8318 4622 8370
rect 4674 8318 4676 8370
rect 4620 8306 4676 8318
rect 4844 6692 4900 6702
rect 4844 6598 4900 6636
rect 4396 4946 4452 4956
rect 4284 4338 4340 4350
rect 4284 4286 4286 4338
rect 4338 4286 4340 4338
rect 1932 4116 1988 4126
rect 1932 4022 1988 4060
rect 4284 3780 4340 4286
rect 4284 3714 4340 3724
rect 4732 4226 4788 4238
rect 4732 4174 4734 4226
rect 4786 4174 4788 4226
rect 1932 3666 1988 3678
rect 1932 3614 1934 3666
rect 1986 3614 1988 3666
rect 1932 1540 1988 3614
rect 4284 3556 4340 3566
rect 4284 3462 4340 3500
rect 4732 3554 4788 4174
rect 4732 3502 4734 3554
rect 4786 3502 4788 3554
rect 4732 3388 4788 3502
rect 1932 1474 1988 1484
rect 4620 3332 4788 3388
rect 4956 3442 5012 9436
rect 5180 9154 5236 9660
rect 5180 9102 5182 9154
rect 5234 9102 5236 9154
rect 5180 9090 5236 9102
rect 5292 9268 5348 9278
rect 6636 9268 6692 10444
rect 5180 8372 5236 8382
rect 5292 8372 5348 9212
rect 5740 9266 6692 9268
rect 5740 9214 6638 9266
rect 6690 9214 6692 9266
rect 5740 9212 6692 9214
rect 5516 9156 5572 9166
rect 5516 9062 5572 9100
rect 5740 9042 5796 9212
rect 5740 8990 5742 9042
rect 5794 8990 5796 9042
rect 5740 8978 5796 8990
rect 5180 8370 5348 8372
rect 5180 8318 5182 8370
rect 5234 8318 5348 8370
rect 5180 8316 5348 8318
rect 5180 8306 5236 8316
rect 5628 8036 5684 8046
rect 5628 7942 5684 7980
rect 5852 7364 5908 9212
rect 6636 9202 6692 9212
rect 6972 10498 7028 10556
rect 7308 10500 7364 11452
rect 7756 11394 7812 16044
rect 7868 14418 7924 14430
rect 7868 14366 7870 14418
rect 7922 14366 7924 14418
rect 7868 13076 7924 14366
rect 7868 13010 7924 13020
rect 7756 11342 7758 11394
rect 7810 11342 7812 11394
rect 6972 10446 6974 10498
rect 7026 10446 7028 10498
rect 6076 8820 6132 8830
rect 5964 8818 6132 8820
rect 5964 8766 6078 8818
rect 6130 8766 6132 8818
rect 5964 8764 6132 8766
rect 5964 8258 6020 8764
rect 6076 8754 6132 8764
rect 5964 8206 5966 8258
rect 6018 8206 6020 8258
rect 5964 8194 6020 8206
rect 5964 7364 6020 7374
rect 5852 7362 6020 7364
rect 5852 7310 5966 7362
rect 6018 7310 6020 7362
rect 5852 7308 6020 7310
rect 5964 7298 6020 7308
rect 6076 7364 6132 7374
rect 6076 5794 6132 7308
rect 6076 5742 6078 5794
rect 6130 5742 6132 5794
rect 6076 5730 6132 5742
rect 5180 4226 5236 4238
rect 5180 4174 5182 4226
rect 5234 4174 5236 4226
rect 5180 3780 5236 4174
rect 5180 3714 5236 3724
rect 5740 4116 5796 4126
rect 5740 3666 5796 4060
rect 5740 3614 5742 3666
rect 5794 3614 5796 3666
rect 5740 3556 5796 3614
rect 5740 3490 5796 3500
rect 4956 3390 4958 3442
rect 5010 3390 5012 3442
rect 4956 3378 5012 3390
rect 3612 924 4004 980
rect 3612 800 3668 924
rect 3584 0 3696 800
rect 3948 756 4004 924
rect 4620 756 4676 3332
rect 6972 2436 7028 10446
rect 7084 10444 7364 10500
rect 7532 11282 7588 11294
rect 7532 11230 7534 11282
rect 7586 11230 7588 11282
rect 7532 10724 7588 11230
rect 7756 11172 7812 11342
rect 7756 11106 7812 11116
rect 7084 9266 7140 10444
rect 7084 9214 7086 9266
rect 7138 9214 7140 9266
rect 7084 9156 7140 9214
rect 7084 9090 7140 9100
rect 7420 9938 7476 9950
rect 7420 9886 7422 9938
rect 7474 9886 7476 9938
rect 7420 8820 7476 9886
rect 7532 9266 7588 10668
rect 7980 10724 8036 17388
rect 8092 17378 8148 17388
rect 8092 16098 8148 16110
rect 8092 16046 8094 16098
rect 8146 16046 8148 16098
rect 8092 15092 8148 16046
rect 8540 16100 8596 20076
rect 8540 16006 8596 16044
rect 8092 15026 8148 15036
rect 8652 13972 8708 22988
rect 9436 21588 9492 23884
rect 9436 21522 9492 21532
rect 8988 21476 9044 21486
rect 8764 21420 8988 21476
rect 8764 20130 8820 21420
rect 8988 21382 9044 21420
rect 8764 20078 8766 20130
rect 8818 20078 8820 20130
rect 8764 20066 8820 20078
rect 8876 20018 8932 20030
rect 8876 19966 8878 20018
rect 8930 19966 8932 20018
rect 8876 19012 8932 19966
rect 9548 20020 9604 24670
rect 9884 24946 9940 26348
rect 9884 24894 9886 24946
rect 9938 24894 9940 24946
rect 9660 23826 9716 23838
rect 9660 23774 9662 23826
rect 9714 23774 9716 23826
rect 9660 23380 9716 23774
rect 9884 23828 9940 24894
rect 10108 24724 10164 27020
rect 10556 26404 10612 27918
rect 10668 28756 10724 28766
rect 10668 26908 10724 28700
rect 11340 28644 11396 29262
rect 11788 29316 11844 29326
rect 11788 29222 11844 29260
rect 13244 29204 13300 29214
rect 13244 29110 13300 29148
rect 13580 28868 13636 29484
rect 13692 29426 13748 31892
rect 13692 29374 13694 29426
rect 13746 29374 13748 29426
rect 13692 29362 13748 29374
rect 13804 30100 13860 30110
rect 13692 28868 13748 28878
rect 13580 28866 13748 28868
rect 13580 28814 13694 28866
rect 13746 28814 13748 28866
rect 13580 28812 13748 28814
rect 13692 28802 13748 28812
rect 13804 28754 13860 30044
rect 13804 28702 13806 28754
rect 13858 28702 13860 28754
rect 13804 28690 13860 28702
rect 11340 28578 11396 28588
rect 11228 28420 11284 28430
rect 11116 28418 11284 28420
rect 11116 28366 11230 28418
rect 11282 28366 11284 28418
rect 11116 28364 11284 28366
rect 11004 27748 11060 27758
rect 11116 27748 11172 28364
rect 11228 28354 11284 28364
rect 11340 27972 11396 27982
rect 11060 27692 11172 27748
rect 11228 27970 11396 27972
rect 11228 27918 11342 27970
rect 11394 27918 11396 27970
rect 11228 27916 11396 27918
rect 11004 27682 11060 27692
rect 10872 27468 11136 27478
rect 10928 27412 10976 27468
rect 11032 27412 11080 27468
rect 10872 27402 11136 27412
rect 11228 27300 11284 27916
rect 11340 27906 11396 27916
rect 10780 27244 11284 27300
rect 11676 27858 11732 27870
rect 11676 27806 11678 27858
rect 11730 27806 11732 27858
rect 10780 27186 10836 27244
rect 10780 27134 10782 27186
rect 10834 27134 10836 27186
rect 10780 27122 10836 27134
rect 10668 26852 11060 26908
rect 11004 26516 11060 26852
rect 11228 26740 11284 26750
rect 11284 26684 11396 26740
rect 11228 26674 11284 26684
rect 11004 26514 11284 26516
rect 11004 26462 11006 26514
rect 11058 26462 11284 26514
rect 11004 26460 11284 26462
rect 11004 26450 11060 26460
rect 10556 26338 10612 26348
rect 10872 25900 11136 25910
rect 10928 25844 10976 25900
rect 11032 25844 11080 25900
rect 10872 25834 11136 25844
rect 11116 25508 11172 25518
rect 11228 25508 11284 26460
rect 11340 26514 11396 26684
rect 11340 26462 11342 26514
rect 11394 26462 11396 26514
rect 11340 26450 11396 26462
rect 11116 25506 11284 25508
rect 11116 25454 11118 25506
rect 11170 25454 11284 25506
rect 11116 25452 11284 25454
rect 11564 26292 11620 26302
rect 11116 25442 11172 25452
rect 10220 25282 10276 25294
rect 10220 25230 10222 25282
rect 10274 25230 10276 25282
rect 10220 24948 10276 25230
rect 10220 24882 10276 24892
rect 10780 25282 10836 25294
rect 10780 25230 10782 25282
rect 10834 25230 10836 25282
rect 10556 24724 10612 24734
rect 10780 24724 10836 25230
rect 10108 24722 10836 24724
rect 10108 24670 10558 24722
rect 10610 24670 10836 24722
rect 10108 24668 10836 24670
rect 9996 23828 10052 23838
rect 9884 23826 10052 23828
rect 9884 23774 9998 23826
rect 10050 23774 10052 23826
rect 9884 23772 10052 23774
rect 9996 23762 10052 23772
rect 9660 23314 9716 23324
rect 10220 22932 10276 22942
rect 9996 21700 10052 21710
rect 9884 21588 9940 21598
rect 9884 20132 9940 21532
rect 9996 20804 10052 21644
rect 9996 20710 10052 20748
rect 10108 20580 10164 20590
rect 10108 20486 10164 20524
rect 9996 20132 10052 20142
rect 9884 20130 10052 20132
rect 9884 20078 9998 20130
rect 10050 20078 10052 20130
rect 9884 20076 10052 20078
rect 9996 20066 10052 20076
rect 9660 20020 9716 20030
rect 9548 19964 9660 20020
rect 9660 19926 9716 19964
rect 10108 20020 10164 20030
rect 10108 19926 10164 19964
rect 10108 19124 10164 19134
rect 9212 19012 9268 19022
rect 8876 19010 9268 19012
rect 8876 18958 9214 19010
rect 9266 18958 9268 19010
rect 8876 18956 9268 18958
rect 8988 16772 9044 16782
rect 8876 15988 8932 15998
rect 8988 15988 9044 16716
rect 8876 15986 9044 15988
rect 8876 15934 8878 15986
rect 8930 15934 9044 15986
rect 8876 15932 9044 15934
rect 8876 15922 8932 15932
rect 9212 15148 9268 18956
rect 9436 16210 9492 16222
rect 9436 16158 9438 16210
rect 9490 16158 9492 16210
rect 9324 16100 9380 16110
rect 9436 16100 9492 16158
rect 9380 16044 9940 16100
rect 9324 16034 9380 16044
rect 9212 15092 9828 15148
rect 8652 13906 8708 13916
rect 8428 13858 8484 13870
rect 8428 13806 8430 13858
rect 8482 13806 8484 13858
rect 8092 13076 8148 13086
rect 8428 13076 8484 13806
rect 8652 13748 8708 13758
rect 8092 13074 8484 13076
rect 8092 13022 8094 13074
rect 8146 13022 8484 13074
rect 8092 13020 8484 13022
rect 8540 13692 8652 13748
rect 8092 13010 8148 13020
rect 8428 12068 8484 12078
rect 8540 12068 8596 13692
rect 8652 13682 8708 13692
rect 8764 13748 8820 13758
rect 9660 13748 9716 13758
rect 8764 13746 9716 13748
rect 8764 13694 8766 13746
rect 8818 13694 9662 13746
rect 9714 13694 9716 13746
rect 8764 13692 9716 13694
rect 8764 13682 8820 13692
rect 9660 13682 9716 13692
rect 8428 12066 8596 12068
rect 8428 12014 8430 12066
rect 8482 12014 8596 12066
rect 8428 12012 8596 12014
rect 8316 11508 8372 11518
rect 8428 11508 8484 12012
rect 8372 11452 8484 11508
rect 8316 11414 8372 11452
rect 8764 11172 8820 11182
rect 8764 11078 8820 11116
rect 7980 10658 8036 10668
rect 8876 10724 8932 10734
rect 9548 10724 9604 10734
rect 8876 10722 9492 10724
rect 8876 10670 8878 10722
rect 8930 10670 9492 10722
rect 8876 10668 9492 10670
rect 8876 10658 8932 10668
rect 8652 10612 8708 10622
rect 8652 10610 8820 10612
rect 8652 10558 8654 10610
rect 8706 10558 8820 10610
rect 8652 10556 8820 10558
rect 8652 10546 8708 10556
rect 8764 9716 8820 10556
rect 9436 9940 9492 10668
rect 9548 10630 9604 10668
rect 9548 9940 9604 9950
rect 9436 9938 9604 9940
rect 9436 9886 9550 9938
rect 9602 9886 9604 9938
rect 9436 9884 9604 9886
rect 9548 9874 9604 9884
rect 8764 9660 9716 9716
rect 7532 9214 7534 9266
rect 7586 9214 7588 9266
rect 7532 9202 7588 9214
rect 7868 9492 7924 9502
rect 7868 9268 7924 9436
rect 7868 9266 8148 9268
rect 7868 9214 7870 9266
rect 7922 9214 8148 9266
rect 7868 9212 8148 9214
rect 7868 9202 7924 9212
rect 7420 8754 7476 8764
rect 8092 7474 8148 9212
rect 9660 9266 9716 9660
rect 9660 9214 9662 9266
rect 9714 9214 9716 9266
rect 9660 9202 9716 9214
rect 8428 9156 8484 9166
rect 8428 9062 8484 9100
rect 8988 9044 9044 9054
rect 8988 9042 9268 9044
rect 8988 8990 8990 9042
rect 9042 8990 9268 9042
rect 8988 8988 9268 8990
rect 8988 8978 9044 8988
rect 9212 8370 9268 8988
rect 9212 8318 9214 8370
rect 9266 8318 9268 8370
rect 8092 7422 8094 7474
rect 8146 7422 8148 7474
rect 8092 7410 8148 7422
rect 8652 7586 8708 7598
rect 8652 7534 8654 7586
rect 8706 7534 8708 7586
rect 7420 7364 7476 7374
rect 7420 7270 7476 7308
rect 8652 7364 8708 7534
rect 8876 7588 8932 7598
rect 8876 7474 8932 7532
rect 8876 7422 8878 7474
rect 8930 7422 8932 7474
rect 8876 7410 8932 7422
rect 8652 7298 8708 7308
rect 7756 7252 7812 7262
rect 7532 7250 7812 7252
rect 7532 7198 7758 7250
rect 7810 7198 7812 7250
rect 7532 7196 7812 7198
rect 7532 5122 7588 7196
rect 7756 7186 7812 7196
rect 9212 6916 9268 8318
rect 9660 7700 9716 7710
rect 9772 7700 9828 15092
rect 9884 11844 9940 16044
rect 10108 15988 10164 19068
rect 10108 15922 10164 15932
rect 9996 14756 10052 14766
rect 9996 13748 10052 14700
rect 10220 13860 10276 22876
rect 10556 21812 10612 24668
rect 11340 24610 11396 24622
rect 11340 24558 11342 24610
rect 11394 24558 11396 24610
rect 10872 24332 11136 24342
rect 10928 24276 10976 24332
rect 11032 24276 11080 24332
rect 10872 24266 11136 24276
rect 11340 23826 11396 24558
rect 11340 23774 11342 23826
rect 11394 23774 11396 23826
rect 11340 23762 11396 23774
rect 10872 22764 11136 22774
rect 10928 22708 10976 22764
rect 11032 22708 11080 22764
rect 10872 22698 11136 22708
rect 10556 21746 10612 21756
rect 11340 22148 11396 22158
rect 10444 21700 10500 21710
rect 10332 21588 10388 21598
rect 10332 21494 10388 21532
rect 10444 21028 10500 21644
rect 10332 20972 10500 21028
rect 10556 21586 10612 21598
rect 10556 21534 10558 21586
rect 10610 21534 10612 21586
rect 10556 21364 10612 21534
rect 10332 20580 10388 20972
rect 10444 20804 10500 20814
rect 10444 20710 10500 20748
rect 10556 20580 10612 21308
rect 10668 21586 10724 21598
rect 10668 21534 10670 21586
rect 10722 21534 10724 21586
rect 10668 20804 10724 21534
rect 11116 21588 11172 21598
rect 11116 21494 11172 21532
rect 11340 21474 11396 22092
rect 11564 21700 11620 26236
rect 11676 25730 11732 27806
rect 13804 27860 13860 27870
rect 12124 27746 12180 27758
rect 12124 27694 12126 27746
rect 12178 27694 12180 27746
rect 12124 27636 12180 27694
rect 11676 25678 11678 25730
rect 11730 25678 11732 25730
rect 11676 25666 11732 25678
rect 11788 26740 11844 26750
rect 11788 26514 11844 26684
rect 11788 26462 11790 26514
rect 11842 26462 11844 26514
rect 11676 24500 11732 24510
rect 11676 23938 11732 24444
rect 11676 23886 11678 23938
rect 11730 23886 11732 23938
rect 11676 23874 11732 23886
rect 11788 21812 11844 26462
rect 12012 25732 12068 25742
rect 12012 25638 12068 25676
rect 11788 21746 11844 21756
rect 11900 22146 11956 22158
rect 11900 22094 11902 22146
rect 11954 22094 11956 22146
rect 11564 21586 11620 21644
rect 11564 21534 11566 21586
rect 11618 21534 11620 21586
rect 11564 21522 11620 21534
rect 11340 21422 11342 21474
rect 11394 21422 11396 21474
rect 10872 21196 11136 21206
rect 10928 21140 10976 21196
rect 11032 21140 11080 21196
rect 10872 21130 11136 21140
rect 10780 20804 10836 20814
rect 10668 20802 10836 20804
rect 10668 20750 10782 20802
rect 10834 20750 10836 20802
rect 10668 20748 10836 20750
rect 10668 20580 10724 20590
rect 10332 20524 10500 20580
rect 10556 20578 10724 20580
rect 10556 20526 10670 20578
rect 10722 20526 10724 20578
rect 10556 20524 10724 20526
rect 10332 20244 10388 20254
rect 10332 19796 10388 20188
rect 10444 20130 10500 20524
rect 10668 20244 10724 20524
rect 10668 20178 10724 20188
rect 10780 20468 10836 20748
rect 10444 20078 10446 20130
rect 10498 20078 10500 20130
rect 10444 20066 10500 20078
rect 10780 20020 10836 20412
rect 11004 20804 11060 20814
rect 10668 19964 10836 20020
rect 10892 20020 10948 20030
rect 11004 20020 11060 20748
rect 11228 20802 11284 20814
rect 11228 20750 11230 20802
rect 11282 20750 11284 20802
rect 11228 20692 11284 20750
rect 11340 20804 11396 21422
rect 11452 21476 11508 21486
rect 11452 21382 11508 21420
rect 11900 21364 11956 22094
rect 11900 21298 11956 21308
rect 12012 21588 12068 21598
rect 11676 20916 11732 20926
rect 11676 20822 11732 20860
rect 11452 20804 11508 20814
rect 11340 20802 11508 20804
rect 11340 20750 11454 20802
rect 11506 20750 11508 20802
rect 11340 20748 11508 20750
rect 11228 20626 11284 20636
rect 10892 20018 11060 20020
rect 10892 19966 10894 20018
rect 10946 19966 11060 20018
rect 10892 19964 11060 19966
rect 10332 19740 10500 19796
rect 10332 16882 10388 16894
rect 10332 16830 10334 16882
rect 10386 16830 10388 16882
rect 10332 16212 10388 16830
rect 10444 16884 10500 19740
rect 10556 19794 10612 19806
rect 10556 19742 10558 19794
rect 10610 19742 10612 19794
rect 10556 19460 10612 19742
rect 10556 19394 10612 19404
rect 10556 16884 10612 16894
rect 10444 16882 10612 16884
rect 10444 16830 10558 16882
rect 10610 16830 10612 16882
rect 10444 16828 10612 16830
rect 10668 16884 10724 19964
rect 10892 19954 10948 19964
rect 11004 19796 11060 19806
rect 11004 19794 11284 19796
rect 11004 19742 11006 19794
rect 11058 19742 11284 19794
rect 11004 19740 11284 19742
rect 11004 19730 11060 19740
rect 10872 19628 11136 19638
rect 10928 19572 10976 19628
rect 11032 19572 11080 19628
rect 10872 19562 11136 19572
rect 10892 19124 10948 19134
rect 10892 19030 10948 19068
rect 11228 18900 11284 19740
rect 11340 19124 11396 19134
rect 11340 19030 11396 19068
rect 11228 18834 11284 18844
rect 10872 18060 11136 18070
rect 10928 18004 10976 18060
rect 11032 18004 11080 18060
rect 10872 17994 11136 18004
rect 10892 16884 10948 16894
rect 10668 16882 10948 16884
rect 10668 16830 10894 16882
rect 10946 16830 10948 16882
rect 10668 16828 10948 16830
rect 10556 16324 10612 16828
rect 10892 16660 10948 16828
rect 11116 16884 11172 16894
rect 11340 16884 11396 16894
rect 11452 16884 11508 20748
rect 11788 20692 11844 20702
rect 11676 20580 11732 20590
rect 11676 20486 11732 20524
rect 11676 20020 11732 20030
rect 11676 19926 11732 19964
rect 11788 19122 11844 20636
rect 11788 19070 11790 19122
rect 11842 19070 11844 19122
rect 11788 19058 11844 19070
rect 11900 20132 11956 20142
rect 11900 18450 11956 20076
rect 11900 18398 11902 18450
rect 11954 18398 11956 18450
rect 11900 18386 11956 18398
rect 11788 17780 11844 17790
rect 11676 17556 11732 17566
rect 11676 17462 11732 17500
rect 11676 17108 11732 17118
rect 11676 17014 11732 17052
rect 11116 16882 11284 16884
rect 11116 16830 11118 16882
rect 11170 16830 11284 16882
rect 11116 16828 11284 16830
rect 11116 16818 11172 16828
rect 10892 16594 10948 16604
rect 11228 16772 11284 16828
rect 11396 16828 11508 16884
rect 11564 16884 11620 16894
rect 11788 16884 11844 17724
rect 12012 17554 12068 21532
rect 12124 21140 12180 27580
rect 12908 27186 12964 27198
rect 12908 27134 12910 27186
rect 12962 27134 12964 27186
rect 12908 25732 12964 27134
rect 12908 25666 12964 25676
rect 12796 25508 12852 25518
rect 12796 25414 12852 25452
rect 13580 25508 13636 25518
rect 12572 25396 12628 25406
rect 12572 25302 12628 25340
rect 13580 25396 13636 25452
rect 13692 25396 13748 25406
rect 13580 25394 13748 25396
rect 13580 25342 13694 25394
rect 13746 25342 13748 25394
rect 13580 25340 13748 25342
rect 13468 24612 13524 24622
rect 13468 24518 13524 24556
rect 13580 23714 13636 25340
rect 13692 25330 13748 25340
rect 13580 23662 13582 23714
rect 13634 23662 13636 23714
rect 13580 22932 13636 23662
rect 13580 22866 13636 22876
rect 13804 22372 13860 27804
rect 14028 26908 14084 32956
rect 14252 32788 14308 32798
rect 14252 32694 14308 32732
rect 14364 32788 14420 32956
rect 14588 32788 14644 32798
rect 14364 32786 14588 32788
rect 14364 32734 14366 32786
rect 14418 32734 14588 32786
rect 14364 32732 14588 32734
rect 14364 32722 14420 32732
rect 14588 32722 14644 32732
rect 14140 32562 14196 32574
rect 14140 32510 14142 32562
rect 14194 32510 14196 32562
rect 14140 31780 14196 32510
rect 14588 32564 14644 32574
rect 14588 32470 14644 32508
rect 14140 31714 14196 31724
rect 14476 30994 14532 31006
rect 14476 30942 14478 30994
rect 14530 30942 14532 30994
rect 14476 30660 14532 30942
rect 14700 30772 14756 33292
rect 14812 33282 14868 33292
rect 15148 33348 15204 33358
rect 15148 33346 15316 33348
rect 15148 33294 15150 33346
rect 15202 33294 15316 33346
rect 15148 33292 15316 33294
rect 15148 33282 15204 33292
rect 14924 32900 14980 32910
rect 14924 32562 14980 32844
rect 15260 32676 15316 33292
rect 15708 33346 15764 33358
rect 15708 33294 15710 33346
rect 15762 33294 15764 33346
rect 15708 33124 15764 33294
rect 15708 33058 15764 33068
rect 15820 33122 15876 34412
rect 16044 34132 16100 34524
rect 16940 34354 16996 34860
rect 17052 34914 17108 35420
rect 17052 34862 17054 34914
rect 17106 34862 17108 34914
rect 17052 34850 17108 34862
rect 16940 34302 16942 34354
rect 16994 34302 16996 34354
rect 16940 34290 16996 34302
rect 17500 34692 17556 35644
rect 17612 35634 17668 35644
rect 17836 35588 17892 35756
rect 19292 35698 19348 35710
rect 19292 35646 19294 35698
rect 19346 35646 19348 35698
rect 18284 35588 18340 35598
rect 17836 35586 18340 35588
rect 17836 35534 18286 35586
rect 18338 35534 18340 35586
rect 17836 35532 18340 35534
rect 17724 35474 17780 35486
rect 17724 35422 17726 35474
rect 17778 35422 17780 35474
rect 17724 35026 17780 35422
rect 18284 35476 18340 35532
rect 19068 35588 19124 35598
rect 19292 35588 19348 35646
rect 19068 35586 19348 35588
rect 19068 35534 19070 35586
rect 19122 35534 19348 35586
rect 19068 35532 19348 35534
rect 20076 35586 20132 35598
rect 20076 35534 20078 35586
rect 20130 35534 20132 35586
rect 18284 35410 18340 35420
rect 18956 35476 19012 35486
rect 17724 34974 17726 35026
rect 17778 34974 17780 35026
rect 17724 34962 17780 34974
rect 18396 35026 18452 35038
rect 18396 34974 18398 35026
rect 18450 34974 18452 35026
rect 18060 34916 18116 34926
rect 18060 34822 18116 34860
rect 17500 34244 17556 34636
rect 17612 34244 17668 34254
rect 17500 34188 17612 34244
rect 17612 34178 17668 34188
rect 18284 34244 18340 34254
rect 15820 33070 15822 33122
rect 15874 33070 15876 33122
rect 15820 33058 15876 33070
rect 15932 34018 15988 34030
rect 15932 33966 15934 34018
rect 15986 33966 15988 34018
rect 15372 32676 15428 32686
rect 15932 32676 15988 33966
rect 15260 32674 15428 32676
rect 15260 32622 15374 32674
rect 15426 32622 15428 32674
rect 15260 32620 15428 32622
rect 14924 32510 14926 32562
rect 14978 32510 14980 32562
rect 14924 31948 14980 32510
rect 15148 32564 15204 32574
rect 15148 32470 15204 32508
rect 15372 32452 15428 32620
rect 15820 32620 15988 32676
rect 16044 33234 16100 34076
rect 17836 34132 17892 34142
rect 17836 34038 17892 34076
rect 18284 34130 18340 34188
rect 18284 34078 18286 34130
rect 18338 34078 18340 34130
rect 18284 34066 18340 34078
rect 18172 34020 18228 34030
rect 16044 33182 16046 33234
rect 16098 33182 16100 33234
rect 15372 32386 15428 32396
rect 15484 32564 15540 32574
rect 15820 32564 15876 32620
rect 15484 32562 15876 32564
rect 15484 32510 15486 32562
rect 15538 32510 15876 32562
rect 15484 32508 15876 32510
rect 14924 31892 15316 31948
rect 15260 31890 15316 31892
rect 15260 31838 15262 31890
rect 15314 31838 15316 31890
rect 15260 31826 15316 31838
rect 15036 31780 15092 31790
rect 15092 31724 15204 31780
rect 15036 31714 15092 31724
rect 14812 31556 14868 31566
rect 14812 30994 14868 31500
rect 14812 30942 14814 30994
rect 14866 30942 14868 30994
rect 14812 30930 14868 30942
rect 14924 30884 14980 30894
rect 14924 30790 14980 30828
rect 14700 30716 14868 30772
rect 14476 30594 14532 30604
rect 14364 30210 14420 30222
rect 14364 30158 14366 30210
rect 14418 30158 14420 30210
rect 14364 30100 14420 30158
rect 14700 30212 14756 30222
rect 14700 30118 14756 30156
rect 14364 30034 14420 30044
rect 14252 29426 14308 29438
rect 14252 29374 14254 29426
rect 14306 29374 14308 29426
rect 14252 28642 14308 29374
rect 14700 28756 14756 28766
rect 14700 28662 14756 28700
rect 14252 28590 14254 28642
rect 14306 28590 14308 28642
rect 14252 28084 14308 28590
rect 14252 28018 14308 28028
rect 14028 26852 14532 26908
rect 14252 24612 14308 24622
rect 13916 24500 13972 24510
rect 13916 24406 13972 24444
rect 14252 24500 14308 24556
rect 14252 24498 14420 24500
rect 14252 24446 14254 24498
rect 14306 24446 14420 24498
rect 14252 24444 14420 24446
rect 14252 24434 14308 24444
rect 13804 22316 13972 22372
rect 12236 22148 12292 22158
rect 12684 22148 12740 22158
rect 13468 22148 13524 22158
rect 12236 22146 12852 22148
rect 12236 22094 12238 22146
rect 12290 22094 12686 22146
rect 12738 22094 12852 22146
rect 12236 22092 12852 22094
rect 12236 22082 12292 22092
rect 12684 22082 12740 22092
rect 12684 21812 12740 21822
rect 12684 21718 12740 21756
rect 12124 21074 12180 21084
rect 12348 21474 12404 21486
rect 12348 21422 12350 21474
rect 12402 21422 12404 21474
rect 12236 20578 12292 20590
rect 12236 20526 12238 20578
rect 12290 20526 12292 20578
rect 12236 20468 12292 20526
rect 12348 20580 12404 21422
rect 12796 21252 12852 22092
rect 13468 22054 13524 22092
rect 13804 22148 13860 22158
rect 13804 22054 13860 22092
rect 13468 21812 13524 21822
rect 13468 21718 13524 21756
rect 13692 21586 13748 21598
rect 13692 21534 13694 21586
rect 13746 21534 13748 21586
rect 13244 21476 13300 21486
rect 13692 21476 13748 21534
rect 13244 21474 13748 21476
rect 13244 21422 13246 21474
rect 13298 21422 13748 21474
rect 13244 21420 13748 21422
rect 13244 21410 13300 21420
rect 13580 21252 13636 21262
rect 12796 21196 13412 21252
rect 12572 20580 12628 20590
rect 12348 20578 12628 20580
rect 12348 20526 12574 20578
rect 12626 20526 12628 20578
rect 12348 20524 12628 20526
rect 12236 20402 12292 20412
rect 12572 20244 12628 20524
rect 12572 20178 12628 20188
rect 13020 20018 13076 20030
rect 13020 19966 13022 20018
rect 13074 19966 13076 20018
rect 12124 19236 12180 19246
rect 12124 19142 12180 19180
rect 12684 19236 12740 19246
rect 12348 19122 12404 19134
rect 12348 19070 12350 19122
rect 12402 19070 12404 19122
rect 12348 18452 12404 19070
rect 12348 18386 12404 18396
rect 12684 19010 12740 19180
rect 12684 18958 12686 19010
rect 12738 18958 12740 19010
rect 12684 18004 12740 18958
rect 13020 18676 13076 19966
rect 13020 18610 13076 18620
rect 12012 17502 12014 17554
rect 12066 17502 12068 17554
rect 12012 17490 12068 17502
rect 12460 17948 12740 18004
rect 12908 18450 12964 18462
rect 12908 18398 12910 18450
rect 12962 18398 12964 18450
rect 12460 17666 12516 17948
rect 12908 17892 12964 18398
rect 13132 18452 13188 18462
rect 13132 18358 13188 18396
rect 12796 17836 12908 17892
rect 12572 17780 12628 17790
rect 12572 17686 12628 17724
rect 12460 17614 12462 17666
rect 12514 17614 12516 17666
rect 11900 16884 11956 16894
rect 11564 16882 11956 16884
rect 11564 16830 11566 16882
rect 11618 16830 11902 16882
rect 11954 16830 11956 16882
rect 11564 16828 11956 16830
rect 11340 16790 11396 16828
rect 11564 16818 11620 16828
rect 11732 16716 11844 16828
rect 11900 16818 11956 16828
rect 12348 16772 12404 16782
rect 11228 16548 11284 16716
rect 12348 16678 12404 16716
rect 10872 16492 11136 16502
rect 10928 16436 10976 16492
rect 11032 16436 11080 16492
rect 11228 16482 11284 16492
rect 12012 16658 12068 16670
rect 12012 16606 12014 16658
rect 12066 16606 12068 16658
rect 10872 16426 11136 16436
rect 11564 16436 11620 16446
rect 10556 16258 10612 16268
rect 10332 16118 10388 16156
rect 11116 16212 11172 16222
rect 11116 16098 11172 16156
rect 11116 16046 11118 16098
rect 11170 16046 11172 16098
rect 11116 16034 11172 16046
rect 11340 15988 11396 15998
rect 11340 15894 11396 15932
rect 11564 15986 11620 16380
rect 11564 15934 11566 15986
rect 11618 15934 11620 15986
rect 11564 15922 11620 15934
rect 11900 16324 11956 16334
rect 10444 15874 10500 15886
rect 10444 15822 10446 15874
rect 10498 15822 10500 15874
rect 10444 15316 10500 15822
rect 10444 15250 10500 15260
rect 11564 15316 11620 15326
rect 11564 15222 11620 15260
rect 10556 15092 10612 15102
rect 10556 13972 10612 15036
rect 10872 14924 11136 14934
rect 10928 14868 10976 14924
rect 11032 14868 11080 14924
rect 10872 14858 11136 14868
rect 10332 13860 10388 13870
rect 10220 13858 10500 13860
rect 10220 13806 10334 13858
rect 10386 13806 10500 13858
rect 10220 13804 10500 13806
rect 10332 13794 10388 13804
rect 9996 13746 10276 13748
rect 9996 13694 9998 13746
rect 10050 13694 10276 13746
rect 9996 13692 10276 13694
rect 9996 13682 10052 13692
rect 10220 13074 10276 13692
rect 10444 13636 10500 13804
rect 10556 13858 10612 13916
rect 10556 13806 10558 13858
rect 10610 13806 10612 13858
rect 10556 13794 10612 13806
rect 11452 13972 11508 13982
rect 11340 13636 11396 13646
rect 10444 13634 11396 13636
rect 10444 13582 11342 13634
rect 11394 13582 11396 13634
rect 10444 13580 11396 13582
rect 10220 13022 10222 13074
rect 10274 13022 10276 13074
rect 10220 13010 10276 13022
rect 9884 11788 10276 11844
rect 10108 10610 10164 10622
rect 10108 10558 10110 10610
rect 10162 10558 10164 10610
rect 10108 10500 10164 10558
rect 10108 10434 10164 10444
rect 10220 9380 10276 11788
rect 10444 11172 10500 11182
rect 10220 9314 10276 9324
rect 10332 9826 10388 9838
rect 10332 9774 10334 9826
rect 10386 9774 10388 9826
rect 9996 8820 10052 8830
rect 9996 8726 10052 8764
rect 9884 8260 9940 8270
rect 9884 8258 10052 8260
rect 9884 8206 9886 8258
rect 9938 8206 10052 8258
rect 9884 8204 10052 8206
rect 9884 8194 9940 8204
rect 9660 7698 9828 7700
rect 9660 7646 9662 7698
rect 9714 7646 9828 7698
rect 9660 7644 9828 7646
rect 9660 7588 9716 7644
rect 9660 7522 9716 7532
rect 9212 6850 9268 6860
rect 9772 6804 9828 7644
rect 9772 6738 9828 6748
rect 8988 6132 9044 6142
rect 8988 5906 9044 6076
rect 8988 5854 8990 5906
rect 9042 5854 9044 5906
rect 8988 5842 9044 5854
rect 9996 6132 10052 8204
rect 10332 6580 10388 9774
rect 10444 8260 10500 11116
rect 10556 10500 10612 10510
rect 10556 10406 10612 10444
rect 10668 9156 10724 13580
rect 11340 13570 11396 13580
rect 11452 13524 11508 13916
rect 11900 13970 11956 16268
rect 12012 15204 12068 16606
rect 12012 15138 12068 15148
rect 12124 16660 12180 16670
rect 11900 13918 11902 13970
rect 11954 13918 11956 13970
rect 11900 13906 11956 13918
rect 11452 13458 11508 13468
rect 11676 13746 11732 13758
rect 11676 13694 11678 13746
rect 11730 13694 11732 13746
rect 10872 13356 11136 13366
rect 10928 13300 10976 13356
rect 11032 13300 11080 13356
rect 10872 13290 11136 13300
rect 11676 12852 11732 13694
rect 12124 13746 12180 16604
rect 12460 16212 12516 17614
rect 12460 16146 12516 16156
rect 12684 17556 12740 17566
rect 12684 16996 12740 17500
rect 12684 16210 12740 16940
rect 12684 16158 12686 16210
rect 12738 16158 12740 16210
rect 12684 16146 12740 16158
rect 12236 15986 12292 15998
rect 12236 15934 12238 15986
rect 12290 15934 12292 15986
rect 12236 15316 12292 15934
rect 12236 15250 12292 15260
rect 12348 15988 12404 15998
rect 12348 14306 12404 15932
rect 12796 15314 12852 17836
rect 12908 17826 12964 17836
rect 12908 17442 12964 17454
rect 12908 17390 12910 17442
rect 12962 17390 12964 17442
rect 12908 16212 12964 17390
rect 12908 16146 12964 16156
rect 13020 16884 13076 16894
rect 12796 15262 12798 15314
rect 12850 15262 12852 15314
rect 12796 15148 12852 15262
rect 12348 14254 12350 14306
rect 12402 14254 12404 14306
rect 12348 14084 12404 14254
rect 12348 14018 12404 14028
rect 12460 15092 12852 15148
rect 12124 13694 12126 13746
rect 12178 13694 12180 13746
rect 12124 13682 12180 13694
rect 12348 13746 12404 13758
rect 12348 13694 12350 13746
rect 12402 13694 12404 13746
rect 11788 12852 11844 12862
rect 11676 12850 11844 12852
rect 11676 12798 11790 12850
rect 11842 12798 11844 12850
rect 11676 12796 11844 12798
rect 10872 11788 11136 11798
rect 10928 11732 10976 11788
rect 11032 11732 11080 11788
rect 10872 11722 11136 11732
rect 11788 11396 11844 12796
rect 12348 12852 12404 13694
rect 12348 12786 12404 12796
rect 11900 12738 11956 12750
rect 11900 12686 11902 12738
rect 11954 12686 11956 12738
rect 11900 12180 11956 12686
rect 12012 12180 12068 12190
rect 11900 12124 12012 12180
rect 12012 12114 12068 12124
rect 12348 12180 12404 12190
rect 12460 12180 12516 15092
rect 13020 14308 13076 16828
rect 13132 15316 13188 15326
rect 13132 15222 13188 15260
rect 13356 14868 13412 21196
rect 13580 20802 13636 21196
rect 13580 20750 13582 20802
rect 13634 20750 13636 20802
rect 13580 20738 13636 20750
rect 13468 20018 13524 20030
rect 13468 19966 13470 20018
rect 13522 19966 13524 20018
rect 13468 17780 13524 19966
rect 13468 17714 13524 17724
rect 13580 17892 13636 17902
rect 13580 17778 13636 17836
rect 13580 17726 13582 17778
rect 13634 17726 13636 17778
rect 13580 17714 13636 17726
rect 13580 16324 13636 16334
rect 13580 16210 13636 16268
rect 13580 16158 13582 16210
rect 13634 16158 13636 16210
rect 13580 16146 13636 16158
rect 13692 15148 13748 21420
rect 13916 19796 13972 22316
rect 14252 22148 14308 22158
rect 14252 22054 14308 22092
rect 13804 19348 13860 19358
rect 13916 19348 13972 19740
rect 13804 19346 13972 19348
rect 13804 19294 13806 19346
rect 13858 19294 13972 19346
rect 13804 19292 13972 19294
rect 14028 21924 14084 21934
rect 13804 19282 13860 19292
rect 13356 14802 13412 14812
rect 13580 15092 13748 15148
rect 13804 18004 13860 18014
rect 12684 14252 13076 14308
rect 12684 13746 12740 14252
rect 13020 13972 13076 13982
rect 13020 13878 13076 13916
rect 12684 13694 12686 13746
rect 12738 13694 12740 13746
rect 12684 13682 12740 13694
rect 13244 13860 13300 13870
rect 12908 13636 12964 13646
rect 12796 13634 12964 13636
rect 12796 13582 12910 13634
rect 12962 13582 12964 13634
rect 12796 13580 12964 13582
rect 12796 12850 12852 13580
rect 12908 13570 12964 13580
rect 12796 12798 12798 12850
rect 12850 12798 12852 12850
rect 12348 12178 12516 12180
rect 12348 12126 12350 12178
rect 12402 12126 12516 12178
rect 12348 12124 12516 12126
rect 12684 12180 12740 12190
rect 12124 12066 12180 12078
rect 12124 12014 12126 12066
rect 12178 12014 12180 12066
rect 12124 11396 12180 12014
rect 11788 11340 11956 11396
rect 11228 11170 11284 11182
rect 11228 11118 11230 11170
rect 11282 11118 11284 11170
rect 11228 10724 11284 11118
rect 11788 11172 11844 11182
rect 11788 10836 11844 11116
rect 11228 10658 11284 10668
rect 11676 10780 11844 10836
rect 11340 10500 11396 10510
rect 10872 10220 11136 10230
rect 10928 10164 10976 10220
rect 11032 10164 11080 10220
rect 10872 10154 11136 10164
rect 10668 9042 10724 9100
rect 10780 9492 10836 9502
rect 10780 9154 10836 9436
rect 10780 9102 10782 9154
rect 10834 9102 10836 9154
rect 10780 9090 10836 9102
rect 10668 8990 10670 9042
rect 10722 8990 10724 9042
rect 10668 8978 10724 8990
rect 11340 8932 11396 10444
rect 11676 10164 11732 10780
rect 11676 10098 11732 10108
rect 11788 10612 11844 10622
rect 11788 9828 11844 10556
rect 11788 9762 11844 9772
rect 11452 9156 11508 9166
rect 11452 9062 11508 9100
rect 11340 8876 11508 8932
rect 10872 8652 11136 8662
rect 10928 8596 10976 8652
rect 11032 8596 11080 8652
rect 10872 8586 11136 8596
rect 10444 8194 10500 8204
rect 10556 8148 10612 8158
rect 10556 8146 10836 8148
rect 10556 8094 10558 8146
rect 10610 8094 10836 8146
rect 10556 8092 10836 8094
rect 10556 8082 10612 8092
rect 10780 7698 10836 8092
rect 10780 7646 10782 7698
rect 10834 7646 10836 7698
rect 10780 7634 10836 7646
rect 11340 7700 11396 7710
rect 11116 7588 11172 7598
rect 11116 7494 11172 7532
rect 10872 7084 11136 7094
rect 10928 7028 10976 7084
rect 11032 7028 11080 7084
rect 10872 7018 11136 7028
rect 11340 6692 11396 7644
rect 11116 6690 11396 6692
rect 11116 6638 11342 6690
rect 11394 6638 11396 6690
rect 11116 6636 11396 6638
rect 11004 6580 11060 6590
rect 10332 6578 11060 6580
rect 10332 6526 11006 6578
rect 11058 6526 11060 6578
rect 10332 6524 11060 6526
rect 10108 6132 10164 6142
rect 10052 6130 10164 6132
rect 10052 6078 10110 6130
rect 10162 6078 10164 6130
rect 10052 6076 10164 6078
rect 8204 5796 8260 5806
rect 7532 5070 7534 5122
rect 7586 5070 7588 5122
rect 7532 5058 7588 5070
rect 7756 5794 8260 5796
rect 7756 5742 8206 5794
rect 8258 5742 8260 5794
rect 7756 5740 8260 5742
rect 7756 5010 7812 5740
rect 8204 5730 8260 5740
rect 8988 5684 9044 5694
rect 8988 5122 9044 5628
rect 9996 5124 10052 6076
rect 10108 6066 10164 6076
rect 10332 5906 10388 6524
rect 11004 6514 11060 6524
rect 11116 6356 11172 6636
rect 11340 6626 11396 6636
rect 10780 6300 11172 6356
rect 10780 6130 10836 6300
rect 10780 6078 10782 6130
rect 10834 6078 10836 6130
rect 10780 6066 10836 6078
rect 11116 6020 11172 6030
rect 11116 5926 11172 5964
rect 10332 5854 10334 5906
rect 10386 5854 10388 5906
rect 10332 5842 10388 5854
rect 10872 5516 11136 5526
rect 10928 5460 10976 5516
rect 11032 5460 11080 5516
rect 10872 5450 11136 5460
rect 8988 5070 8990 5122
rect 9042 5070 9044 5122
rect 8988 5058 9044 5070
rect 9660 5122 10052 5124
rect 9660 5070 9998 5122
rect 10050 5070 10052 5122
rect 9660 5068 10052 5070
rect 7756 4958 7758 5010
rect 7810 4958 7812 5010
rect 7756 4946 7812 4958
rect 9212 4900 9268 4910
rect 9212 4806 9268 4844
rect 9660 4338 9716 5068
rect 9996 5058 10052 5068
rect 10780 5012 10836 5022
rect 10780 4918 10836 4956
rect 10332 4900 10388 4910
rect 10332 4450 10388 4844
rect 10332 4398 10334 4450
rect 10386 4398 10388 4450
rect 10332 4386 10388 4398
rect 9660 4286 9662 4338
rect 9714 4286 9716 4338
rect 9660 4274 9716 4286
rect 10872 3948 11136 3958
rect 10928 3892 10976 3948
rect 11032 3892 11080 3948
rect 10872 3882 11136 3892
rect 6972 2370 7028 2380
rect 7644 3444 7700 3482
rect 7868 3444 7924 3454
rect 7644 3442 7924 3444
rect 7644 3390 7646 3442
rect 7698 3390 7870 3442
rect 7922 3390 7924 3442
rect 7644 3388 7924 3390
rect 7644 800 7700 3388
rect 7868 3378 7924 3388
rect 8204 3444 8260 3482
rect 11452 3388 11508 8876
rect 11788 8818 11844 8830
rect 11788 8766 11790 8818
rect 11842 8766 11844 8818
rect 11788 7588 11844 8766
rect 11788 7522 11844 7532
rect 11564 5684 11620 5694
rect 11564 5590 11620 5628
rect 11900 5682 11956 11340
rect 12124 11330 12180 11340
rect 12012 11282 12068 11294
rect 12012 11230 12014 11282
rect 12066 11230 12068 11282
rect 12012 10724 12068 11230
rect 12012 10658 12068 10668
rect 12124 11170 12180 11182
rect 12124 11118 12126 11170
rect 12178 11118 12180 11170
rect 12124 10388 12180 11118
rect 12348 10610 12404 12124
rect 12684 12086 12740 12124
rect 12684 11844 12740 11854
rect 12572 10612 12628 10622
rect 12348 10558 12350 10610
rect 12402 10558 12404 10610
rect 12348 10546 12404 10558
rect 12460 10610 12628 10612
rect 12460 10558 12574 10610
rect 12626 10558 12628 10610
rect 12460 10556 12628 10558
rect 12460 10388 12516 10556
rect 12572 10546 12628 10556
rect 12124 10332 12516 10388
rect 12012 10164 12068 10174
rect 12012 7364 12068 10108
rect 12460 9826 12516 9838
rect 12460 9774 12462 9826
rect 12514 9774 12516 9826
rect 12124 9604 12180 9614
rect 12460 9604 12516 9774
rect 12124 9602 12516 9604
rect 12124 9550 12126 9602
rect 12178 9550 12516 9602
rect 12124 9548 12516 9550
rect 12124 9538 12180 9548
rect 12348 9380 12404 9390
rect 12348 9154 12404 9324
rect 12348 9102 12350 9154
rect 12402 9102 12404 9154
rect 12348 9090 12404 9102
rect 12124 8818 12180 8830
rect 12124 8766 12126 8818
rect 12178 8766 12180 8818
rect 12124 7700 12180 8766
rect 12460 8596 12516 9548
rect 12460 8530 12516 8540
rect 12684 9154 12740 11788
rect 12796 11620 12852 12798
rect 13020 12852 13076 12862
rect 12908 12738 12964 12750
rect 12908 12686 12910 12738
rect 12962 12686 12964 12738
rect 12908 12068 12964 12686
rect 12908 12002 12964 12012
rect 13020 11844 13076 12796
rect 13020 11778 13076 11788
rect 12796 11564 13076 11620
rect 12796 11396 12852 11406
rect 12796 11282 12852 11340
rect 12796 11230 12798 11282
rect 12850 11230 12852 11282
rect 12796 10612 12852 11230
rect 12796 10546 12852 10556
rect 12908 11170 12964 11182
rect 12908 11118 12910 11170
rect 12962 11118 12964 11170
rect 12908 10500 12964 11118
rect 12908 10434 12964 10444
rect 12684 9102 12686 9154
rect 12738 9102 12740 9154
rect 12124 7634 12180 7644
rect 12572 8484 12628 8494
rect 12012 7298 12068 7308
rect 11900 5630 11902 5682
rect 11954 5630 11956 5682
rect 11900 4228 11956 5630
rect 12460 6018 12516 6030
rect 12460 5966 12462 6018
rect 12514 5966 12516 6018
rect 12460 4788 12516 5966
rect 12460 4722 12516 4732
rect 12460 4228 12516 4238
rect 11900 4226 12516 4228
rect 11900 4174 12462 4226
rect 12514 4174 12516 4226
rect 11900 4172 12516 4174
rect 12460 4162 12516 4172
rect 12572 4004 12628 8428
rect 12684 8370 12740 9102
rect 12796 9938 12852 9950
rect 12796 9886 12798 9938
rect 12850 9886 12852 9938
rect 12796 9156 12852 9886
rect 12796 9090 12852 9100
rect 12684 8318 12686 8370
rect 12738 8318 12740 8370
rect 12684 8306 12740 8318
rect 12684 5908 12740 5918
rect 12684 5814 12740 5852
rect 12908 5236 12964 5246
rect 13020 5236 13076 11564
rect 13244 9266 13300 13804
rect 13580 11060 13636 15092
rect 13692 14084 13748 14094
rect 13692 11844 13748 14028
rect 13804 12850 13860 17948
rect 14028 17444 14084 21868
rect 14140 21812 14196 21822
rect 14140 21718 14196 21756
rect 14364 21364 14420 24444
rect 14364 21298 14420 21308
rect 14476 21812 14532 26852
rect 14588 25508 14644 25518
rect 14588 24834 14644 25452
rect 14812 25172 14868 30716
rect 15036 30100 15092 30110
rect 14924 29426 14980 29438
rect 14924 29374 14926 29426
rect 14978 29374 14980 29426
rect 14924 28756 14980 29374
rect 14924 28690 14980 28700
rect 14924 28084 14980 28094
rect 14924 26290 14980 28028
rect 15036 28082 15092 30044
rect 15148 29538 15204 31724
rect 15484 31220 15540 32508
rect 15932 32452 15988 32462
rect 15932 32358 15988 32396
rect 16044 32228 16100 33182
rect 16268 33234 16324 33246
rect 16268 33182 16270 33234
rect 16322 33182 16324 33234
rect 16268 32788 16324 33182
rect 16716 33124 16772 33134
rect 16268 32722 16324 32732
rect 16380 33012 16436 33022
rect 16380 32786 16436 32956
rect 16380 32734 16382 32786
rect 16434 32734 16436 32786
rect 16380 32452 16436 32734
rect 16380 32386 16436 32396
rect 16716 32340 16772 33068
rect 16716 32274 16772 32284
rect 15372 31164 15540 31220
rect 15708 32172 16100 32228
rect 15260 30772 15316 30782
rect 15260 30098 15316 30716
rect 15260 30046 15262 30098
rect 15314 30046 15316 30098
rect 15260 30034 15316 30046
rect 15372 29876 15428 31164
rect 15148 29486 15150 29538
rect 15202 29486 15204 29538
rect 15148 29474 15204 29486
rect 15260 29820 15428 29876
rect 15484 30994 15540 31006
rect 15484 30942 15486 30994
rect 15538 30942 15540 30994
rect 15484 30100 15540 30942
rect 15596 30212 15652 30222
rect 15596 30118 15652 30156
rect 15036 28030 15038 28082
rect 15090 28030 15092 28082
rect 15036 28018 15092 28030
rect 14924 26238 14926 26290
rect 14978 26238 14980 26290
rect 14924 26226 14980 26238
rect 15260 25732 15316 29820
rect 15484 29652 15540 30044
rect 15484 29586 15540 29596
rect 15596 29428 15652 29438
rect 15484 29426 15652 29428
rect 15484 29374 15598 29426
rect 15650 29374 15652 29426
rect 15484 29372 15652 29374
rect 15708 29428 15764 32172
rect 18172 31948 18228 33964
rect 18396 33124 18452 34974
rect 18956 35026 19012 35420
rect 18956 34974 18958 35026
rect 19010 34974 19012 35026
rect 18956 34962 19012 34974
rect 19068 34244 19124 35532
rect 20076 34692 20132 35534
rect 20076 34636 20468 34692
rect 20412 34354 20468 34636
rect 20532 34524 20796 34534
rect 20588 34468 20636 34524
rect 20692 34468 20740 34524
rect 20532 34458 20796 34468
rect 20412 34302 20414 34354
rect 20466 34302 20468 34354
rect 20412 34290 20468 34302
rect 18844 34188 19124 34244
rect 18508 34018 18564 34030
rect 18508 33966 18510 34018
rect 18562 33966 18564 34018
rect 18508 33348 18564 33966
rect 18508 33282 18564 33292
rect 18732 34020 18788 34030
rect 18620 33236 18676 33246
rect 18620 33142 18676 33180
rect 18732 33234 18788 33964
rect 18732 33182 18734 33234
rect 18786 33182 18788 33234
rect 18732 33170 18788 33182
rect 18508 33124 18564 33134
rect 18396 33122 18564 33124
rect 18396 33070 18510 33122
rect 18562 33070 18564 33122
rect 18396 33068 18564 33070
rect 18844 33124 18900 34188
rect 20524 34132 20580 34142
rect 20524 34038 20580 34076
rect 19516 34020 19572 34030
rect 19516 33926 19572 33964
rect 20860 33684 20916 37324
rect 21308 36596 21364 39200
rect 21644 37492 21700 37502
rect 21308 36594 21588 36596
rect 21308 36542 21310 36594
rect 21362 36542 21588 36594
rect 21308 36540 21588 36542
rect 21308 36530 21364 36540
rect 21532 36482 21588 36540
rect 21532 36430 21534 36482
rect 21586 36430 21588 36482
rect 21532 36418 21588 36430
rect 21532 35140 21588 35150
rect 21532 34914 21588 35084
rect 21532 34862 21534 34914
rect 21586 34862 21588 34914
rect 21532 34850 21588 34862
rect 20636 33628 20916 33684
rect 21420 34132 21476 34142
rect 19740 33572 19796 33582
rect 19740 33460 19796 33516
rect 19292 33458 19796 33460
rect 19292 33406 19742 33458
rect 19794 33406 19796 33458
rect 19292 33404 19796 33406
rect 18956 33346 19012 33358
rect 18956 33294 18958 33346
rect 19010 33294 19012 33346
rect 18956 33236 19012 33294
rect 19292 33346 19348 33404
rect 19740 33394 19796 33404
rect 19292 33294 19294 33346
rect 19346 33294 19348 33346
rect 18956 33180 19236 33236
rect 18844 33068 19124 33124
rect 18172 31892 18452 31948
rect 18396 31890 18452 31892
rect 18396 31838 18398 31890
rect 18450 31838 18452 31890
rect 16156 31666 16212 31678
rect 16156 31614 16158 31666
rect 16210 31614 16212 31666
rect 15932 31554 15988 31566
rect 15932 31502 15934 31554
rect 15986 31502 15988 31554
rect 15932 31332 15988 31502
rect 16044 31556 16100 31566
rect 16044 31462 16100 31500
rect 15932 31276 16100 31332
rect 15820 30994 15876 31006
rect 15820 30942 15822 30994
rect 15874 30942 15876 30994
rect 15820 30436 15876 30942
rect 15820 30380 15988 30436
rect 15932 30098 15988 30380
rect 15932 30046 15934 30098
rect 15986 30046 15988 30098
rect 15820 29986 15876 29998
rect 15820 29934 15822 29986
rect 15874 29934 15876 29986
rect 15820 29540 15876 29934
rect 15932 29988 15988 30046
rect 16044 30100 16100 31276
rect 16156 30324 16212 31614
rect 17836 31668 17892 31678
rect 17836 31220 17892 31612
rect 18396 31332 18452 31838
rect 18508 31892 18564 33068
rect 18956 32564 19012 32574
rect 18508 31826 18564 31836
rect 18844 32562 19012 32564
rect 18844 32510 18958 32562
rect 19010 32510 19012 32562
rect 18844 32508 19012 32510
rect 18844 31778 18900 32508
rect 18956 32498 19012 32508
rect 18844 31726 18846 31778
rect 18898 31726 18900 31778
rect 18844 31668 18900 31726
rect 18396 31266 18452 31276
rect 18508 31612 18900 31668
rect 18956 31892 19012 31902
rect 17948 31220 18004 31230
rect 17836 31218 18004 31220
rect 17836 31166 17950 31218
rect 18002 31166 18004 31218
rect 17836 31164 18004 31166
rect 17948 31154 18004 31164
rect 18508 31218 18564 31612
rect 18508 31166 18510 31218
rect 18562 31166 18564 31218
rect 18508 31154 18564 31166
rect 16380 31106 16436 31118
rect 16380 31054 16382 31106
rect 16434 31054 16436 31106
rect 16380 30996 16436 31054
rect 17948 30996 18004 31006
rect 18396 30996 18452 31006
rect 18620 30996 18676 31006
rect 16380 30940 16660 30996
rect 16268 30884 16324 30894
rect 16268 30882 16548 30884
rect 16268 30830 16270 30882
rect 16322 30830 16548 30882
rect 16268 30828 16548 30830
rect 16268 30818 16324 30828
rect 16492 30436 16548 30828
rect 16492 30342 16548 30380
rect 16156 30258 16212 30268
rect 16604 30212 16660 30940
rect 16492 30156 16660 30212
rect 16828 30882 16884 30894
rect 16828 30830 16830 30882
rect 16882 30830 16884 30882
rect 16380 30100 16436 30110
rect 16044 30044 16380 30100
rect 16380 30006 16436 30044
rect 15932 29922 15988 29932
rect 16268 29652 16324 29662
rect 16268 29558 16324 29596
rect 15820 29484 15988 29540
rect 15932 29428 15988 29484
rect 16492 29428 16548 30156
rect 15708 29372 15876 29428
rect 15932 29426 16548 29428
rect 15932 29374 16494 29426
rect 16546 29374 16548 29426
rect 15932 29372 16548 29374
rect 14924 25676 15316 25732
rect 15372 29314 15428 29326
rect 15372 29262 15374 29314
rect 15426 29262 15428 29314
rect 15372 27858 15428 29262
rect 15484 28420 15540 29372
rect 15596 29362 15652 29372
rect 15708 29204 15764 29214
rect 15708 28530 15764 29148
rect 15708 28478 15710 28530
rect 15762 28478 15764 28530
rect 15708 28466 15764 28478
rect 15596 28420 15652 28430
rect 15484 28364 15596 28420
rect 15596 28354 15652 28364
rect 15372 27806 15374 27858
rect 15426 27806 15428 27858
rect 14924 25506 14980 25676
rect 14924 25454 14926 25506
rect 14978 25454 14980 25506
rect 14924 25442 14980 25454
rect 14812 25106 14868 25116
rect 14588 24782 14590 24834
rect 14642 24782 14644 24834
rect 14588 24770 14644 24782
rect 14812 24948 14868 24958
rect 14812 24834 14868 24892
rect 14812 24782 14814 24834
rect 14866 24782 14868 24834
rect 14812 24276 14868 24782
rect 14812 24210 14868 24220
rect 15372 24164 15428 27806
rect 15596 27748 15652 27758
rect 15596 27654 15652 27692
rect 15820 26908 15876 29372
rect 16156 29092 16212 29102
rect 16156 28642 16212 29036
rect 16156 28590 16158 28642
rect 16210 28590 16212 28642
rect 16156 28578 16212 28590
rect 16268 27748 16324 27758
rect 16268 27654 16324 27692
rect 15820 26852 16324 26908
rect 16044 26178 16100 26190
rect 16044 26126 16046 26178
rect 16098 26126 16100 26178
rect 15484 25620 15540 25630
rect 15484 25526 15540 25564
rect 15820 25620 15876 25630
rect 15876 25564 15988 25620
rect 15820 25554 15876 25564
rect 15708 25508 15764 25518
rect 15484 25172 15540 25182
rect 15484 24834 15540 25116
rect 15708 24836 15764 25452
rect 15484 24782 15486 24834
rect 15538 24782 15540 24834
rect 15484 24770 15540 24782
rect 15596 24780 15764 24836
rect 15820 24948 15876 24958
rect 15148 24108 15428 24164
rect 15484 24612 15540 24622
rect 15484 24276 15540 24556
rect 15036 23044 15092 23054
rect 15036 22950 15092 22988
rect 14476 21252 14532 21756
rect 14476 21186 14532 21196
rect 14924 22036 14980 22046
rect 14252 20692 14308 20702
rect 14252 20690 14756 20692
rect 14252 20638 14254 20690
rect 14306 20638 14756 20690
rect 14252 20636 14756 20638
rect 14252 20626 14308 20636
rect 14476 20018 14532 20030
rect 14476 19966 14478 20018
rect 14530 19966 14532 20018
rect 14364 19012 14420 19022
rect 14364 18918 14420 18956
rect 14252 18676 14308 18686
rect 14252 17780 14308 18620
rect 14476 18452 14532 19966
rect 14700 19346 14756 20636
rect 14812 19906 14868 19918
rect 14812 19854 14814 19906
rect 14866 19854 14868 19906
rect 14812 19460 14868 19854
rect 14812 19394 14868 19404
rect 14700 19294 14702 19346
rect 14754 19294 14756 19346
rect 14700 19282 14756 19294
rect 14812 19124 14868 19134
rect 14812 19030 14868 19068
rect 14588 19010 14644 19022
rect 14588 18958 14590 19010
rect 14642 18958 14644 19010
rect 14588 18788 14644 18958
rect 14588 18732 14868 18788
rect 14700 18564 14756 18574
rect 14588 18452 14644 18462
rect 14476 18450 14644 18452
rect 14476 18398 14590 18450
rect 14642 18398 14644 18450
rect 14476 18396 14644 18398
rect 14588 18340 14644 18396
rect 14588 18274 14644 18284
rect 14700 18338 14756 18508
rect 14700 18286 14702 18338
rect 14754 18286 14756 18338
rect 14700 18274 14756 18286
rect 14252 17666 14308 17724
rect 14700 17780 14756 17790
rect 14700 17686 14756 17724
rect 14252 17614 14254 17666
rect 14306 17614 14308 17666
rect 14252 17602 14308 17614
rect 14028 17388 14196 17444
rect 14028 17220 14084 17230
rect 13916 15316 13972 15326
rect 13916 14642 13972 15260
rect 13916 14590 13918 14642
rect 13970 14590 13972 14642
rect 13916 14578 13972 14590
rect 13916 13860 13972 13870
rect 13916 13766 13972 13804
rect 14028 13858 14084 17164
rect 14140 15148 14196 17388
rect 14476 16770 14532 16782
rect 14476 16718 14478 16770
rect 14530 16718 14532 16770
rect 14476 16212 14532 16718
rect 14588 16212 14644 16222
rect 14476 16210 14644 16212
rect 14476 16158 14590 16210
rect 14642 16158 14644 16210
rect 14476 16156 14644 16158
rect 14588 16146 14644 16156
rect 14364 16100 14420 16110
rect 14364 15988 14420 16044
rect 14476 15988 14532 15998
rect 14364 15986 14532 15988
rect 14364 15934 14478 15986
rect 14530 15934 14532 15986
rect 14364 15932 14532 15934
rect 14476 15922 14532 15932
rect 14252 15876 14308 15886
rect 14700 15876 14756 15886
rect 14812 15876 14868 18732
rect 14924 17220 14980 21980
rect 15148 21810 15204 24108
rect 15260 23940 15316 23950
rect 15484 23940 15540 24220
rect 15260 23938 15540 23940
rect 15260 23886 15262 23938
rect 15314 23886 15540 23938
rect 15260 23884 15540 23886
rect 15260 23874 15316 23884
rect 15372 23604 15428 23614
rect 15372 23492 15428 23548
rect 15148 21758 15150 21810
rect 15202 21758 15204 21810
rect 15148 21746 15204 21758
rect 15260 23436 15428 23492
rect 15260 21588 15316 23436
rect 15596 23380 15652 24780
rect 15820 24722 15876 24892
rect 15820 24670 15822 24722
rect 15874 24670 15876 24722
rect 15820 23604 15876 24670
rect 15820 23538 15876 23548
rect 15708 23380 15764 23390
rect 15932 23380 15988 25564
rect 16044 25508 16100 26126
rect 16044 25506 16212 25508
rect 16044 25454 16046 25506
rect 16098 25454 16212 25506
rect 16044 25452 16212 25454
rect 16044 25442 16100 25452
rect 16156 24610 16212 25452
rect 16156 24558 16158 24610
rect 16210 24558 16212 24610
rect 16156 23940 16212 24558
rect 16268 24050 16324 26852
rect 16268 23998 16270 24050
rect 16322 23998 16324 24050
rect 16268 23986 16324 23998
rect 16156 23874 16212 23884
rect 15596 23378 15764 23380
rect 15596 23326 15710 23378
rect 15762 23326 15764 23378
rect 15596 23324 15764 23326
rect 15708 23314 15764 23324
rect 15820 23324 15988 23380
rect 16268 23380 16324 23390
rect 15484 23266 15540 23278
rect 15484 23214 15486 23266
rect 15538 23214 15540 23266
rect 15372 23156 15428 23166
rect 15372 23062 15428 23100
rect 15484 23044 15540 23214
rect 15484 21924 15540 22988
rect 15484 21858 15540 21868
rect 15596 21700 15652 21710
rect 15596 21606 15652 21644
rect 15148 21532 15316 21588
rect 15708 21586 15764 21598
rect 15708 21534 15710 21586
rect 15762 21534 15764 21586
rect 15036 19794 15092 19806
rect 15036 19742 15038 19794
rect 15090 19742 15092 19794
rect 15036 19460 15092 19742
rect 15036 19394 15092 19404
rect 15148 19012 15204 21532
rect 15708 20580 15764 21534
rect 15708 20514 15764 20524
rect 15820 20356 15876 23324
rect 16268 23286 16324 23324
rect 16044 23268 16100 23278
rect 16044 23174 16100 23212
rect 15932 23156 15988 23166
rect 15932 22372 15988 23100
rect 15932 22306 15988 22316
rect 16268 22260 16324 22270
rect 16268 22166 16324 22204
rect 15932 21588 15988 21598
rect 15932 21494 15988 21532
rect 16380 21252 16436 29372
rect 16492 29362 16548 29372
rect 16716 29988 16772 29998
rect 16716 29428 16772 29932
rect 16716 29334 16772 29372
rect 16604 29316 16660 29326
rect 16604 29222 16660 29260
rect 16828 28980 16884 30830
rect 16828 28914 16884 28924
rect 17052 30884 17108 30894
rect 17052 28642 17108 30828
rect 17724 30772 17780 30782
rect 17612 30770 17780 30772
rect 17612 30718 17726 30770
rect 17778 30718 17780 30770
rect 17612 30716 17780 30718
rect 17388 30436 17444 30446
rect 17276 30212 17332 30222
rect 17276 30118 17332 30156
rect 17388 29650 17444 30380
rect 17612 30100 17668 30716
rect 17724 30706 17780 30716
rect 17948 30434 18004 30940
rect 18060 30994 18452 30996
rect 18060 30942 18398 30994
rect 18450 30942 18452 30994
rect 18060 30940 18452 30942
rect 18060 30882 18116 30940
rect 18396 30930 18452 30940
rect 18508 30994 18676 30996
rect 18508 30942 18622 30994
rect 18674 30942 18676 30994
rect 18508 30940 18676 30942
rect 18060 30830 18062 30882
rect 18114 30830 18116 30882
rect 18060 30818 18116 30830
rect 17948 30382 17950 30434
rect 18002 30382 18004 30434
rect 17948 30370 18004 30382
rect 17388 29598 17390 29650
rect 17442 29598 17444 29650
rect 17388 29586 17444 29598
rect 17500 29652 17556 29662
rect 17500 29558 17556 29596
rect 17612 29426 17668 30044
rect 17612 29374 17614 29426
rect 17666 29374 17668 29426
rect 17052 28590 17054 28642
rect 17106 28590 17108 28642
rect 17052 28578 17108 28590
rect 17500 29092 17556 29102
rect 17164 28420 17220 28430
rect 17164 28326 17220 28364
rect 16828 27860 16884 27870
rect 16828 27746 16884 27804
rect 16828 27694 16830 27746
rect 16882 27694 16884 27746
rect 16828 27682 16884 27694
rect 16492 27636 16548 27646
rect 16492 27542 16548 27580
rect 17388 27074 17444 27086
rect 17388 27022 17390 27074
rect 17442 27022 17444 27074
rect 16492 26964 16548 27002
rect 16828 26964 16884 27002
rect 16492 26962 16828 26964
rect 16492 26910 16494 26962
rect 16546 26910 16828 26962
rect 16492 26908 16828 26910
rect 16492 26402 16548 26908
rect 16828 26898 16884 26908
rect 17164 26962 17220 26974
rect 17164 26910 17166 26962
rect 17218 26910 17220 26962
rect 16492 26350 16494 26402
rect 16546 26350 16548 26402
rect 16492 26338 16548 26350
rect 16828 26292 16884 26302
rect 17164 26292 17220 26910
rect 17388 26964 17444 27022
rect 17388 26898 17444 26908
rect 16828 26290 17220 26292
rect 16828 26238 16830 26290
rect 16882 26238 17220 26290
rect 16828 26236 17220 26238
rect 16604 26178 16660 26190
rect 16604 26126 16606 26178
rect 16658 26126 16660 26178
rect 16380 21186 16436 21196
rect 16492 25732 16548 25742
rect 16492 22260 16548 25676
rect 16604 24612 16660 26126
rect 16716 25508 16772 25518
rect 16716 25414 16772 25452
rect 16716 24948 16772 24958
rect 16828 24948 16884 26236
rect 16772 24892 16884 24948
rect 16716 24882 16772 24892
rect 17500 24834 17556 29036
rect 17612 28084 17668 29374
rect 17836 30210 17892 30222
rect 17836 30158 17838 30210
rect 17890 30158 17892 30210
rect 17836 29538 17892 30158
rect 17836 29486 17838 29538
rect 17890 29486 17892 29538
rect 17836 29316 17892 29486
rect 17836 29250 17892 29260
rect 18284 29316 18340 29326
rect 18284 28642 18340 29260
rect 18284 28590 18286 28642
rect 18338 28590 18340 28642
rect 18284 28578 18340 28590
rect 18396 28420 18452 28430
rect 17724 28084 17780 28094
rect 17612 28082 17780 28084
rect 17612 28030 17726 28082
rect 17778 28030 17780 28082
rect 17612 28028 17780 28030
rect 17724 28018 17780 28028
rect 17836 27860 17892 27870
rect 17836 27766 17892 27804
rect 18172 27858 18228 27870
rect 18172 27806 18174 27858
rect 18226 27806 18228 27858
rect 17500 24782 17502 24834
rect 17554 24782 17556 24834
rect 16604 24546 16660 24556
rect 16716 24722 16772 24734
rect 16716 24670 16718 24722
rect 16770 24670 16772 24722
rect 16716 24500 16772 24670
rect 16716 24434 16772 24444
rect 17500 24388 17556 24782
rect 17500 24322 17556 24332
rect 17612 27636 17668 27646
rect 16716 23940 16772 23950
rect 16716 23846 16772 23884
rect 17500 23938 17556 23950
rect 17500 23886 17502 23938
rect 17554 23886 17556 23938
rect 17500 23380 17556 23886
rect 17500 23314 17556 23324
rect 16604 23044 16660 23054
rect 16604 22950 16660 22988
rect 17276 22372 17332 22382
rect 17276 22370 17444 22372
rect 17276 22318 17278 22370
rect 17330 22318 17444 22370
rect 17276 22316 17444 22318
rect 17276 22306 17332 22316
rect 16604 22260 16660 22270
rect 16492 22258 16660 22260
rect 16492 22206 16606 22258
rect 16658 22206 16660 22258
rect 16492 22204 16660 22206
rect 16380 20914 16436 20926
rect 16380 20862 16382 20914
rect 16434 20862 16436 20914
rect 16380 20692 16436 20862
rect 16380 20626 16436 20636
rect 15820 20300 16324 20356
rect 16268 20130 16324 20300
rect 16268 20078 16270 20130
rect 16322 20078 16324 20130
rect 16268 20066 16324 20078
rect 16044 20020 16100 20030
rect 15260 20018 16100 20020
rect 15260 19966 16046 20018
rect 16098 19966 16100 20018
rect 15260 19964 16100 19966
rect 15260 19234 15316 19964
rect 16044 19954 16100 19964
rect 16380 20020 16436 20030
rect 16380 19926 16436 19964
rect 16268 19908 16324 19918
rect 16156 19796 16212 19806
rect 15820 19684 15876 19694
rect 15260 19182 15262 19234
rect 15314 19182 15316 19234
rect 15260 19170 15316 19182
rect 15708 19234 15764 19246
rect 15708 19182 15710 19234
rect 15762 19182 15764 19234
rect 15148 18956 15540 19012
rect 15372 18340 15428 18350
rect 15036 18228 15092 18238
rect 15036 18134 15092 18172
rect 15372 17780 15428 18284
rect 14924 17154 14980 17164
rect 15148 17778 15428 17780
rect 15148 17726 15374 17778
rect 15426 17726 15428 17778
rect 15148 17724 15428 17726
rect 15148 16100 15204 17724
rect 15372 17714 15428 17724
rect 15260 16884 15316 16894
rect 15260 16882 15428 16884
rect 15260 16830 15262 16882
rect 15314 16830 15428 16882
rect 15260 16828 15428 16830
rect 15260 16818 15316 16828
rect 15036 16044 15204 16100
rect 14252 15874 14420 15876
rect 14252 15822 14254 15874
rect 14306 15822 14420 15874
rect 14252 15820 14420 15822
rect 14252 15810 14308 15820
rect 14364 15652 14420 15820
rect 14756 15820 14868 15876
rect 14924 15874 14980 15886
rect 14924 15822 14926 15874
rect 14978 15822 14980 15874
rect 14700 15782 14756 15820
rect 14924 15652 14980 15822
rect 14364 15596 14980 15652
rect 15036 15540 15092 16044
rect 15260 15986 15316 15998
rect 15260 15934 15262 15986
rect 15314 15934 15316 15986
rect 14924 15484 15092 15540
rect 15148 15874 15204 15886
rect 15148 15822 15150 15874
rect 15202 15822 15204 15874
rect 14588 15316 14644 15326
rect 14588 15222 14644 15260
rect 14700 15204 14756 15242
rect 14140 15092 14420 15148
rect 14700 15138 14756 15148
rect 14028 13806 14030 13858
rect 14082 13806 14084 13858
rect 14028 13794 14084 13806
rect 13916 13524 13972 13534
rect 13916 13430 13972 13468
rect 13804 12798 13806 12850
rect 13858 12798 13860 12850
rect 13804 12786 13860 12798
rect 14028 12852 14084 12862
rect 14028 12758 14084 12796
rect 14252 12738 14308 12750
rect 14252 12686 14254 12738
rect 14306 12686 14308 12738
rect 14252 12178 14308 12686
rect 14252 12126 14254 12178
rect 14306 12126 14308 12178
rect 14252 12114 14308 12126
rect 13804 11844 13860 11854
rect 13692 11788 13804 11844
rect 13804 11282 13860 11788
rect 13804 11230 13806 11282
rect 13858 11230 13860 11282
rect 13804 11218 13860 11230
rect 14028 11282 14084 11294
rect 14028 11230 14030 11282
rect 14082 11230 14084 11282
rect 14028 11172 14084 11230
rect 14028 11106 14084 11116
rect 14252 11170 14308 11182
rect 14252 11118 14254 11170
rect 14306 11118 14308 11170
rect 13580 11004 13860 11060
rect 13580 9828 13636 9838
rect 13580 9734 13636 9772
rect 13244 9214 13246 9266
rect 13298 9214 13300 9266
rect 13244 9202 13300 9214
rect 13468 9154 13524 9166
rect 13468 9102 13470 9154
rect 13522 9102 13524 9154
rect 13468 8484 13524 9102
rect 13580 9156 13636 9166
rect 13580 9062 13636 9100
rect 13468 8418 13524 8428
rect 13580 8034 13636 8046
rect 13580 7982 13582 8034
rect 13634 7982 13636 8034
rect 13580 7700 13636 7982
rect 13132 6916 13188 6926
rect 13132 6132 13188 6860
rect 13580 6692 13636 7644
rect 13804 7476 13860 11004
rect 14252 10610 14308 11118
rect 14252 10558 14254 10610
rect 14306 10558 14308 10610
rect 14252 10546 14308 10558
rect 14252 9940 14308 9950
rect 14252 9846 14308 9884
rect 13916 9380 13972 9390
rect 13916 8372 13972 9324
rect 14028 9156 14084 9166
rect 14028 9062 14084 9100
rect 14028 8372 14084 8382
rect 13916 8370 14084 8372
rect 13916 8318 14030 8370
rect 14082 8318 14084 8370
rect 13916 8316 14084 8318
rect 13804 7410 13860 7420
rect 14028 7140 14084 8316
rect 14028 7074 14084 7084
rect 14252 7700 14308 7710
rect 14252 6802 14308 7644
rect 14252 6750 14254 6802
rect 14306 6750 14308 6802
rect 14252 6738 14308 6750
rect 14364 6804 14420 15092
rect 14700 14532 14756 14542
rect 14924 14532 14980 15484
rect 15036 15204 15092 15214
rect 15036 15090 15092 15148
rect 15036 15038 15038 15090
rect 15090 15038 15092 15090
rect 15036 15026 15092 15038
rect 15148 14532 15204 15822
rect 15260 15428 15316 15934
rect 15260 15362 15316 15372
rect 14700 14530 14980 14532
rect 14700 14478 14702 14530
rect 14754 14478 14980 14530
rect 14700 14476 14980 14478
rect 14700 14466 14756 14476
rect 14924 14420 14980 14476
rect 14924 14354 14980 14364
rect 15036 14476 15204 14532
rect 15036 14196 15092 14476
rect 15260 14420 15316 14430
rect 15148 14308 15204 14318
rect 15260 14308 15316 14364
rect 15148 14306 15316 14308
rect 15148 14254 15150 14306
rect 15202 14254 15316 14306
rect 15148 14252 15316 14254
rect 15148 14242 15204 14252
rect 14924 14140 15092 14196
rect 14924 13524 14980 14140
rect 14924 13458 14980 13468
rect 15036 13412 15092 13422
rect 14588 12962 14644 12974
rect 14588 12910 14590 12962
rect 14642 12910 14644 12962
rect 14588 12740 14644 12910
rect 15036 12740 15092 13356
rect 15372 13300 15428 16828
rect 15484 15876 15540 18956
rect 15708 17668 15764 19182
rect 15708 17574 15764 17612
rect 15708 17332 15764 17342
rect 15708 16996 15764 17276
rect 15708 16930 15764 16940
rect 15596 16882 15652 16894
rect 15596 16830 15598 16882
rect 15650 16830 15652 16882
rect 15596 16100 15652 16830
rect 15596 16034 15652 16044
rect 15708 16772 15764 16782
rect 15708 16098 15764 16716
rect 15708 16046 15710 16098
rect 15762 16046 15764 16098
rect 15708 16034 15764 16046
rect 15820 16212 15876 19628
rect 16044 19012 16100 19022
rect 16044 18918 16100 18956
rect 15932 18788 15988 18798
rect 15932 17556 15988 18732
rect 16156 18676 16212 19740
rect 16268 19122 16324 19852
rect 16492 19460 16548 22204
rect 16604 22194 16660 22204
rect 17052 22260 17108 22270
rect 16828 22146 16884 22158
rect 16828 22094 16830 22146
rect 16882 22094 16884 22146
rect 16828 21924 16884 22094
rect 16828 21858 16884 21868
rect 16940 22146 16996 22158
rect 16940 22094 16942 22146
rect 16994 22094 16996 22146
rect 16604 21812 16660 21822
rect 16604 21718 16660 21756
rect 16940 21700 16996 22094
rect 16940 21634 16996 21644
rect 17052 22146 17108 22204
rect 17052 22094 17054 22146
rect 17106 22094 17108 22146
rect 16716 21252 16772 21262
rect 16772 21196 16884 21252
rect 16716 21186 16772 21196
rect 16716 20692 16772 20702
rect 16604 20356 16660 20366
rect 16604 19684 16660 20300
rect 16716 20130 16772 20636
rect 16828 20580 16884 21196
rect 16940 20916 16996 20926
rect 16940 20802 16996 20860
rect 16940 20750 16942 20802
rect 16994 20750 16996 20802
rect 16940 20738 16996 20750
rect 16828 20524 16996 20580
rect 16716 20078 16718 20130
rect 16770 20078 16772 20130
rect 16716 20066 16772 20078
rect 16604 19618 16660 19628
rect 16828 19794 16884 19806
rect 16828 19742 16830 19794
rect 16882 19742 16884 19794
rect 16492 19404 16660 19460
rect 16268 19070 16270 19122
rect 16322 19070 16324 19122
rect 16268 19058 16324 19070
rect 16492 19234 16548 19246
rect 16492 19182 16494 19234
rect 16546 19182 16548 19234
rect 16380 19010 16436 19022
rect 16380 18958 16382 19010
rect 16434 18958 16436 19010
rect 16380 18900 16436 18958
rect 16380 18834 16436 18844
rect 16156 18620 16436 18676
rect 16156 18340 16212 18350
rect 16156 18246 16212 18284
rect 16156 17892 16212 17902
rect 16156 17556 16212 17836
rect 15932 17462 15988 17500
rect 16044 17554 16212 17556
rect 16044 17502 16158 17554
rect 16210 17502 16212 17554
rect 16044 17500 16212 17502
rect 15820 16100 15876 16156
rect 15932 16100 15988 16110
rect 15820 16098 15988 16100
rect 15820 16046 15934 16098
rect 15986 16046 15988 16098
rect 15820 16044 15988 16046
rect 15932 16034 15988 16044
rect 16044 15988 16100 17500
rect 16156 17490 16212 17500
rect 16268 17444 16324 17454
rect 16268 17350 16324 17388
rect 16380 17332 16436 18620
rect 16492 18116 16548 19182
rect 16492 18050 16548 18060
rect 16492 17556 16548 17566
rect 16604 17556 16660 19404
rect 16828 19124 16884 19742
rect 16940 19234 16996 20524
rect 16940 19182 16942 19234
rect 16994 19182 16996 19234
rect 16940 19170 16996 19182
rect 16716 18676 16772 18686
rect 16716 17778 16772 18620
rect 16828 18564 16884 19068
rect 17052 19012 17108 22094
rect 17388 21700 17444 22316
rect 17276 21588 17332 21598
rect 17276 20914 17332 21532
rect 17276 20862 17278 20914
rect 17330 20862 17332 20914
rect 17276 20850 17332 20862
rect 17276 20692 17332 20702
rect 17164 20580 17220 20590
rect 17164 19908 17220 20524
rect 17164 19842 17220 19852
rect 17276 20578 17332 20636
rect 17276 20526 17278 20578
rect 17330 20526 17332 20578
rect 17276 19796 17332 20526
rect 17276 19730 17332 19740
rect 17388 19794 17444 21644
rect 17500 19908 17556 19918
rect 17500 19814 17556 19852
rect 17388 19742 17390 19794
rect 17442 19742 17444 19794
rect 17388 19730 17444 19742
rect 17612 19572 17668 27580
rect 18172 27412 18228 27806
rect 18172 27346 18228 27356
rect 18284 27636 18340 27646
rect 18284 27298 18340 27580
rect 18284 27246 18286 27298
rect 18338 27246 18340 27298
rect 18284 27234 18340 27246
rect 18396 26908 18452 28364
rect 18508 27186 18564 30940
rect 18620 30930 18676 30940
rect 18620 30210 18676 30222
rect 18620 30158 18622 30210
rect 18674 30158 18676 30210
rect 18620 29652 18676 30158
rect 18620 29586 18676 29596
rect 18732 27972 18788 27982
rect 18508 27134 18510 27186
rect 18562 27134 18564 27186
rect 18508 27122 18564 27134
rect 18620 27524 18676 27534
rect 18620 27074 18676 27468
rect 18620 27022 18622 27074
rect 18674 27022 18676 27074
rect 18620 27010 18676 27022
rect 17724 26852 17780 26862
rect 18396 26852 18564 26908
rect 17724 26850 18004 26852
rect 17724 26798 17726 26850
rect 17778 26798 18004 26850
rect 17724 26796 18004 26798
rect 17724 26786 17780 26796
rect 17948 26292 18004 26796
rect 18060 26292 18116 26302
rect 17948 26290 18116 26292
rect 17948 26238 18062 26290
rect 18114 26238 18116 26290
rect 17948 26236 18116 26238
rect 17948 25506 18004 25518
rect 17948 25454 17950 25506
rect 18002 25454 18004 25506
rect 17724 24612 17780 24622
rect 17724 24518 17780 24556
rect 17948 24612 18004 25454
rect 17948 24052 18004 24556
rect 17948 23986 18004 23996
rect 18060 23154 18116 26236
rect 18396 26178 18452 26190
rect 18396 26126 18398 26178
rect 18450 26126 18452 26178
rect 18172 26068 18228 26078
rect 18172 23378 18228 26012
rect 18396 24724 18452 26126
rect 18508 25618 18564 26852
rect 18732 26516 18788 27916
rect 18956 26516 19012 31836
rect 19068 31444 19124 33068
rect 19180 32450 19236 33180
rect 19292 32900 19348 33294
rect 20524 33236 20580 33246
rect 20300 33124 20356 33134
rect 20300 33030 20356 33068
rect 20412 33124 20468 33134
rect 20524 33124 20580 33180
rect 20412 33122 20580 33124
rect 20412 33070 20414 33122
rect 20466 33070 20580 33122
rect 20412 33068 20580 33070
rect 20636 33234 20692 33628
rect 20860 33460 20916 33470
rect 20636 33182 20638 33234
rect 20690 33182 20692 33234
rect 20636 33124 20692 33182
rect 20748 33236 20804 33246
rect 20860 33236 20916 33404
rect 21420 33458 21476 34076
rect 21644 33796 21700 37436
rect 22092 36932 22148 36942
rect 22092 36594 22148 36876
rect 22092 36542 22094 36594
rect 22146 36542 22148 36594
rect 22092 36530 22148 36542
rect 23660 36596 23716 36606
rect 23772 36596 23828 39200
rect 23660 36594 24612 36596
rect 23660 36542 23662 36594
rect 23714 36542 24612 36594
rect 23660 36540 24612 36542
rect 23660 36530 23716 36540
rect 24556 36482 24612 36540
rect 24556 36430 24558 36482
rect 24610 36430 24612 36482
rect 24556 36418 24612 36430
rect 24780 36484 24836 36494
rect 22092 36372 22148 36382
rect 21868 35700 21924 35710
rect 21868 34916 21924 35644
rect 21868 34850 21924 34860
rect 22092 34580 22148 36316
rect 24108 36372 24164 36382
rect 24108 36278 24164 36316
rect 24780 35922 24836 36428
rect 24780 35870 24782 35922
rect 24834 35870 24836 35922
rect 24780 35858 24836 35870
rect 25116 36482 25172 36494
rect 25116 36430 25118 36482
rect 25170 36430 25172 36482
rect 22316 35586 22372 35598
rect 22316 35534 22318 35586
rect 22370 35534 22372 35586
rect 22204 34804 22260 34814
rect 22204 34710 22260 34748
rect 22092 34524 22260 34580
rect 21420 33406 21422 33458
rect 21474 33406 21476 33458
rect 21420 33394 21476 33406
rect 21532 33740 21700 33796
rect 21868 34018 21924 34030
rect 21868 33966 21870 34018
rect 21922 33966 21924 34018
rect 20748 33234 20916 33236
rect 20748 33182 20750 33234
rect 20802 33182 20916 33234
rect 20748 33180 20916 33182
rect 20748 33170 20804 33180
rect 20412 33058 20468 33068
rect 20636 33058 20692 33068
rect 20532 32956 20796 32966
rect 20588 32900 20636 32956
rect 20692 32900 20740 32956
rect 20532 32890 20796 32900
rect 19292 32834 19348 32844
rect 19516 32674 19572 32686
rect 19516 32622 19518 32674
rect 19570 32622 19572 32674
rect 19292 32564 19348 32574
rect 19292 32470 19348 32508
rect 19180 32398 19182 32450
rect 19234 32398 19236 32450
rect 19180 32386 19236 32398
rect 19516 32452 19572 32622
rect 19964 32564 20020 32574
rect 19516 32386 19572 32396
rect 19740 32508 19964 32564
rect 19068 31378 19124 31388
rect 19404 31332 19460 31342
rect 19068 30324 19124 30334
rect 19068 30230 19124 30268
rect 19292 30212 19348 30222
rect 19180 30100 19236 30110
rect 19068 29988 19124 29998
rect 19068 29426 19124 29932
rect 19180 29650 19236 30044
rect 19180 29598 19182 29650
rect 19234 29598 19236 29650
rect 19180 29586 19236 29598
rect 19068 29374 19070 29426
rect 19122 29374 19124 29426
rect 19068 29362 19124 29374
rect 19292 29426 19348 30156
rect 19404 29764 19460 31276
rect 19628 31106 19684 31118
rect 19628 31054 19630 31106
rect 19682 31054 19684 31106
rect 19516 30994 19572 31006
rect 19516 30942 19518 30994
rect 19570 30942 19572 30994
rect 19516 30212 19572 30942
rect 19516 30118 19572 30156
rect 19628 29988 19684 31054
rect 19628 29922 19684 29932
rect 19404 29708 19572 29764
rect 19292 29374 19294 29426
rect 19346 29374 19348 29426
rect 19292 29362 19348 29374
rect 19292 29092 19348 29102
rect 19180 29036 19292 29092
rect 19068 28642 19124 28654
rect 19068 28590 19070 28642
rect 19122 28590 19124 28642
rect 19068 27860 19124 28590
rect 19068 27794 19124 27804
rect 19068 27188 19124 27198
rect 19180 27188 19236 29036
rect 19292 29026 19348 29036
rect 19292 28084 19348 28094
rect 19292 27636 19348 28028
rect 19292 27570 19348 27580
rect 19068 27186 19236 27188
rect 19068 27134 19070 27186
rect 19122 27134 19236 27186
rect 19068 27132 19236 27134
rect 19068 27122 19124 27132
rect 18620 26460 18788 26516
rect 18844 26460 19012 26516
rect 18620 25956 18676 26460
rect 18732 26180 18788 26190
rect 18732 26086 18788 26124
rect 18732 25956 18788 25966
rect 18620 25900 18732 25956
rect 18732 25890 18788 25900
rect 18508 25566 18510 25618
rect 18562 25566 18564 25618
rect 18508 25554 18564 25566
rect 18732 24724 18788 24734
rect 18396 24668 18732 24724
rect 18732 24630 18788 24668
rect 18732 24276 18788 24286
rect 18396 24052 18452 24062
rect 18452 23996 18564 24052
rect 18396 23986 18452 23996
rect 18508 23938 18564 23996
rect 18508 23886 18510 23938
rect 18562 23886 18564 23938
rect 18508 23874 18564 23886
rect 18172 23326 18174 23378
rect 18226 23326 18228 23378
rect 18172 23314 18228 23326
rect 18060 23102 18062 23154
rect 18114 23102 18116 23154
rect 18060 23090 18116 23102
rect 18732 23154 18788 24220
rect 18732 23102 18734 23154
rect 18786 23102 18788 23154
rect 18732 23090 18788 23102
rect 18172 22932 18228 22942
rect 18844 22932 18900 26460
rect 19516 26404 19572 29708
rect 19740 29540 19796 32508
rect 19964 32470 20020 32508
rect 20412 32452 20468 32462
rect 20412 32358 20468 32396
rect 20412 31890 20468 31902
rect 20412 31838 20414 31890
rect 20466 31838 20468 31890
rect 20300 31778 20356 31790
rect 20300 31726 20302 31778
rect 20354 31726 20356 31778
rect 19852 31108 19908 31118
rect 19852 31014 19908 31052
rect 20076 31108 20132 31118
rect 20076 31014 20132 31052
rect 20188 31106 20244 31118
rect 20188 31054 20190 31106
rect 20242 31054 20244 31106
rect 20076 30772 20132 30782
rect 20076 30434 20132 30716
rect 20188 30548 20244 31054
rect 20188 30482 20244 30492
rect 20076 30382 20078 30434
rect 20130 30382 20132 30434
rect 20076 30370 20132 30382
rect 20188 30212 20244 30222
rect 19740 29484 20020 29540
rect 19740 29316 19796 29326
rect 19740 29222 19796 29260
rect 19628 28644 19684 28654
rect 19628 28642 19908 28644
rect 19628 28590 19630 28642
rect 19682 28590 19908 28642
rect 19628 28588 19908 28590
rect 19628 28578 19684 28588
rect 19852 28082 19908 28588
rect 19852 28030 19854 28082
rect 19906 28030 19908 28082
rect 19852 28018 19908 28030
rect 19628 27858 19684 27870
rect 19628 27806 19630 27858
rect 19682 27806 19684 27858
rect 19628 27524 19684 27806
rect 19628 27458 19684 27468
rect 19964 27300 20020 29484
rect 20188 28754 20244 30156
rect 20300 30100 20356 31726
rect 20412 31218 20468 31838
rect 20532 31388 20796 31398
rect 20588 31332 20636 31388
rect 20692 31332 20740 31388
rect 20532 31322 20796 31332
rect 20412 31166 20414 31218
rect 20466 31166 20468 31218
rect 20412 31154 20468 31166
rect 20748 30882 20804 30894
rect 20748 30830 20750 30882
rect 20802 30830 20804 30882
rect 20748 30548 20804 30830
rect 20748 30482 20804 30492
rect 20300 30034 20356 30044
rect 20524 30100 20580 30110
rect 20524 30006 20580 30044
rect 20532 29820 20796 29830
rect 20588 29764 20636 29820
rect 20692 29764 20740 29820
rect 20532 29754 20796 29764
rect 20300 29652 20356 29662
rect 20300 29538 20356 29596
rect 20748 29652 20804 29662
rect 20748 29558 20804 29596
rect 20300 29486 20302 29538
rect 20354 29486 20356 29538
rect 20300 29474 20356 29486
rect 20412 29540 20468 29550
rect 20636 29540 20692 29550
rect 20412 29538 20580 29540
rect 20412 29486 20414 29538
rect 20466 29486 20580 29538
rect 20412 29484 20580 29486
rect 20412 29474 20468 29484
rect 20524 29204 20580 29484
rect 20636 29446 20692 29484
rect 20860 29316 20916 33180
rect 21532 33234 21588 33740
rect 21868 33460 21924 33966
rect 21868 33394 21924 33404
rect 22092 33346 22148 33358
rect 22092 33294 22094 33346
rect 22146 33294 22148 33346
rect 21532 33182 21534 33234
rect 21586 33182 21588 33234
rect 21308 33122 21364 33134
rect 21308 33070 21310 33122
rect 21362 33070 21364 33122
rect 20972 33012 21028 33022
rect 20972 32788 21028 32956
rect 20972 32694 21028 32732
rect 21308 32676 21364 33070
rect 21532 33012 21588 33182
rect 21644 33236 21700 33246
rect 21644 33142 21700 33180
rect 22092 33124 22148 33294
rect 22092 33058 22148 33068
rect 21532 32946 21588 32956
rect 21308 32610 21364 32620
rect 21420 30994 21476 31006
rect 21420 30942 21422 30994
rect 21474 30942 21476 30994
rect 21308 30884 21364 30894
rect 21308 30548 21364 30828
rect 21420 30772 21476 30942
rect 21420 30706 21476 30716
rect 21308 30492 21476 30548
rect 21196 30100 21252 30110
rect 20524 29138 20580 29148
rect 20636 29260 20916 29316
rect 20972 29538 21028 29550
rect 20972 29486 20974 29538
rect 21026 29486 21028 29538
rect 20636 28980 20692 29260
rect 20188 28702 20190 28754
rect 20242 28702 20244 28754
rect 20188 28690 20244 28702
rect 20300 28924 20692 28980
rect 20748 28980 20804 28990
rect 20076 27972 20132 27982
rect 20076 27878 20132 27916
rect 20188 27858 20244 27870
rect 20188 27806 20190 27858
rect 20242 27806 20244 27858
rect 20188 27412 20244 27806
rect 20188 27346 20244 27356
rect 19964 27244 20132 27300
rect 19964 27076 20020 27086
rect 19852 26516 19908 26526
rect 19740 26460 19852 26516
rect 19516 26348 19684 26404
rect 19404 26292 19460 26302
rect 19404 26198 19460 26236
rect 19180 26178 19236 26190
rect 19628 26180 19684 26348
rect 19180 26126 19182 26178
rect 19234 26126 19236 26178
rect 19068 26068 19124 26078
rect 19068 25974 19124 26012
rect 18956 25956 19012 25966
rect 18956 23548 19012 25900
rect 19180 24722 19236 26126
rect 19516 26124 19684 26180
rect 19180 24670 19182 24722
rect 19234 24670 19236 24722
rect 19180 24658 19236 24670
rect 19404 24724 19460 24734
rect 19404 24630 19460 24668
rect 19068 24500 19124 24510
rect 19068 23938 19124 24444
rect 19068 23886 19070 23938
rect 19122 23886 19124 23938
rect 19068 23874 19124 23886
rect 18956 23492 19236 23548
rect 18172 22370 18228 22876
rect 18508 22876 18900 22932
rect 19068 23268 19124 23278
rect 18172 22318 18174 22370
rect 18226 22318 18228 22370
rect 18172 22306 18228 22318
rect 18284 22484 18340 22494
rect 18284 22370 18340 22428
rect 18284 22318 18286 22370
rect 18338 22318 18340 22370
rect 18284 22306 18340 22318
rect 18508 22370 18564 22876
rect 18508 22318 18510 22370
rect 18562 22318 18564 22370
rect 18508 22306 18564 22318
rect 18732 22596 18788 22606
rect 18732 22370 18788 22540
rect 18732 22318 18734 22370
rect 18786 22318 18788 22370
rect 18732 22306 18788 22318
rect 18396 22148 18452 22158
rect 18396 22054 18452 22092
rect 18396 21924 18452 21934
rect 18284 21586 18340 21598
rect 18284 21534 18286 21586
rect 18338 21534 18340 21586
rect 17836 21474 17892 21486
rect 17836 21422 17838 21474
rect 17890 21422 17892 21474
rect 17836 21140 17892 21422
rect 17836 21074 17892 21084
rect 18284 21364 18340 21534
rect 17836 20916 17892 20926
rect 17836 20822 17892 20860
rect 18284 20804 18340 21308
rect 18284 20738 18340 20748
rect 18396 21586 18452 21868
rect 18508 21812 18564 21822
rect 18508 21718 18564 21756
rect 18732 21700 18788 21710
rect 18732 21606 18788 21644
rect 18396 21534 18398 21586
rect 18450 21534 18452 21586
rect 18284 20580 18340 20590
rect 18396 20580 18452 21534
rect 18620 21586 18676 21598
rect 18620 21534 18622 21586
rect 18674 21534 18676 21586
rect 18620 21140 18676 21534
rect 18620 21074 18676 21084
rect 18508 20580 18564 20590
rect 18396 20524 18508 20580
rect 18284 20486 18340 20524
rect 17948 19908 18004 19918
rect 17948 19906 18116 19908
rect 17948 19854 17950 19906
rect 18002 19854 18116 19906
rect 17948 19852 18116 19854
rect 17948 19842 18004 19852
rect 17836 19794 17892 19806
rect 17836 19742 17838 19794
rect 17890 19742 17892 19794
rect 17836 19684 17892 19742
rect 17836 19628 18004 19684
rect 16828 18498 16884 18508
rect 16940 18956 17108 19012
rect 17164 19516 17668 19572
rect 16828 18340 16884 18350
rect 16940 18340 16996 18956
rect 17164 18788 17220 19516
rect 16884 18284 16996 18340
rect 17052 18732 17220 18788
rect 17276 19234 17332 19246
rect 17276 19182 17278 19234
rect 17330 19182 17332 19234
rect 16828 18246 16884 18284
rect 17052 18116 17108 18732
rect 17276 18452 17332 19182
rect 17836 19124 17892 19134
rect 17724 19068 17836 19124
rect 16716 17726 16718 17778
rect 16770 17726 16772 17778
rect 16716 17714 16772 17726
rect 16828 18060 17108 18116
rect 17164 18396 17332 18452
rect 17388 18900 17444 18910
rect 17388 18450 17444 18844
rect 17388 18398 17390 18450
rect 17442 18398 17444 18450
rect 17164 18228 17220 18396
rect 17388 18386 17444 18398
rect 17724 18562 17780 19068
rect 17836 19058 17892 19068
rect 17724 18510 17726 18562
rect 17778 18510 17780 18562
rect 17724 18228 17780 18510
rect 16492 17554 16660 17556
rect 16492 17502 16494 17554
rect 16546 17502 16660 17554
rect 16492 17500 16660 17502
rect 16716 17556 16772 17566
rect 16492 17490 16548 17500
rect 16716 17462 16772 17500
rect 16380 17276 16548 17332
rect 16268 16996 16324 17006
rect 16268 16902 16324 16940
rect 16156 16882 16212 16894
rect 16156 16830 16158 16882
rect 16210 16830 16212 16882
rect 16156 16210 16212 16830
rect 16380 16884 16436 16894
rect 16380 16790 16436 16828
rect 16156 16158 16158 16210
rect 16210 16158 16212 16210
rect 16156 16146 16212 16158
rect 16156 15988 16212 15998
rect 16044 15986 16212 15988
rect 16044 15934 16158 15986
rect 16210 15934 16212 15986
rect 16044 15932 16212 15934
rect 16156 15922 16212 15932
rect 16268 15876 16324 15886
rect 16492 15876 16548 17276
rect 15484 15820 15876 15876
rect 15708 15540 15764 15550
rect 15372 13244 15540 13300
rect 14588 12738 15092 12740
rect 14588 12686 15038 12738
rect 15090 12686 15092 12738
rect 14588 12684 15092 12686
rect 14588 11394 14644 12684
rect 15036 12674 15092 12684
rect 15260 13188 15316 13198
rect 14588 11342 14590 11394
rect 14642 11342 14644 11394
rect 14364 6738 14420 6748
rect 14476 9828 14532 9838
rect 14476 8260 14532 9772
rect 14588 9268 14644 11342
rect 15148 11844 15204 11854
rect 14924 9268 14980 9278
rect 14588 9266 14980 9268
rect 14588 9214 14926 9266
rect 14978 9214 14980 9266
rect 14588 9212 14980 9214
rect 14924 9202 14980 9212
rect 14588 8260 14644 8270
rect 14476 8258 14644 8260
rect 14476 8206 14590 8258
rect 14642 8206 14644 8258
rect 14476 8204 14644 8206
rect 13692 6692 13748 6702
rect 13580 6690 13748 6692
rect 13580 6638 13694 6690
rect 13746 6638 13748 6690
rect 13580 6636 13748 6638
rect 13692 6626 13748 6636
rect 13468 6468 13524 6478
rect 13468 6466 13748 6468
rect 13468 6414 13470 6466
rect 13522 6414 13748 6466
rect 13468 6412 13748 6414
rect 13468 6402 13524 6412
rect 13132 6038 13188 6076
rect 13580 5908 13636 5918
rect 13580 5794 13636 5852
rect 13580 5742 13582 5794
rect 13634 5742 13636 5794
rect 13580 5730 13636 5742
rect 12964 5180 13076 5236
rect 12908 5142 12964 5180
rect 12796 5012 12852 5022
rect 12796 4562 12852 4956
rect 13580 4900 13636 4910
rect 12796 4510 12798 4562
rect 12850 4510 12852 4562
rect 12796 4498 12852 4510
rect 13132 4898 13636 4900
rect 13132 4846 13582 4898
rect 13634 4846 13636 4898
rect 13132 4844 13636 4846
rect 13132 4450 13188 4844
rect 13580 4834 13636 4844
rect 13692 4788 13748 6412
rect 14252 6132 14308 6142
rect 14252 5684 14308 6076
rect 14252 5618 14308 5628
rect 13916 5236 13972 5246
rect 14476 5236 14532 8204
rect 14588 8194 14644 8204
rect 15148 7252 15204 11788
rect 15260 11394 15316 13132
rect 15484 13076 15540 13244
rect 15708 13188 15764 15484
rect 15820 15148 15876 15820
rect 16268 15874 16548 15876
rect 16268 15822 16270 15874
rect 16322 15822 16548 15874
rect 16268 15820 16548 15822
rect 16716 17220 16772 17230
rect 16156 15428 16212 15438
rect 16156 15334 16212 15372
rect 15820 15092 15988 15148
rect 15932 15090 15988 15092
rect 15932 15038 15934 15090
rect 15986 15038 15988 15090
rect 15932 15026 15988 15038
rect 15932 14196 15988 14206
rect 15932 13858 15988 14140
rect 15932 13806 15934 13858
rect 15986 13806 15988 13858
rect 15932 13794 15988 13806
rect 15708 13122 15764 13132
rect 15820 13746 15876 13758
rect 15820 13694 15822 13746
rect 15874 13694 15876 13746
rect 15372 13020 15540 13076
rect 15372 11508 15428 13020
rect 15484 12738 15540 12750
rect 15484 12686 15486 12738
rect 15538 12686 15540 12738
rect 15484 11844 15540 12686
rect 15820 12740 15876 13694
rect 16044 13748 16100 13758
rect 16044 13654 16100 13692
rect 16268 13524 16324 15820
rect 16716 15652 16772 17164
rect 16828 17106 16884 18060
rect 17164 17892 17220 18172
rect 17164 17826 17220 17836
rect 17388 18172 17780 18228
rect 17836 18900 17892 18910
rect 17388 17890 17444 18172
rect 17388 17838 17390 17890
rect 17442 17838 17444 17890
rect 17388 17826 17444 17838
rect 17500 17892 17556 17902
rect 17500 17798 17556 17836
rect 17724 17892 17780 17902
rect 17836 17892 17892 18844
rect 17724 17890 17892 17892
rect 17724 17838 17726 17890
rect 17778 17838 17892 17890
rect 17724 17836 17892 17838
rect 17724 17826 17780 17836
rect 17948 17668 18004 19628
rect 18060 19236 18116 19852
rect 18172 19460 18228 19470
rect 18172 19458 18452 19460
rect 18172 19406 18174 19458
rect 18226 19406 18452 19458
rect 18172 19404 18452 19406
rect 18172 19394 18228 19404
rect 18396 19236 18452 19404
rect 18060 19180 18228 19236
rect 18060 18450 18116 18462
rect 18060 18398 18062 18450
rect 18114 18398 18116 18450
rect 18060 18004 18116 18398
rect 18060 17938 18116 17948
rect 18172 17780 18228 19180
rect 18284 19124 18340 19134
rect 18284 19030 18340 19068
rect 18396 18900 18452 19180
rect 18396 18834 18452 18844
rect 18508 18676 18564 20524
rect 18956 20580 19012 20590
rect 18956 20486 19012 20524
rect 18732 20468 18788 20478
rect 18620 19236 18676 19246
rect 18620 19142 18676 19180
rect 18732 19012 18788 20412
rect 19068 20468 19124 23212
rect 19068 20402 19124 20412
rect 19180 20132 19236 23492
rect 19404 22484 19460 22494
rect 19516 22484 19572 26124
rect 19740 25620 19796 26460
rect 19852 26450 19908 26460
rect 19852 26292 19908 26302
rect 19852 26198 19908 26236
rect 19852 25620 19908 25630
rect 19740 25618 19908 25620
rect 19740 25566 19854 25618
rect 19906 25566 19908 25618
rect 19740 25564 19908 25566
rect 19852 25554 19908 25564
rect 19740 24948 19796 24958
rect 19628 24834 19684 24846
rect 19628 24782 19630 24834
rect 19682 24782 19684 24834
rect 19628 24612 19684 24782
rect 19740 24836 19796 24892
rect 19740 24834 19908 24836
rect 19740 24782 19742 24834
rect 19794 24782 19908 24834
rect 19740 24780 19908 24782
rect 19740 24770 19796 24780
rect 19628 24556 19796 24612
rect 19628 24388 19684 24398
rect 19628 23378 19684 24332
rect 19628 23326 19630 23378
rect 19682 23326 19684 23378
rect 19628 23314 19684 23326
rect 19740 23268 19796 24556
rect 19852 24276 19908 24780
rect 19852 24210 19908 24220
rect 19964 24164 20020 27020
rect 20076 26292 20132 27244
rect 20076 26226 20132 26236
rect 20076 26068 20132 26078
rect 20076 25506 20132 26012
rect 20076 25454 20078 25506
rect 20130 25454 20132 25506
rect 20076 25442 20132 25454
rect 20188 24836 20244 24846
rect 20188 24610 20244 24780
rect 20300 24722 20356 28924
rect 20748 28754 20804 28924
rect 20972 28868 21028 29486
rect 20972 28802 21028 28812
rect 21084 29426 21140 29438
rect 21084 29374 21086 29426
rect 21138 29374 21140 29426
rect 20748 28702 20750 28754
rect 20802 28702 20804 28754
rect 20748 28690 20804 28702
rect 21084 28756 21140 29374
rect 21084 28690 21140 28700
rect 20860 28644 20916 28654
rect 20532 28252 20796 28262
rect 20588 28196 20636 28252
rect 20692 28196 20740 28252
rect 20532 28186 20796 28196
rect 20748 28084 20804 28094
rect 20748 27858 20804 28028
rect 20748 27806 20750 27858
rect 20802 27806 20804 27858
rect 20524 27748 20580 27758
rect 20524 27188 20580 27692
rect 20524 27122 20580 27132
rect 20748 27076 20804 27806
rect 20748 27010 20804 27020
rect 20532 26684 20796 26694
rect 20588 26628 20636 26684
rect 20692 26628 20740 26684
rect 20532 26618 20796 26628
rect 20636 26402 20692 26414
rect 20636 26350 20638 26402
rect 20690 26350 20692 26402
rect 20636 26068 20692 26350
rect 20636 26002 20692 26012
rect 20748 25508 20804 25518
rect 20748 25414 20804 25452
rect 20532 25116 20796 25126
rect 20588 25060 20636 25116
rect 20692 25060 20740 25116
rect 20532 25050 20796 25060
rect 20300 24670 20302 24722
rect 20354 24670 20356 24722
rect 20300 24658 20356 24670
rect 20524 24722 20580 24734
rect 20524 24670 20526 24722
rect 20578 24670 20580 24722
rect 20188 24558 20190 24610
rect 20242 24558 20244 24610
rect 19964 24108 20132 24164
rect 19852 24050 19908 24062
rect 19852 23998 19854 24050
rect 19906 23998 19908 24050
rect 19852 23380 19908 23998
rect 19852 23324 20020 23380
rect 19740 23202 19796 23212
rect 19460 22428 19572 22484
rect 19852 23156 19908 23166
rect 19852 22596 19908 23100
rect 19852 22482 19908 22540
rect 19852 22430 19854 22482
rect 19906 22430 19908 22482
rect 19404 22390 19460 22428
rect 19852 22418 19908 22430
rect 19964 22036 20020 23324
rect 19852 21980 20020 22036
rect 19292 21812 19348 21822
rect 19348 21756 19572 21812
rect 19292 21746 19348 21756
rect 19516 21698 19572 21756
rect 19516 21646 19518 21698
rect 19570 21646 19572 21698
rect 19516 21634 19572 21646
rect 19292 21588 19348 21598
rect 19292 21494 19348 21532
rect 19404 21586 19460 21598
rect 19404 21534 19406 21586
rect 19458 21534 19460 21586
rect 19404 21476 19460 21534
rect 19404 21410 19460 21420
rect 19628 21140 19684 21150
rect 19292 20580 19348 20590
rect 19404 20580 19460 20590
rect 19292 20578 19404 20580
rect 19292 20526 19294 20578
rect 19346 20526 19404 20578
rect 19292 20524 19404 20526
rect 19292 20514 19348 20524
rect 19180 20076 19348 20132
rect 18956 19122 19012 19134
rect 18956 19070 18958 19122
rect 19010 19070 19012 19122
rect 18172 17714 18228 17724
rect 18396 18620 18564 18676
rect 18620 18956 18788 19012
rect 18844 19010 18900 19022
rect 18844 18958 18846 19010
rect 18898 18958 18900 19010
rect 17388 17612 18004 17668
rect 16828 17054 16830 17106
rect 16882 17054 16884 17106
rect 16828 17042 16884 17054
rect 16940 17554 16996 17566
rect 16940 17502 16942 17554
rect 16994 17502 16996 17554
rect 16828 16212 16884 16222
rect 16828 15764 16884 16156
rect 16940 15988 16996 17502
rect 17052 17444 17108 17454
rect 17052 16098 17108 17388
rect 17052 16046 17054 16098
rect 17106 16046 17108 16098
rect 17052 16034 17108 16046
rect 17164 16884 17220 16894
rect 16940 15922 16996 15932
rect 16828 15708 17108 15764
rect 16716 15596 16996 15652
rect 16604 15316 16660 15326
rect 16604 15202 16660 15260
rect 16604 15150 16606 15202
rect 16658 15150 16660 15202
rect 16492 15090 16548 15102
rect 16492 15038 16494 15090
rect 16546 15038 16548 15090
rect 16492 13970 16548 15038
rect 16492 13918 16494 13970
rect 16546 13918 16548 13970
rect 16492 13906 16548 13918
rect 15932 13468 16324 13524
rect 15932 12962 15988 13468
rect 15932 12910 15934 12962
rect 15986 12910 15988 12962
rect 15932 12898 15988 12910
rect 16268 13076 16324 13086
rect 16268 12962 16324 13020
rect 16268 12910 16270 12962
rect 16322 12910 16324 12962
rect 16268 12898 16324 12910
rect 16380 12962 16436 12974
rect 16380 12910 16382 12962
rect 16434 12910 16436 12962
rect 15820 12674 15876 12684
rect 16044 12738 16100 12750
rect 16044 12686 16046 12738
rect 16098 12686 16100 12738
rect 15484 11778 15540 11788
rect 15708 12180 15764 12190
rect 15708 11508 15764 12124
rect 15820 12068 15876 12078
rect 15820 11974 15876 12012
rect 15372 11452 15652 11508
rect 15708 11452 15876 11508
rect 15260 11342 15262 11394
rect 15314 11342 15316 11394
rect 15260 11330 15316 11342
rect 15484 11284 15540 11294
rect 15484 11190 15540 11228
rect 15372 11170 15428 11182
rect 15372 11118 15374 11170
rect 15426 11118 15428 11170
rect 15372 9940 15428 11118
rect 15484 10610 15540 10622
rect 15484 10558 15486 10610
rect 15538 10558 15540 10610
rect 15484 10276 15540 10558
rect 15484 10210 15540 10220
rect 15372 9874 15428 9884
rect 15596 8428 15652 11452
rect 15708 10500 15764 10510
rect 15708 10406 15764 10444
rect 15708 10276 15764 10286
rect 15820 10276 15876 11452
rect 15932 11394 15988 11406
rect 15932 11342 15934 11394
rect 15986 11342 15988 11394
rect 15932 10836 15988 11342
rect 16044 11284 16100 12686
rect 16156 12740 16212 12750
rect 16156 12646 16212 12684
rect 16268 12068 16324 12078
rect 16268 11954 16324 12012
rect 16268 11902 16270 11954
rect 16322 11902 16324 11954
rect 16268 11890 16324 11902
rect 16380 11396 16436 12910
rect 16604 12852 16660 15150
rect 16716 14756 16772 14766
rect 16716 14530 16772 14700
rect 16716 14478 16718 14530
rect 16770 14478 16772 14530
rect 16716 14466 16772 14478
rect 16828 14532 16884 14542
rect 16492 12796 16660 12852
rect 16492 12180 16548 12796
rect 16492 12114 16548 12124
rect 16716 12628 16772 12638
rect 16268 11340 16436 11396
rect 16492 11506 16548 11518
rect 16492 11454 16494 11506
rect 16546 11454 16548 11506
rect 16492 11396 16548 11454
rect 16156 11284 16212 11294
rect 16044 11282 16212 11284
rect 16044 11230 16158 11282
rect 16210 11230 16212 11282
rect 16044 11228 16212 11230
rect 15932 10770 15988 10780
rect 16044 10388 16100 10398
rect 16044 10294 16100 10332
rect 15764 10220 15876 10276
rect 15708 10210 15764 10220
rect 16156 8596 16212 11228
rect 16268 9940 16324 11340
rect 16492 11330 16548 11340
rect 16716 11394 16772 12572
rect 16828 12516 16884 14476
rect 16940 14306 16996 15596
rect 16940 14254 16942 14306
rect 16994 14254 16996 14306
rect 16940 13972 16996 14254
rect 16940 13906 16996 13916
rect 16940 13076 16996 13086
rect 17052 13076 17108 15708
rect 17164 14642 17220 16828
rect 17388 15652 17444 17612
rect 18284 17554 18340 17566
rect 18284 17502 18286 17554
rect 18338 17502 18340 17554
rect 17612 16882 17668 16894
rect 17612 16830 17614 16882
rect 17666 16830 17668 16882
rect 17612 16324 17668 16830
rect 18060 16770 18116 16782
rect 18060 16718 18062 16770
rect 18114 16718 18116 16770
rect 18060 16436 18116 16718
rect 18284 16548 18340 17502
rect 18396 17220 18452 18620
rect 18620 18452 18676 18956
rect 18620 18386 18676 18396
rect 18508 18340 18564 18350
rect 18508 17556 18564 18284
rect 18620 18226 18676 18238
rect 18620 18174 18622 18226
rect 18674 18174 18676 18226
rect 18620 17780 18676 18174
rect 18620 17724 18788 17780
rect 18620 17556 18676 17566
rect 18508 17554 18676 17556
rect 18508 17502 18622 17554
rect 18674 17502 18676 17554
rect 18508 17500 18676 17502
rect 18620 17490 18676 17500
rect 18396 17154 18452 17164
rect 18732 16996 18788 17724
rect 18844 17778 18900 18958
rect 18956 18676 19012 19070
rect 18956 18610 19012 18620
rect 19068 18564 19124 18574
rect 19068 18470 19124 18508
rect 18844 17726 18846 17778
rect 18898 17726 18900 17778
rect 18844 17714 18900 17726
rect 18956 18452 19012 18462
rect 18844 17444 18900 17454
rect 18844 17350 18900 17388
rect 18844 16996 18900 17006
rect 18732 16940 18844 16996
rect 18844 16930 18900 16940
rect 18844 16772 18900 16782
rect 18620 16770 18900 16772
rect 18620 16718 18846 16770
rect 18898 16718 18900 16770
rect 18620 16716 18900 16718
rect 18284 16492 18564 16548
rect 18060 16380 18452 16436
rect 17500 16268 18340 16324
rect 17500 16210 17556 16268
rect 17500 16158 17502 16210
rect 17554 16158 17556 16210
rect 17500 16146 17556 16158
rect 17836 16100 17892 16110
rect 17164 14590 17166 14642
rect 17218 14590 17220 14642
rect 17164 14578 17220 14590
rect 17276 15596 17444 15652
rect 17612 16098 17892 16100
rect 17612 16046 17838 16098
rect 17890 16046 17892 16098
rect 17612 16044 17892 16046
rect 17276 14532 17332 15596
rect 17612 15540 17668 16044
rect 17836 16034 17892 16044
rect 17500 15484 17668 15540
rect 17948 15988 18004 15998
rect 17388 15426 17444 15438
rect 17388 15374 17390 15426
rect 17442 15374 17444 15426
rect 17388 14756 17444 15374
rect 17388 14690 17444 14700
rect 17388 14532 17444 14542
rect 17276 14530 17444 14532
rect 17276 14478 17390 14530
rect 17442 14478 17444 14530
rect 17276 14476 17444 14478
rect 17164 14308 17220 14318
rect 17164 14214 17220 14252
rect 17388 13746 17444 14476
rect 17500 14532 17556 15484
rect 17612 15314 17668 15326
rect 17612 15262 17614 15314
rect 17666 15262 17668 15314
rect 17612 14980 17668 15262
rect 17948 15314 18004 15932
rect 17948 15262 17950 15314
rect 18002 15262 18004 15314
rect 17948 15148 18004 15262
rect 18284 15314 18340 16268
rect 18284 15262 18286 15314
rect 18338 15262 18340 15314
rect 18284 15250 18340 15262
rect 17612 14914 17668 14924
rect 17724 15090 17780 15102
rect 17724 15038 17726 15090
rect 17778 15038 17780 15090
rect 17500 14466 17556 14476
rect 17724 14532 17780 15038
rect 17724 14466 17780 14476
rect 17836 15092 18004 15148
rect 18396 15204 18452 16380
rect 18396 15138 18452 15148
rect 17836 14308 17892 15092
rect 18060 14980 18116 14990
rect 17388 13694 17390 13746
rect 17442 13694 17444 13746
rect 17388 13682 17444 13694
rect 17500 14252 17892 14308
rect 17948 14308 18004 14318
rect 17500 13524 17556 14252
rect 17948 14214 18004 14252
rect 17836 13972 17892 13982
rect 17836 13878 17892 13916
rect 16996 13020 17108 13076
rect 17388 13468 17556 13524
rect 17612 13746 17668 13758
rect 17612 13694 17614 13746
rect 17666 13694 17668 13746
rect 17612 13524 17668 13694
rect 17724 13748 17780 13758
rect 17724 13654 17780 13692
rect 17948 13746 18004 13758
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 16940 12982 16996 13020
rect 17276 12852 17332 12862
rect 17388 12852 17444 13468
rect 17612 13458 17668 13468
rect 17836 13636 17892 13646
rect 17836 13188 17892 13580
rect 17276 12850 17444 12852
rect 17276 12798 17278 12850
rect 17330 12798 17444 12850
rect 17276 12796 17444 12798
rect 17500 13132 17892 13188
rect 17500 12962 17556 13132
rect 17948 13076 18004 13694
rect 18060 13636 18116 14924
rect 18396 14980 18452 14990
rect 18284 14644 18340 14654
rect 18284 14550 18340 14588
rect 18396 14530 18452 14924
rect 18396 14478 18398 14530
rect 18450 14478 18452 14530
rect 18396 14466 18452 14478
rect 18060 13570 18116 13580
rect 18172 14306 18228 14318
rect 18172 14254 18174 14306
rect 18226 14254 18228 14306
rect 18172 13188 18228 14254
rect 18284 13524 18340 13534
rect 18340 13468 18452 13524
rect 18284 13458 18340 13468
rect 18172 13132 18340 13188
rect 18284 13076 18340 13132
rect 17500 12910 17502 12962
rect 17554 12910 17556 12962
rect 17276 12740 17332 12796
rect 17276 12674 17332 12684
rect 16828 12450 16884 12460
rect 17276 11620 17332 11630
rect 17276 11506 17332 11564
rect 17276 11454 17278 11506
rect 17330 11454 17332 11506
rect 17276 11442 17332 11454
rect 16716 11342 16718 11394
rect 16770 11342 16772 11394
rect 16716 11330 16772 11342
rect 16828 11396 16884 11406
rect 16828 11302 16884 11340
rect 16940 11284 16996 11294
rect 16380 11172 16436 11182
rect 16380 11078 16436 11116
rect 16828 10052 16884 10062
rect 16940 10052 16996 11228
rect 17500 11172 17556 12910
rect 17724 13020 18228 13076
rect 17724 12850 17780 13020
rect 17724 12798 17726 12850
rect 17778 12798 17780 12850
rect 17724 12786 17780 12798
rect 17836 12852 17892 12862
rect 17836 12758 17892 12796
rect 18060 12850 18116 12862
rect 18060 12798 18062 12850
rect 18114 12798 18116 12850
rect 17948 12628 18004 12638
rect 18060 12628 18116 12798
rect 18004 12572 18116 12628
rect 17948 12562 18004 12572
rect 17612 12290 17668 12302
rect 17612 12238 17614 12290
rect 17666 12238 17668 12290
rect 17612 11620 17668 12238
rect 17612 11554 17668 11564
rect 17500 11106 17556 11116
rect 18060 11172 18116 11182
rect 17276 10836 17332 10846
rect 18060 10836 18116 11116
rect 17276 10742 17332 10780
rect 17948 10834 18116 10836
rect 17948 10782 18062 10834
rect 18114 10782 18116 10834
rect 17948 10780 18116 10782
rect 17500 10722 17556 10734
rect 17500 10670 17502 10722
rect 17554 10670 17556 10722
rect 17500 10500 17556 10670
rect 17500 10434 17556 10444
rect 17612 10610 17668 10622
rect 17612 10558 17614 10610
rect 17666 10558 17668 10610
rect 16828 10050 16996 10052
rect 16828 9998 16830 10050
rect 16882 9998 16996 10050
rect 16828 9996 16996 9998
rect 17388 10276 17444 10286
rect 17388 10050 17444 10220
rect 17388 9998 17390 10050
rect 17442 9998 17444 10050
rect 16828 9986 16884 9996
rect 16380 9940 16436 9950
rect 16716 9940 16772 9950
rect 16268 9938 16772 9940
rect 16268 9886 16382 9938
rect 16434 9886 16718 9938
rect 16770 9886 16772 9938
rect 16268 9884 16772 9886
rect 16380 9874 16436 9884
rect 16716 9874 16772 9884
rect 17388 9938 17444 9998
rect 17388 9886 17390 9938
rect 17442 9886 17444 9938
rect 17388 9874 17444 9886
rect 17612 9716 17668 10558
rect 17948 10050 18004 10780
rect 18060 10770 18116 10780
rect 17948 9998 17950 10050
rect 18002 9998 18004 10050
rect 17948 9986 18004 9998
rect 17836 9716 17892 9726
rect 17612 9660 17836 9716
rect 17836 9622 17892 9660
rect 16156 8530 16212 8540
rect 17276 8596 17332 8606
rect 17332 8540 17444 8596
rect 17276 8530 17332 8540
rect 15596 8372 15876 8428
rect 15372 8148 15428 8158
rect 15372 8146 15652 8148
rect 15372 8094 15374 8146
rect 15426 8094 15652 8146
rect 15372 8092 15652 8094
rect 15372 8082 15428 8092
rect 15596 7698 15652 8092
rect 15596 7646 15598 7698
rect 15650 7646 15652 7698
rect 15596 7634 15652 7646
rect 15148 7186 15204 7196
rect 15820 6132 15876 8372
rect 17388 8148 17444 8540
rect 17500 8372 17556 8382
rect 18172 8372 18228 13020
rect 18284 12962 18340 13020
rect 18284 12910 18286 12962
rect 18338 12910 18340 12962
rect 18284 12898 18340 12910
rect 18396 12852 18452 13468
rect 18508 12964 18564 16492
rect 18620 15314 18676 16716
rect 18844 16706 18900 16716
rect 18732 16548 18788 16558
rect 18732 16322 18788 16492
rect 18956 16436 19012 18396
rect 19180 18116 19236 18126
rect 18956 16370 19012 16380
rect 19068 17554 19124 17566
rect 19068 17502 19070 17554
rect 19122 17502 19124 17554
rect 18732 16270 18734 16322
rect 18786 16270 18788 16322
rect 18732 16258 18788 16270
rect 18956 16100 19012 16110
rect 18956 16006 19012 16044
rect 18620 15262 18622 15314
rect 18674 15262 18676 15314
rect 18620 14530 18676 15262
rect 19068 14980 19124 17502
rect 19180 16882 19236 18060
rect 19180 16830 19182 16882
rect 19234 16830 19236 16882
rect 19180 16818 19236 16830
rect 19292 16658 19348 20076
rect 19292 16606 19294 16658
rect 19346 16606 19348 16658
rect 19292 16594 19348 16606
rect 19292 16436 19348 16446
rect 19068 14914 19124 14924
rect 19180 15202 19236 15214
rect 19180 15150 19182 15202
rect 19234 15150 19236 15202
rect 18620 14478 18622 14530
rect 18674 14478 18676 14530
rect 18620 14466 18676 14478
rect 18844 14644 18900 14654
rect 18844 14418 18900 14588
rect 18956 14532 19012 14542
rect 18956 14438 19012 14476
rect 18844 14366 18846 14418
rect 18898 14366 18900 14418
rect 18844 14354 18900 14366
rect 19180 13972 19236 15150
rect 19180 13906 19236 13916
rect 18620 13188 18676 13198
rect 18620 13186 19012 13188
rect 18620 13134 18622 13186
rect 18674 13134 19012 13186
rect 18620 13132 19012 13134
rect 18620 13122 18676 13132
rect 18508 12908 18788 12964
rect 18396 12796 18564 12852
rect 18508 12738 18564 12796
rect 18508 12686 18510 12738
rect 18562 12686 18564 12738
rect 18284 12516 18340 12526
rect 18284 11844 18340 12460
rect 18284 11506 18340 11788
rect 18396 11732 18452 11742
rect 18396 11618 18452 11676
rect 18396 11566 18398 11618
rect 18450 11566 18452 11618
rect 18396 11554 18452 11566
rect 18284 11454 18286 11506
rect 18338 11454 18340 11506
rect 18284 11442 18340 11454
rect 18508 10948 18564 12686
rect 18620 12178 18676 12190
rect 18620 12126 18622 12178
rect 18674 12126 18676 12178
rect 18620 12068 18676 12126
rect 18620 12002 18676 12012
rect 18620 11284 18676 11294
rect 18620 11190 18676 11228
rect 18284 10892 18564 10948
rect 18284 8708 18340 10892
rect 18732 10836 18788 12908
rect 18844 12852 18900 12862
rect 18844 12758 18900 12796
rect 18956 12850 19012 13132
rect 18956 12798 18958 12850
rect 19010 12798 19012 12850
rect 18956 12786 19012 12798
rect 19180 12738 19236 12750
rect 19180 12686 19182 12738
rect 19234 12686 19236 12738
rect 19180 12628 19236 12686
rect 18844 12572 19236 12628
rect 18844 12178 18900 12572
rect 19292 12516 19348 16380
rect 18956 12460 19348 12516
rect 18956 12290 19012 12460
rect 19404 12404 19460 20524
rect 19516 19908 19572 19918
rect 19516 15428 19572 19852
rect 19628 18450 19684 21084
rect 19740 20580 19796 20590
rect 19740 20486 19796 20524
rect 19628 18398 19630 18450
rect 19682 18398 19684 18450
rect 19628 17556 19684 18398
rect 19740 17556 19796 17566
rect 19628 17554 19796 17556
rect 19628 17502 19742 17554
rect 19794 17502 19796 17554
rect 19628 17500 19796 17502
rect 19740 17490 19796 17500
rect 19852 17332 19908 21980
rect 19964 21812 20020 21822
rect 20076 21812 20132 24108
rect 20188 23828 20244 24558
rect 20524 23940 20580 24670
rect 20524 23874 20580 23884
rect 20188 23762 20244 23772
rect 20532 23548 20796 23558
rect 19964 21810 20132 21812
rect 19964 21758 19966 21810
rect 20018 21758 20132 21810
rect 19964 21756 20132 21758
rect 20188 23492 20244 23502
rect 20588 23492 20636 23548
rect 20692 23492 20740 23548
rect 20532 23482 20796 23492
rect 19964 21746 20020 21756
rect 20188 21252 20244 23436
rect 20300 22932 20356 22942
rect 20300 22482 20356 22876
rect 20300 22430 20302 22482
rect 20354 22430 20356 22482
rect 20300 22418 20356 22430
rect 20532 21980 20796 21990
rect 20588 21924 20636 21980
rect 20692 21924 20740 21980
rect 20532 21914 20796 21924
rect 20300 21700 20356 21710
rect 20300 21606 20356 21644
rect 20188 21186 20244 21196
rect 20636 21586 20692 21598
rect 20636 21534 20638 21586
rect 20690 21534 20692 21586
rect 20636 21028 20692 21534
rect 20636 20962 20692 20972
rect 20748 20916 20804 20926
rect 20860 20916 20916 28588
rect 21196 28532 21252 30044
rect 20972 28476 21252 28532
rect 21308 28642 21364 28654
rect 21308 28590 21310 28642
rect 21362 28590 21364 28642
rect 20972 26178 21028 28476
rect 21308 28084 21364 28590
rect 21308 28018 21364 28028
rect 21084 27860 21140 27870
rect 21084 27746 21140 27804
rect 21084 27694 21086 27746
rect 21138 27694 21140 27746
rect 21084 27682 21140 27694
rect 21420 27188 21476 30492
rect 21756 30210 21812 30222
rect 22092 30212 22148 30222
rect 21756 30158 21758 30210
rect 21810 30158 21812 30210
rect 21644 29764 21700 29774
rect 21532 29204 21588 29214
rect 21532 28084 21588 29148
rect 21644 28980 21700 29708
rect 21756 29652 21812 30158
rect 21756 29586 21812 29596
rect 21868 30210 22148 30212
rect 21868 30158 22094 30210
rect 22146 30158 22148 30210
rect 21868 30156 22148 30158
rect 21644 28642 21700 28924
rect 21644 28590 21646 28642
rect 21698 28590 21700 28642
rect 21644 28578 21700 28590
rect 21756 28084 21812 28094
rect 21532 28082 21812 28084
rect 21532 28030 21758 28082
rect 21810 28030 21812 28082
rect 21532 28028 21812 28030
rect 21756 28018 21812 28028
rect 21868 27972 21924 30156
rect 22092 30146 22148 30156
rect 21868 27878 21924 27916
rect 21980 29988 22036 29998
rect 21980 28866 22036 29932
rect 22092 29540 22148 29550
rect 22092 29446 22148 29484
rect 22204 29316 22260 34524
rect 22316 34132 22372 35534
rect 23660 35586 23716 35598
rect 23660 35534 23662 35586
rect 23714 35534 23716 35586
rect 23436 34468 23492 34478
rect 22316 34066 22372 34076
rect 22988 34132 23044 34142
rect 22988 34038 23044 34076
rect 23436 34130 23492 34412
rect 23660 34356 23716 35534
rect 25004 35140 25060 35150
rect 23660 34290 23716 34300
rect 24220 34804 24276 34814
rect 24220 34354 24276 34748
rect 24444 34692 24500 34702
rect 24444 34598 24500 34636
rect 25004 34690 25060 35084
rect 25004 34638 25006 34690
rect 25058 34638 25060 34690
rect 25004 34580 25060 34638
rect 24556 34524 25060 34580
rect 24220 34302 24222 34354
rect 24274 34302 24276 34354
rect 24220 34290 24276 34302
rect 24444 34356 24500 34366
rect 24444 34242 24500 34300
rect 24444 34190 24446 34242
rect 24498 34190 24500 34242
rect 23884 34132 23940 34142
rect 23436 34078 23438 34130
rect 23490 34078 23492 34130
rect 23436 34066 23492 34078
rect 23660 34130 23940 34132
rect 23660 34078 23886 34130
rect 23938 34078 23940 34130
rect 23660 34076 23940 34078
rect 23548 33460 23604 33470
rect 22876 33348 22932 33358
rect 22876 33122 22932 33292
rect 23548 33346 23604 33404
rect 23660 33458 23716 34076
rect 23884 34066 23940 34076
rect 24108 34130 24164 34142
rect 24108 34078 24110 34130
rect 24162 34078 24164 34130
rect 24108 34020 24164 34078
rect 24108 33954 24164 33964
rect 23660 33406 23662 33458
rect 23714 33406 23716 33458
rect 23660 33394 23716 33406
rect 23548 33294 23550 33346
rect 23602 33294 23604 33346
rect 23548 33282 23604 33294
rect 23324 33124 23380 33134
rect 22876 33070 22878 33122
rect 22930 33070 22932 33122
rect 22876 33012 22932 33070
rect 22540 32676 22596 32686
rect 22540 32450 22596 32620
rect 22540 32398 22542 32450
rect 22594 32398 22596 32450
rect 22428 31778 22484 31790
rect 22428 31726 22430 31778
rect 22482 31726 22484 31778
rect 22428 30436 22484 31726
rect 22428 30370 22484 30380
rect 22540 29988 22596 32398
rect 22876 31948 22932 32956
rect 22988 33068 23324 33124
rect 22988 32786 23044 33068
rect 23324 33030 23380 33068
rect 23772 33122 23828 33134
rect 23772 33070 23774 33122
rect 23826 33070 23828 33122
rect 23772 33012 23828 33070
rect 24332 33124 24388 33134
rect 24332 33030 24388 33068
rect 23772 32946 23828 32956
rect 22988 32734 22990 32786
rect 23042 32734 23044 32786
rect 22988 32722 23044 32734
rect 23660 32676 23716 32686
rect 23660 32674 24052 32676
rect 23660 32622 23662 32674
rect 23714 32622 24052 32674
rect 23660 32620 24052 32622
rect 23660 32610 23716 32620
rect 22652 31892 22932 31948
rect 23660 32450 23716 32462
rect 23660 32398 23662 32450
rect 23714 32398 23716 32450
rect 23324 31892 23380 31902
rect 22652 31556 22708 31892
rect 23324 31798 23380 31836
rect 22764 31780 22820 31790
rect 22764 31686 22820 31724
rect 23548 31778 23604 31790
rect 23548 31726 23550 31778
rect 23602 31726 23604 31778
rect 22876 31668 22932 31678
rect 22876 31666 23044 31668
rect 22876 31614 22878 31666
rect 22930 31614 23044 31666
rect 22876 31612 23044 31614
rect 22876 31602 22932 31612
rect 22652 31500 22820 31556
rect 22540 29922 22596 29932
rect 22652 30324 22708 30334
rect 21980 28814 21982 28866
rect 22034 28814 22036 28866
rect 21308 27132 21476 27188
rect 21532 27636 21588 27646
rect 21084 26964 21140 26974
rect 21084 26740 21140 26908
rect 21084 26674 21140 26684
rect 20972 26126 20974 26178
rect 21026 26126 21028 26178
rect 20972 26114 21028 26126
rect 21196 26290 21252 26302
rect 21196 26238 21198 26290
rect 21250 26238 21252 26290
rect 21196 26068 21252 26238
rect 21196 26002 21252 26012
rect 21308 24836 21364 27132
rect 21308 24770 21364 24780
rect 21420 26964 21476 26974
rect 21420 24162 21476 26908
rect 21532 26962 21588 27580
rect 21532 26910 21534 26962
rect 21586 26910 21588 26962
rect 21532 26898 21588 26910
rect 21644 27076 21700 27086
rect 21644 26962 21700 27020
rect 21644 26910 21646 26962
rect 21698 26910 21700 26962
rect 21644 26898 21700 26910
rect 21756 26962 21812 26974
rect 21756 26910 21758 26962
rect 21810 26910 21812 26962
rect 21756 26908 21812 26910
rect 21868 26962 21924 26974
rect 21868 26910 21870 26962
rect 21922 26910 21924 26962
rect 21868 26908 21924 26910
rect 21756 26852 21924 26908
rect 21868 26740 21924 26750
rect 21756 26290 21812 26302
rect 21756 26238 21758 26290
rect 21810 26238 21812 26290
rect 21644 25508 21700 25518
rect 21644 25414 21700 25452
rect 21420 24110 21422 24162
rect 21474 24110 21476 24162
rect 21420 24098 21476 24110
rect 21756 24052 21812 26238
rect 21756 23986 21812 23996
rect 21868 24050 21924 26684
rect 21980 25284 22036 28814
rect 22092 29260 22260 29316
rect 22428 29876 22484 29886
rect 22428 29426 22484 29820
rect 22428 29374 22430 29426
rect 22482 29374 22484 29426
rect 22092 28644 22148 29260
rect 22428 29092 22484 29374
rect 22428 29026 22484 29036
rect 22092 28578 22148 28588
rect 22540 28644 22596 28654
rect 22316 28308 22372 28318
rect 22092 26964 22148 26974
rect 22204 26964 22260 27002
rect 22092 26962 22260 26964
rect 22092 26910 22094 26962
rect 22146 26910 22206 26962
rect 22258 26910 22260 26962
rect 22092 26908 22260 26910
rect 22092 26898 22148 26908
rect 22092 26516 22148 26526
rect 22092 26422 22148 26460
rect 21980 25218 22036 25228
rect 22204 25172 22260 26908
rect 22316 25396 22372 28252
rect 22316 25302 22372 25340
rect 22428 26068 22484 26078
rect 22092 25116 22260 25172
rect 22092 24388 22148 25116
rect 22428 25060 22484 26012
rect 22092 24162 22148 24332
rect 22092 24110 22094 24162
rect 22146 24110 22148 24162
rect 22092 24098 22148 24110
rect 22204 25004 22484 25060
rect 21868 23998 21870 24050
rect 21922 23998 21924 24050
rect 21308 23940 21364 23950
rect 21308 23846 21364 23884
rect 21756 23828 21812 23838
rect 21420 23714 21476 23726
rect 21420 23662 21422 23714
rect 21474 23662 21476 23714
rect 21420 23604 21476 23662
rect 21420 23538 21476 23548
rect 21756 23492 21812 23772
rect 21868 23716 21924 23998
rect 21868 23650 21924 23660
rect 21980 23940 22036 23950
rect 21756 23436 21924 23492
rect 21196 23044 21252 23054
rect 21084 21474 21140 21486
rect 21084 21422 21086 21474
rect 21138 21422 21140 21474
rect 21084 21028 21140 21422
rect 21084 20962 21140 20972
rect 20748 20914 20916 20916
rect 20748 20862 20750 20914
rect 20802 20862 20916 20914
rect 20748 20860 20916 20862
rect 20748 20850 20804 20860
rect 19964 20804 20020 20814
rect 19964 18674 20020 20748
rect 20860 20804 20916 20860
rect 20860 20738 20916 20748
rect 20532 20412 20796 20422
rect 20588 20356 20636 20412
rect 20692 20356 20740 20412
rect 20532 20346 20796 20356
rect 20188 19908 20244 19918
rect 20188 19814 20244 19852
rect 19964 18622 19966 18674
rect 20018 18622 20020 18674
rect 19964 18610 20020 18622
rect 20188 19012 20244 19022
rect 20748 19012 20804 19022
rect 20076 18452 20132 18462
rect 20076 17890 20132 18396
rect 20188 18450 20244 18956
rect 20188 18398 20190 18450
rect 20242 18398 20244 18450
rect 20188 18004 20244 18398
rect 20412 19010 20804 19012
rect 20412 18958 20750 19010
rect 20802 18958 20804 19010
rect 20412 18956 20804 18958
rect 20412 18450 20468 18956
rect 20748 18946 20804 18956
rect 20532 18844 20796 18854
rect 20588 18788 20636 18844
rect 20692 18788 20740 18844
rect 20532 18778 20796 18788
rect 20412 18398 20414 18450
rect 20466 18398 20468 18450
rect 20300 18340 20356 18350
rect 20300 18246 20356 18284
rect 20188 17938 20244 17948
rect 20076 17838 20078 17890
rect 20130 17838 20132 17890
rect 20076 17826 20132 17838
rect 20300 17666 20356 17678
rect 20300 17614 20302 17666
rect 20354 17614 20356 17666
rect 20300 17556 20356 17614
rect 20300 17490 20356 17500
rect 19516 15362 19572 15372
rect 19628 17276 19908 17332
rect 19964 17444 20020 17454
rect 18956 12238 18958 12290
rect 19010 12238 19012 12290
rect 18956 12226 19012 12238
rect 19068 12348 19460 12404
rect 19516 12964 19572 12974
rect 18844 12126 18846 12178
rect 18898 12126 18900 12178
rect 18844 11956 18900 12126
rect 18844 11890 18900 11900
rect 19068 11396 19124 12348
rect 19404 12180 19460 12190
rect 19516 12180 19572 12908
rect 19404 12178 19572 12180
rect 19404 12126 19406 12178
rect 19458 12126 19572 12178
rect 19404 12124 19572 12126
rect 19404 12114 19460 12124
rect 19292 12068 19348 12078
rect 19180 11620 19236 11630
rect 19180 11526 19236 11564
rect 19292 11618 19348 12012
rect 19292 11566 19294 11618
rect 19346 11566 19348 11618
rect 19292 11554 19348 11566
rect 19516 11956 19572 11966
rect 19516 11618 19572 11900
rect 19516 11566 19518 11618
rect 19570 11566 19572 11618
rect 19516 11554 19572 11566
rect 19068 11340 19236 11396
rect 18732 10780 19124 10836
rect 18508 10500 18564 10510
rect 18564 10444 18788 10500
rect 18508 10406 18564 10444
rect 18284 8642 18340 8652
rect 18284 8372 18340 8382
rect 17500 8370 18340 8372
rect 17500 8318 17502 8370
rect 17554 8318 18286 8370
rect 18338 8318 18340 8370
rect 17500 8316 18340 8318
rect 17500 8306 17556 8316
rect 18284 8306 18340 8316
rect 18732 8148 18788 10444
rect 18844 9044 18900 9054
rect 18844 8950 18900 8988
rect 18956 8708 19012 8718
rect 18844 8148 18900 8158
rect 17388 8092 17892 8148
rect 15932 8036 15988 8046
rect 15932 7586 15988 7980
rect 17500 7700 17556 7710
rect 17500 7606 17556 7644
rect 15932 7534 15934 7586
rect 15986 7534 15988 7586
rect 15932 7522 15988 7534
rect 15820 6018 15876 6076
rect 15820 5966 15822 6018
rect 15874 5966 15876 6018
rect 15820 5954 15876 5966
rect 16044 6804 16100 6814
rect 14588 5908 14644 5918
rect 14588 5814 14644 5852
rect 15036 5794 15092 5806
rect 15036 5742 15038 5794
rect 15090 5742 15092 5794
rect 13916 5142 13972 5180
rect 14028 5180 14476 5236
rect 13692 4722 13748 4732
rect 13132 4398 13134 4450
rect 13186 4398 13188 4450
rect 13132 4386 13188 4398
rect 14028 4338 14084 5180
rect 14476 5170 14532 5180
rect 14700 5460 14756 5470
rect 14700 5122 14756 5404
rect 15036 5460 15092 5742
rect 15036 5394 15092 5404
rect 15148 5684 15204 5694
rect 14700 5070 14702 5122
rect 14754 5070 14756 5122
rect 14700 5058 14756 5070
rect 14476 5010 14532 5022
rect 14476 4958 14478 5010
rect 14530 4958 14532 5010
rect 14476 4788 14532 4958
rect 14476 4722 14532 4732
rect 14700 4452 14756 4462
rect 14700 4358 14756 4396
rect 14028 4286 14030 4338
rect 14082 4286 14084 4338
rect 14028 4274 14084 4286
rect 12236 3948 12628 4004
rect 8204 3378 8260 3388
rect 11340 3332 11508 3388
rect 11676 3444 11732 3482
rect 11900 3444 11956 3454
rect 11676 3442 11956 3444
rect 11676 3390 11678 3442
rect 11730 3390 11902 3442
rect 11954 3390 11956 3442
rect 11676 3388 11956 3390
rect 11340 2996 11396 3332
rect 11340 2930 11396 2940
rect 11676 800 11732 3388
rect 11900 3378 11956 3388
rect 12236 3442 12292 3948
rect 12236 3390 12238 3442
rect 12290 3390 12292 3442
rect 12236 3378 12292 3390
rect 15148 2772 15204 5628
rect 15708 5684 15764 5694
rect 15708 5122 15764 5628
rect 15708 5070 15710 5122
rect 15762 5070 15764 5122
rect 15708 5058 15764 5070
rect 15372 4898 15428 4910
rect 15372 4846 15374 4898
rect 15426 4846 15428 4898
rect 15372 4452 15428 4846
rect 15372 4386 15428 4396
rect 15148 2706 15204 2716
rect 15708 3444 15764 3482
rect 15932 3444 15988 3454
rect 15708 3442 15988 3444
rect 15708 3390 15710 3442
rect 15762 3390 15934 3442
rect 15986 3390 15988 3442
rect 15708 3388 15988 3390
rect 16044 3444 16100 6748
rect 16156 6020 16212 6030
rect 16828 6020 16884 6030
rect 16156 6018 16324 6020
rect 16156 5966 16158 6018
rect 16210 5966 16324 6018
rect 16156 5964 16324 5966
rect 16156 5954 16212 5964
rect 16268 5124 16324 5964
rect 16828 6018 17108 6020
rect 16828 5966 16830 6018
rect 16882 5966 17108 6018
rect 16828 5964 17108 5966
rect 16828 5954 16884 5964
rect 16268 5030 16324 5068
rect 16604 5906 16660 5918
rect 16604 5854 16606 5906
rect 16658 5854 16660 5906
rect 16604 4564 16660 5854
rect 16604 4498 16660 4508
rect 16716 5796 16772 5806
rect 16716 4452 16772 5740
rect 17052 5234 17108 5964
rect 17836 5908 17892 8092
rect 18732 8146 18900 8148
rect 18732 8094 18846 8146
rect 18898 8094 18900 8146
rect 18732 8092 18900 8094
rect 17948 8036 18004 8046
rect 17948 7942 18004 7980
rect 18732 7700 18788 8092
rect 18844 8082 18900 8092
rect 18732 7634 18788 7644
rect 18508 6018 18564 6030
rect 18508 5966 18510 6018
rect 18562 5966 18564 6018
rect 17052 5182 17054 5234
rect 17106 5182 17108 5234
rect 17052 5170 17108 5182
rect 17164 5906 17892 5908
rect 17164 5854 17838 5906
rect 17890 5854 17892 5906
rect 17164 5852 17892 5854
rect 17164 5012 17220 5852
rect 17836 5842 17892 5852
rect 18396 5906 18452 5918
rect 18396 5854 18398 5906
rect 18450 5854 18452 5906
rect 18396 5796 18452 5854
rect 18396 5730 18452 5740
rect 17500 5684 17556 5694
rect 17500 5590 17556 5628
rect 16716 4386 16772 4396
rect 16828 4956 17220 5012
rect 17948 5236 18004 5246
rect 16828 4226 16884 4956
rect 17612 4564 17668 4574
rect 17612 4470 17668 4508
rect 17948 4338 18004 5180
rect 18508 4788 18564 5966
rect 18956 5236 19012 8652
rect 19068 8596 19124 10780
rect 19068 8530 19124 8540
rect 19068 8260 19124 8270
rect 19068 8166 19124 8204
rect 19180 6468 19236 11340
rect 19628 10500 19684 17276
rect 19740 16884 19796 16894
rect 19740 12180 19796 16828
rect 19852 16884 19908 16894
rect 19964 16884 20020 17388
rect 20412 17108 20468 18398
rect 20748 18562 20804 18574
rect 20748 18510 20750 18562
rect 20802 18510 20804 18562
rect 20748 18340 20804 18510
rect 20860 18562 20916 18574
rect 20860 18510 20862 18562
rect 20914 18510 20916 18562
rect 20860 18452 20916 18510
rect 20860 18386 20916 18396
rect 21084 18450 21140 18462
rect 21084 18398 21086 18450
rect 21138 18398 21140 18450
rect 20748 18274 20804 18284
rect 21084 18340 21140 18398
rect 21084 18274 21140 18284
rect 20748 18004 20804 18014
rect 20748 17668 20804 17948
rect 20748 17574 20804 17612
rect 20532 17276 20796 17286
rect 20588 17220 20636 17276
rect 20692 17220 20740 17276
rect 20532 17210 20796 17220
rect 20412 17052 20692 17108
rect 20412 16884 20468 16894
rect 19852 16882 20468 16884
rect 19852 16830 19854 16882
rect 19906 16830 20414 16882
rect 20466 16830 20468 16882
rect 19852 16828 20468 16830
rect 19852 16818 19908 16828
rect 19852 15988 19908 15998
rect 19852 15894 19908 15932
rect 20188 15876 20244 15886
rect 20188 15782 20244 15820
rect 20412 15204 20468 16828
rect 20636 15876 20692 17052
rect 20636 15810 20692 15820
rect 20532 15708 20796 15718
rect 20588 15652 20636 15708
rect 20692 15652 20740 15708
rect 20532 15642 20796 15652
rect 20412 15138 20468 15148
rect 21196 15148 21252 22988
rect 21420 21588 21476 21598
rect 21420 20914 21476 21532
rect 21868 21362 21924 23436
rect 21980 23266 22036 23884
rect 22204 23716 22260 25004
rect 21980 23214 21982 23266
rect 22034 23214 22036 23266
rect 21980 23202 22036 23214
rect 22092 23660 22260 23716
rect 22316 24722 22372 24734
rect 22316 24670 22318 24722
rect 22370 24670 22372 24722
rect 22092 23042 22148 23660
rect 22204 23492 22260 23502
rect 22204 23378 22260 23436
rect 22204 23326 22206 23378
rect 22258 23326 22260 23378
rect 22204 23314 22260 23326
rect 22092 22990 22094 23042
rect 22146 22990 22148 23042
rect 22092 22978 22148 22990
rect 22204 22596 22260 22606
rect 22316 22596 22372 24670
rect 22540 24276 22596 28588
rect 22652 28532 22708 30268
rect 22764 29988 22820 31500
rect 22876 31106 22932 31118
rect 22876 31054 22878 31106
rect 22930 31054 22932 31106
rect 22876 30212 22932 31054
rect 22876 30146 22932 30156
rect 22764 29932 22932 29988
rect 22764 29650 22820 29662
rect 22764 29598 22766 29650
rect 22818 29598 22820 29650
rect 22764 28644 22820 29598
rect 22876 29316 22932 29932
rect 22988 29428 23044 31612
rect 23548 31556 23604 31726
rect 23660 31780 23716 32398
rect 23660 31714 23716 31724
rect 23884 32338 23940 32350
rect 23884 32286 23886 32338
rect 23938 32286 23940 32338
rect 23884 31780 23940 32286
rect 23884 31714 23940 31724
rect 23548 30996 23604 31500
rect 23548 30930 23604 30940
rect 23884 31554 23940 31566
rect 23884 31502 23886 31554
rect 23938 31502 23940 31554
rect 23884 30996 23940 31502
rect 23884 30930 23940 30940
rect 23436 30882 23492 30894
rect 23436 30830 23438 30882
rect 23490 30830 23492 30882
rect 23324 30436 23380 30446
rect 23324 30322 23380 30380
rect 23324 30270 23326 30322
rect 23378 30270 23380 30322
rect 23324 30258 23380 30270
rect 23436 29652 23492 30830
rect 23772 30212 23828 30222
rect 23436 29586 23492 29596
rect 23548 30210 23828 30212
rect 23548 30158 23774 30210
rect 23826 30158 23828 30210
rect 23548 30156 23828 30158
rect 23436 29428 23492 29438
rect 22988 29426 23492 29428
rect 22988 29374 23438 29426
rect 23490 29374 23492 29426
rect 22988 29372 23492 29374
rect 23436 29362 23492 29372
rect 22876 29260 23044 29316
rect 22764 28578 22820 28588
rect 22876 28980 22932 28990
rect 22652 28466 22708 28476
rect 22876 28308 22932 28924
rect 22876 28242 22932 28252
rect 22876 27972 22932 27982
rect 22876 27878 22932 27916
rect 22988 27748 23044 29260
rect 23100 28868 23156 28878
rect 23100 28420 23156 28812
rect 23100 27970 23156 28364
rect 23100 27918 23102 27970
rect 23154 27918 23156 27970
rect 23100 27906 23156 27918
rect 23212 28756 23268 28766
rect 23212 27860 23268 28700
rect 23548 28532 23604 30156
rect 23772 30146 23828 30156
rect 23996 30212 24052 32620
rect 24220 31778 24276 31790
rect 24220 31726 24222 31778
rect 24274 31726 24276 31778
rect 24220 31556 24276 31726
rect 24220 31490 24276 31500
rect 24108 31106 24164 31118
rect 24108 31054 24110 31106
rect 24162 31054 24164 31106
rect 24108 30436 24164 31054
rect 24108 30370 24164 30380
rect 24444 30212 24500 34190
rect 23996 30118 24052 30156
rect 24108 30156 24500 30212
rect 23324 28476 23604 28532
rect 23660 29876 23716 29886
rect 23324 28082 23380 28476
rect 23324 28030 23326 28082
rect 23378 28030 23380 28082
rect 23324 28018 23380 28030
rect 23436 27860 23492 27870
rect 23212 27858 23492 27860
rect 23212 27806 23438 27858
rect 23490 27806 23492 27858
rect 23212 27804 23492 27806
rect 23436 27794 23492 27804
rect 22988 27692 23156 27748
rect 22652 26964 22708 27002
rect 22652 26898 22708 26908
rect 23100 26908 23156 27692
rect 23548 27076 23604 27086
rect 22764 26852 22820 26862
rect 22764 26850 22932 26852
rect 22764 26798 22766 26850
rect 22818 26798 22932 26850
rect 22764 26796 22932 26798
rect 22764 26786 22820 26796
rect 22652 26178 22708 26190
rect 22652 26126 22654 26178
rect 22706 26126 22708 26178
rect 22652 25508 22708 26126
rect 22652 25442 22708 25452
rect 22540 24210 22596 24220
rect 22764 23826 22820 23838
rect 22764 23774 22766 23826
rect 22818 23774 22820 23826
rect 22428 23716 22484 23726
rect 22764 23716 22820 23774
rect 22428 23714 22820 23716
rect 22428 23662 22430 23714
rect 22482 23662 22820 23714
rect 22428 23660 22820 23662
rect 22428 23378 22484 23660
rect 22428 23326 22430 23378
rect 22482 23326 22484 23378
rect 22428 23314 22484 23326
rect 22764 23266 22820 23660
rect 22876 23378 22932 26796
rect 22988 26850 23044 26862
rect 23100 26852 23380 26908
rect 22988 26798 22990 26850
rect 23042 26798 23044 26850
rect 22988 25508 23044 26798
rect 22988 25442 23044 25452
rect 23100 24052 23156 24062
rect 23324 24052 23380 26852
rect 23548 25506 23604 27020
rect 23660 26514 23716 29820
rect 23884 28644 23940 28654
rect 23660 26462 23662 26514
rect 23714 26462 23716 26514
rect 23660 26450 23716 26462
rect 23772 28420 23828 28430
rect 23548 25454 23550 25506
rect 23602 25454 23604 25506
rect 23548 25442 23604 25454
rect 23548 24724 23604 24762
rect 23548 24658 23604 24668
rect 22988 23828 23044 23838
rect 22988 23604 23044 23772
rect 23100 23714 23156 23996
rect 23100 23662 23102 23714
rect 23154 23662 23156 23714
rect 23100 23650 23156 23662
rect 23212 23996 23380 24052
rect 23436 24500 23492 24510
rect 22988 23538 23044 23548
rect 22876 23326 22878 23378
rect 22930 23326 22932 23378
rect 22876 23314 22932 23326
rect 23212 23268 23268 23996
rect 23436 23940 23492 24444
rect 23772 23940 23828 28364
rect 23884 24610 23940 28588
rect 23884 24558 23886 24610
rect 23938 24558 23940 24610
rect 23884 24546 23940 24558
rect 23996 27748 24052 27758
rect 23436 23846 23492 23884
rect 23660 23884 23828 23940
rect 23884 24388 23940 24398
rect 22764 23214 22766 23266
rect 22818 23214 22820 23266
rect 22764 23202 22820 23214
rect 22988 23212 23268 23268
rect 23324 23828 23380 23838
rect 22204 22594 22372 22596
rect 22204 22542 22206 22594
rect 22258 22542 22372 22594
rect 22204 22540 22372 22542
rect 22204 22530 22260 22540
rect 22092 22372 22148 22382
rect 22092 22278 22148 22316
rect 21868 21310 21870 21362
rect 21922 21310 21924 21362
rect 21868 21298 21924 21310
rect 21980 22148 22036 22158
rect 21420 20862 21422 20914
rect 21474 20862 21476 20914
rect 21420 20850 21476 20862
rect 21308 20802 21364 20814
rect 21308 20750 21310 20802
rect 21362 20750 21364 20802
rect 21308 20692 21364 20750
rect 21308 20626 21364 20636
rect 21532 20804 21588 20814
rect 21532 18788 21588 20748
rect 21868 20802 21924 20814
rect 21868 20750 21870 20802
rect 21922 20750 21924 20802
rect 21756 20692 21812 20702
rect 21756 20598 21812 20636
rect 21868 19908 21924 20750
rect 21868 19842 21924 19852
rect 21980 19684 22036 22092
rect 22204 22148 22260 22158
rect 22876 22148 22932 22158
rect 22204 22146 22932 22148
rect 22204 22094 22206 22146
rect 22258 22094 22878 22146
rect 22930 22094 22932 22146
rect 22204 22092 22932 22094
rect 22204 22082 22260 22092
rect 22092 21474 22148 21486
rect 22428 21476 22484 21486
rect 22092 21422 22094 21474
rect 22146 21422 22148 21474
rect 22092 20692 22148 21422
rect 22092 20626 22148 20636
rect 22316 21420 22428 21476
rect 21980 19618 22036 19628
rect 22204 20578 22260 20590
rect 22204 20526 22206 20578
rect 22258 20526 22260 20578
rect 21868 19572 21924 19582
rect 21756 19348 21812 19358
rect 21868 19348 21924 19516
rect 21756 19346 21924 19348
rect 21756 19294 21758 19346
rect 21810 19294 21924 19346
rect 21756 19292 21924 19294
rect 21756 19282 21812 19292
rect 22204 19234 22260 20526
rect 22316 20356 22372 21420
rect 22428 21382 22484 21420
rect 22540 21362 22596 21374
rect 22540 21310 22542 21362
rect 22594 21310 22596 21362
rect 22540 21252 22596 21310
rect 22428 21196 22596 21252
rect 22428 20690 22484 21196
rect 22428 20638 22430 20690
rect 22482 20638 22484 20690
rect 22428 20626 22484 20638
rect 22540 20690 22596 20702
rect 22540 20638 22542 20690
rect 22594 20638 22596 20690
rect 22540 20356 22596 20638
rect 22316 20300 22484 20356
rect 22316 19906 22372 19918
rect 22316 19854 22318 19906
rect 22370 19854 22372 19906
rect 22316 19572 22372 19854
rect 22316 19506 22372 19516
rect 22204 19182 22206 19234
rect 22258 19182 22260 19234
rect 22204 19170 22260 19182
rect 22316 19346 22372 19358
rect 22316 19294 22318 19346
rect 22370 19294 22372 19346
rect 21644 19124 21700 19134
rect 21644 19030 21700 19068
rect 21980 19124 22036 19134
rect 21868 19012 21924 19022
rect 21868 18918 21924 18956
rect 21980 18900 22036 19068
rect 21532 18732 21924 18788
rect 21420 18450 21476 18462
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 21420 17556 21476 18398
rect 21532 17778 21588 18732
rect 21868 18674 21924 18732
rect 21868 18622 21870 18674
rect 21922 18622 21924 18674
rect 21868 18610 21924 18622
rect 21756 18564 21812 18574
rect 21532 17726 21534 17778
rect 21586 17726 21588 17778
rect 21532 17714 21588 17726
rect 21644 18450 21700 18462
rect 21644 18398 21646 18450
rect 21698 18398 21700 18450
rect 21644 17668 21700 18398
rect 21644 17602 21700 17612
rect 21420 17490 21476 17500
rect 21532 15540 21588 15550
rect 21532 15314 21588 15484
rect 21532 15262 21534 15314
rect 21586 15262 21588 15314
rect 21196 15092 21476 15148
rect 20860 14980 20916 14990
rect 20188 14308 20244 14318
rect 20076 14084 20132 14094
rect 20076 13074 20132 14028
rect 20076 13022 20078 13074
rect 20130 13022 20132 13074
rect 20076 12852 20132 13022
rect 19964 12740 20020 12750
rect 19852 12180 19908 12190
rect 19740 12178 19908 12180
rect 19740 12126 19854 12178
rect 19906 12126 19908 12178
rect 19740 12124 19908 12126
rect 19740 11732 19796 12124
rect 19852 12114 19908 12124
rect 19964 11732 20020 12684
rect 20076 12180 20132 12796
rect 20076 12114 20132 12124
rect 20188 13636 20244 14252
rect 20532 14140 20796 14150
rect 20588 14084 20636 14140
rect 20692 14084 20740 14140
rect 20532 14074 20796 14084
rect 20860 13860 20916 14924
rect 21308 14308 21364 14318
rect 21308 14214 21364 14252
rect 20076 11956 20132 11966
rect 20076 11862 20132 11900
rect 19964 11676 20132 11732
rect 19740 11666 19796 11676
rect 19964 11172 20020 11182
rect 19628 10434 19684 10444
rect 19740 11170 20020 11172
rect 19740 11118 19966 11170
rect 20018 11118 20020 11170
rect 19740 11116 20020 11118
rect 19740 9940 19796 11116
rect 19964 11106 20020 11116
rect 19852 10724 19908 10734
rect 19852 10500 19908 10668
rect 19964 10724 20020 10734
rect 20076 10724 20132 11676
rect 20188 10834 20244 13580
rect 20524 13636 20580 13646
rect 20412 13074 20468 13086
rect 20412 13022 20414 13074
rect 20466 13022 20468 13074
rect 20300 12852 20356 12862
rect 20300 12758 20356 12796
rect 20412 12404 20468 13022
rect 20524 12962 20580 13580
rect 20524 12910 20526 12962
rect 20578 12910 20580 12962
rect 20524 12898 20580 12910
rect 20860 12962 20916 13804
rect 20860 12910 20862 12962
rect 20914 12910 20916 12962
rect 20860 12898 20916 12910
rect 21084 13634 21140 13646
rect 21084 13582 21086 13634
rect 21138 13582 21140 13634
rect 21084 12964 21140 13582
rect 21084 12908 21364 12964
rect 21196 12740 21252 12750
rect 21084 12738 21252 12740
rect 21084 12686 21198 12738
rect 21250 12686 21252 12738
rect 21084 12684 21252 12686
rect 20532 12572 20796 12582
rect 20588 12516 20636 12572
rect 20692 12516 20740 12572
rect 20532 12506 20796 12516
rect 20412 12348 20692 12404
rect 20636 12290 20692 12348
rect 20972 12292 21028 12302
rect 20636 12238 20638 12290
rect 20690 12238 20692 12290
rect 20636 12226 20692 12238
rect 20748 12290 21028 12292
rect 20748 12238 20974 12290
rect 21026 12238 21028 12290
rect 20748 12236 21028 12238
rect 20412 12180 20468 12190
rect 20188 10782 20190 10834
rect 20242 10782 20244 10834
rect 20188 10770 20244 10782
rect 20300 12178 20468 12180
rect 20300 12126 20414 12178
rect 20466 12126 20468 12178
rect 20300 12124 20468 12126
rect 19964 10722 20132 10724
rect 19964 10670 19966 10722
rect 20018 10670 20132 10722
rect 19964 10668 20132 10670
rect 19964 10658 20020 10668
rect 19852 10434 19908 10444
rect 20300 10052 20356 12124
rect 20412 12114 20468 12124
rect 20524 11956 20580 11966
rect 20748 11956 20804 12236
rect 20524 11954 20804 11956
rect 20524 11902 20526 11954
rect 20578 11902 20804 11954
rect 20524 11900 20804 11902
rect 20860 11956 20916 11966
rect 20524 11890 20580 11900
rect 20860 11396 20916 11900
rect 20972 11732 21028 12236
rect 20972 11666 21028 11676
rect 20860 11330 20916 11340
rect 20412 11284 20468 11294
rect 21084 11284 21140 12684
rect 21196 12674 21252 12684
rect 21308 12738 21364 12908
rect 21308 12686 21310 12738
rect 21362 12686 21364 12738
rect 21308 12292 21364 12686
rect 20412 10722 20468 11228
rect 20972 11228 21140 11284
rect 21196 12236 21364 12292
rect 20532 11004 20796 11014
rect 20588 10948 20636 11004
rect 20692 10948 20740 11004
rect 20532 10938 20796 10948
rect 20972 10834 21028 11228
rect 21196 11060 21252 12236
rect 21308 12066 21364 12078
rect 21308 12014 21310 12066
rect 21362 12014 21364 12066
rect 21308 11788 21364 12014
rect 21420 11956 21476 15092
rect 21532 14530 21588 15262
rect 21532 14478 21534 14530
rect 21586 14478 21588 14530
rect 21532 14466 21588 14478
rect 21756 15538 21812 18508
rect 21980 18452 22036 18844
rect 21756 15486 21758 15538
rect 21810 15486 21812 15538
rect 21532 13748 21588 13758
rect 21532 13076 21588 13692
rect 21756 13636 21812 15486
rect 21868 18396 22036 18452
rect 21868 14196 21924 18396
rect 21980 18228 22036 18238
rect 21980 18134 22036 18172
rect 22092 17668 22148 17678
rect 22092 17442 22148 17612
rect 22092 17390 22094 17442
rect 22146 17390 22148 17442
rect 22092 16548 22148 17390
rect 22316 17332 22372 19294
rect 22316 17266 22372 17276
rect 22092 16482 22148 16492
rect 22092 16212 22148 16222
rect 22092 16118 22148 16156
rect 22204 15540 22260 15550
rect 22092 14644 22148 14654
rect 22204 14644 22260 15484
rect 22428 15148 22484 20300
rect 22540 20290 22596 20300
rect 22652 19346 22708 22092
rect 22876 22082 22932 22092
rect 22652 19294 22654 19346
rect 22706 19294 22708 19346
rect 22652 19282 22708 19294
rect 22764 21924 22820 21934
rect 22540 18562 22596 18574
rect 22540 18510 22542 18562
rect 22594 18510 22596 18562
rect 22540 18452 22596 18510
rect 22540 18386 22596 18396
rect 22652 18340 22708 18350
rect 22540 18228 22596 18238
rect 22540 17890 22596 18172
rect 22652 18226 22708 18284
rect 22652 18174 22654 18226
rect 22706 18174 22708 18226
rect 22652 18162 22708 18174
rect 22540 17838 22542 17890
rect 22594 17838 22596 17890
rect 22540 17826 22596 17838
rect 22764 17780 22820 21868
rect 22988 21812 23044 23212
rect 22988 21718 23044 21756
rect 22988 21362 23044 21374
rect 22988 21310 22990 21362
rect 23042 21310 23044 21362
rect 22988 20914 23044 21310
rect 22988 20862 22990 20914
rect 23042 20862 23044 20914
rect 22988 20850 23044 20862
rect 23100 20020 23156 20030
rect 23100 19926 23156 19964
rect 23324 19796 23380 23772
rect 23436 23716 23492 23726
rect 23436 23378 23492 23660
rect 23436 23326 23438 23378
rect 23490 23326 23492 23378
rect 23436 23314 23492 23326
rect 23548 22146 23604 22158
rect 23548 22094 23550 22146
rect 23602 22094 23604 22146
rect 23548 22036 23604 22094
rect 23548 21970 23604 21980
rect 23436 21588 23492 21598
rect 23436 21494 23492 21532
rect 23548 20578 23604 20590
rect 23548 20526 23550 20578
rect 23602 20526 23604 20578
rect 23548 20356 23604 20526
rect 23548 20290 23604 20300
rect 23548 19908 23604 19918
rect 23548 19814 23604 19852
rect 23324 19730 23380 19740
rect 23436 19794 23492 19806
rect 23436 19742 23438 19794
rect 23490 19742 23492 19794
rect 23100 19460 23156 19470
rect 22092 14642 22260 14644
rect 22092 14590 22094 14642
rect 22146 14590 22260 14642
rect 22092 14588 22260 14590
rect 22316 15092 22484 15148
rect 22652 17724 22820 17780
rect 22876 19234 22932 19246
rect 22876 19182 22878 19234
rect 22930 19182 22932 19234
rect 22876 18452 22932 19182
rect 22876 17778 22932 18396
rect 22876 17726 22878 17778
rect 22930 17726 22932 17778
rect 22092 14578 22148 14588
rect 21868 14130 21924 14140
rect 21756 13570 21812 13580
rect 22092 14084 22148 14094
rect 21980 13524 22036 13534
rect 21532 12962 21588 13020
rect 21532 12910 21534 12962
rect 21586 12910 21588 12962
rect 21532 12898 21588 12910
rect 21756 13076 21812 13086
rect 21756 12850 21812 13020
rect 21756 12798 21758 12850
rect 21810 12798 21812 12850
rect 21756 12740 21812 12798
rect 21756 12674 21812 12684
rect 21756 12068 21812 12078
rect 21420 11900 21700 11956
rect 21308 11732 21588 11788
rect 21308 11508 21364 11518
rect 21308 11414 21364 11452
rect 20972 10782 20974 10834
rect 21026 10782 21028 10834
rect 20972 10770 21028 10782
rect 21084 11004 21252 11060
rect 21532 11394 21588 11732
rect 21532 11342 21534 11394
rect 21586 11342 21588 11394
rect 20412 10670 20414 10722
rect 20466 10670 20468 10722
rect 20412 10388 20468 10670
rect 20524 10612 20580 10622
rect 20860 10612 20916 10622
rect 20524 10610 20916 10612
rect 20524 10558 20526 10610
rect 20578 10558 20862 10610
rect 20914 10558 20916 10610
rect 20524 10556 20916 10558
rect 20524 10546 20580 10556
rect 20860 10546 20916 10556
rect 20412 10332 20580 10388
rect 19740 9874 19796 9884
rect 19852 9996 20300 10052
rect 19852 9826 19908 9996
rect 20300 9958 20356 9996
rect 19852 9774 19854 9826
rect 19906 9774 19908 9826
rect 19852 9762 19908 9774
rect 20188 9828 20244 9838
rect 20412 9828 20468 9838
rect 20188 9826 20468 9828
rect 20188 9774 20190 9826
rect 20242 9774 20414 9826
rect 20466 9774 20468 9826
rect 20188 9772 20468 9774
rect 20188 9762 20244 9772
rect 20412 9762 20468 9772
rect 19292 9716 19348 9726
rect 19628 9716 19684 9726
rect 19292 9714 19628 9716
rect 19292 9662 19294 9714
rect 19346 9662 19628 9714
rect 19292 9660 19628 9662
rect 19292 9650 19348 9660
rect 19628 9622 19684 9660
rect 19740 9602 19796 9614
rect 20524 9604 20580 10332
rect 21084 10164 21140 11004
rect 21196 10836 21252 10846
rect 21420 10836 21476 10846
rect 21196 10834 21420 10836
rect 21196 10782 21198 10834
rect 21250 10782 21420 10834
rect 21196 10780 21420 10782
rect 21196 10770 21252 10780
rect 21420 10770 21476 10780
rect 21532 10388 21588 11342
rect 21532 10322 21588 10332
rect 21196 10164 21252 10174
rect 21084 10108 21196 10164
rect 21196 10098 21252 10108
rect 21308 10052 21364 10062
rect 21532 10052 21588 10062
rect 21308 9958 21364 9996
rect 21420 9996 21532 10052
rect 20748 9940 20804 9950
rect 20748 9826 20804 9884
rect 21420 9938 21476 9996
rect 21420 9886 21422 9938
rect 21474 9886 21476 9938
rect 21420 9874 21476 9886
rect 20748 9774 20750 9826
rect 20802 9774 20804 9826
rect 20748 9762 20804 9774
rect 19740 9550 19742 9602
rect 19794 9550 19796 9602
rect 19516 9156 19572 9166
rect 19740 9156 19796 9550
rect 20412 9548 20580 9604
rect 20636 9604 20692 9642
rect 19516 9154 19796 9156
rect 19516 9102 19518 9154
rect 19570 9102 19796 9154
rect 19516 9100 19796 9102
rect 19852 9492 19908 9502
rect 19516 9090 19572 9100
rect 19628 8596 19684 8606
rect 19516 8260 19572 8270
rect 19516 7698 19572 8204
rect 19516 7646 19518 7698
rect 19570 7646 19572 7698
rect 19516 7588 19572 7646
rect 19516 7522 19572 7532
rect 19180 6402 19236 6412
rect 19292 5796 19348 5806
rect 19292 5702 19348 5740
rect 19180 5236 19236 5246
rect 19012 5234 19236 5236
rect 19012 5182 19182 5234
rect 19234 5182 19236 5234
rect 19012 5180 19236 5182
rect 18956 5142 19012 5180
rect 19180 5170 19236 5180
rect 18508 4450 18564 4732
rect 18508 4398 18510 4450
rect 18562 4398 18564 4450
rect 18508 4386 18564 4398
rect 17948 4286 17950 4338
rect 18002 4286 18004 4338
rect 17948 4274 18004 4286
rect 18732 4340 18788 4350
rect 18732 4246 18788 4284
rect 19404 4340 19460 4350
rect 19404 4246 19460 4284
rect 16828 4174 16830 4226
rect 16882 4174 16884 4226
rect 16828 4162 16884 4174
rect 16268 3444 16324 3454
rect 16044 3442 16324 3444
rect 16044 3390 16270 3442
rect 16322 3390 16324 3442
rect 16044 3388 16324 3390
rect 15708 800 15764 3388
rect 15932 3378 15988 3388
rect 16268 3378 16324 3388
rect 19628 3332 19684 8540
rect 19852 8370 19908 9436
rect 19852 8318 19854 8370
rect 19906 8318 19908 8370
rect 19852 8306 19908 8318
rect 19964 9044 20020 9054
rect 19740 6580 19796 6590
rect 19964 6580 20020 8988
rect 20412 8820 20468 9548
rect 20636 9538 20692 9548
rect 20532 9436 20796 9446
rect 20588 9380 20636 9436
rect 20692 9380 20740 9436
rect 20532 9370 20796 9380
rect 20412 8754 20468 8764
rect 20748 9156 20804 9166
rect 20748 8372 20804 9100
rect 21532 8932 21588 9996
rect 21644 9156 21700 11900
rect 21756 11618 21812 12012
rect 21756 11566 21758 11618
rect 21810 11566 21812 11618
rect 21756 10836 21812 11566
rect 21756 10770 21812 10780
rect 21756 10498 21812 10510
rect 21756 10446 21758 10498
rect 21810 10446 21812 10498
rect 21756 10164 21812 10446
rect 21756 10098 21812 10108
rect 21868 9940 21924 9950
rect 21980 9940 22036 13468
rect 21924 9884 22036 9940
rect 21868 9846 21924 9884
rect 22092 9716 22148 14028
rect 22204 12068 22260 12078
rect 22204 11974 22260 12012
rect 22204 11620 22260 11630
rect 22204 11506 22260 11564
rect 22204 11454 22206 11506
rect 22258 11454 22260 11506
rect 22204 11442 22260 11454
rect 22316 11172 22372 15092
rect 22652 14980 22708 17724
rect 22876 17714 22932 17726
rect 22988 19012 23044 19022
rect 22764 17556 22820 17566
rect 22988 17556 23044 18956
rect 23100 18788 23156 19404
rect 23100 18722 23156 18732
rect 23324 19234 23380 19246
rect 23324 19182 23326 19234
rect 23378 19182 23380 19234
rect 23324 18340 23380 19182
rect 23436 19012 23492 19742
rect 23436 18946 23492 18956
rect 23436 18788 23492 18798
rect 23436 18450 23492 18732
rect 23436 18398 23438 18450
rect 23490 18398 23492 18450
rect 23436 18386 23492 18398
rect 23660 18452 23716 23884
rect 23772 23716 23828 23726
rect 23884 23716 23940 24332
rect 23772 23714 23940 23716
rect 23772 23662 23774 23714
rect 23826 23662 23940 23714
rect 23772 23660 23940 23662
rect 23772 23604 23828 23660
rect 23772 23538 23828 23548
rect 23996 22596 24052 27692
rect 24108 25618 24164 30156
rect 24220 29538 24276 29550
rect 24220 29486 24222 29538
rect 24274 29486 24276 29538
rect 24220 29316 24276 29486
rect 24220 29250 24276 29260
rect 24556 28644 24612 34524
rect 24780 33460 24836 33470
rect 24780 33366 24836 33404
rect 25116 32900 25172 36430
rect 26236 36484 26292 39200
rect 28700 37268 28756 39200
rect 31164 37268 31220 39200
rect 33628 37268 33684 39200
rect 34972 37268 35028 37278
rect 28700 37212 29204 37268
rect 31164 37212 31668 37268
rect 33628 37212 33908 37268
rect 26236 36418 26292 36428
rect 26348 37044 26404 37054
rect 26348 36594 26404 36988
rect 26348 36542 26350 36594
rect 26402 36542 26404 36594
rect 25340 36260 25396 36270
rect 25340 35698 25396 36204
rect 25900 36258 25956 36270
rect 25900 36206 25902 36258
rect 25954 36206 25956 36258
rect 25900 35812 25956 36206
rect 25900 35746 25956 35756
rect 25340 35646 25342 35698
rect 25394 35646 25396 35698
rect 25340 35140 25396 35646
rect 26348 35700 26404 36542
rect 29148 36596 29204 37212
rect 27356 36484 27412 36494
rect 27356 36390 27412 36428
rect 28252 36484 28308 36494
rect 27020 36372 27076 36382
rect 27020 36278 27076 36316
rect 26684 36260 26740 36270
rect 27692 36260 27748 36270
rect 26348 35634 26404 35644
rect 26572 36258 26740 36260
rect 26572 36206 26686 36258
rect 26738 36206 26740 36258
rect 26572 36204 26740 36206
rect 26012 35588 26068 35598
rect 25340 35074 25396 35084
rect 25452 35586 26068 35588
rect 25452 35534 26014 35586
rect 26066 35534 26068 35586
rect 25452 35532 26068 35534
rect 25452 35138 25508 35532
rect 26012 35522 26068 35532
rect 25452 35086 25454 35138
rect 25506 35086 25508 35138
rect 25452 35074 25508 35086
rect 26572 35140 26628 36204
rect 26684 36194 26740 36204
rect 27580 36258 27748 36260
rect 27580 36206 27694 36258
rect 27746 36206 27748 36258
rect 27580 36204 27748 36206
rect 26572 34916 26628 35084
rect 27356 35140 27412 35150
rect 26572 34914 26740 34916
rect 26572 34862 26574 34914
rect 26626 34862 26740 34914
rect 26572 34860 26740 34862
rect 26572 34850 26628 34860
rect 25340 34804 25396 34814
rect 25900 34804 25956 34814
rect 25340 34802 25508 34804
rect 25340 34750 25342 34802
rect 25394 34750 25508 34802
rect 25340 34748 25508 34750
rect 25340 34738 25396 34748
rect 25340 34020 25396 34030
rect 25340 33926 25396 33964
rect 25452 33458 25508 34748
rect 25788 34802 25956 34804
rect 25788 34750 25902 34802
rect 25954 34750 25956 34802
rect 25788 34748 25956 34750
rect 25452 33406 25454 33458
rect 25506 33406 25508 33458
rect 25452 33394 25508 33406
rect 25564 34020 25620 34030
rect 25340 33346 25396 33358
rect 25340 33294 25342 33346
rect 25394 33294 25396 33346
rect 25228 33234 25284 33246
rect 25228 33182 25230 33234
rect 25282 33182 25284 33234
rect 25228 33124 25284 33182
rect 25228 33058 25284 33068
rect 25116 32834 25172 32844
rect 25228 32674 25284 32686
rect 25228 32622 25230 32674
rect 25282 32622 25284 32674
rect 25228 32452 25284 32622
rect 25228 32386 25284 32396
rect 25340 32450 25396 33294
rect 25564 33348 25620 33964
rect 25564 33234 25620 33292
rect 25564 33182 25566 33234
rect 25618 33182 25620 33234
rect 25564 33170 25620 33182
rect 25788 33124 25844 34748
rect 25900 34738 25956 34748
rect 26348 34356 26404 34366
rect 26684 34356 26740 34860
rect 26348 34354 26740 34356
rect 26348 34302 26350 34354
rect 26402 34302 26740 34354
rect 26348 34300 26740 34302
rect 26796 34914 26852 34926
rect 26796 34862 26798 34914
rect 26850 34862 26852 34914
rect 26796 34356 26852 34862
rect 27356 34802 27412 35084
rect 27356 34750 27358 34802
rect 27410 34750 27412 34802
rect 27356 34738 27412 34750
rect 27468 34802 27524 34814
rect 27468 34750 27470 34802
rect 27522 34750 27524 34802
rect 27132 34692 27188 34702
rect 27132 34598 27188 34636
rect 27468 34580 27524 34750
rect 27244 34524 27468 34580
rect 27132 34356 27188 34366
rect 27244 34356 27300 34524
rect 27468 34514 27524 34524
rect 26796 34354 27300 34356
rect 26796 34302 27134 34354
rect 27186 34302 27300 34354
rect 26796 34300 27300 34302
rect 26348 34290 26404 34300
rect 25900 34132 25956 34142
rect 26684 34132 26740 34300
rect 27132 34290 27188 34300
rect 26796 34132 26852 34142
rect 26684 34130 26852 34132
rect 26684 34078 26798 34130
rect 26850 34078 26852 34130
rect 26684 34076 26852 34078
rect 25900 34038 25956 34076
rect 26796 34066 26852 34076
rect 27244 33458 27300 34300
rect 27244 33406 27246 33458
rect 27298 33406 27300 33458
rect 27244 33394 27300 33406
rect 26684 33348 26740 33358
rect 25676 33122 25844 33124
rect 25676 33070 25790 33122
rect 25842 33070 25844 33122
rect 25676 33068 25844 33070
rect 25452 32564 25508 32574
rect 25452 32470 25508 32508
rect 25340 32398 25342 32450
rect 25394 32398 25396 32450
rect 25340 32386 25396 32398
rect 25452 32004 25508 32014
rect 24668 31892 24724 31902
rect 25452 31892 25508 31948
rect 24668 31778 24724 31836
rect 25228 31890 25508 31892
rect 25228 31838 25454 31890
rect 25506 31838 25508 31890
rect 25228 31836 25508 31838
rect 24668 31726 24670 31778
rect 24722 31726 24724 31778
rect 24668 30994 24724 31726
rect 25004 31780 25060 31790
rect 25004 31666 25060 31724
rect 25004 31614 25006 31666
rect 25058 31614 25060 31666
rect 25004 31108 25060 31614
rect 25004 31042 25060 31052
rect 25228 30996 25284 31836
rect 25452 31826 25508 31836
rect 25676 31332 25732 33068
rect 25788 33058 25844 33068
rect 26348 33124 26404 33134
rect 26348 32676 26404 33068
rect 26684 32788 26740 33292
rect 26684 32722 26740 32732
rect 27468 32900 27524 32910
rect 26348 32610 26404 32620
rect 25788 32564 25844 32574
rect 26124 32564 26180 32574
rect 25788 32562 25956 32564
rect 25788 32510 25790 32562
rect 25842 32510 25956 32562
rect 25788 32508 25956 32510
rect 25788 32498 25844 32508
rect 24668 30942 24670 30994
rect 24722 30942 24724 30994
rect 24668 30884 24724 30942
rect 24668 30818 24724 30828
rect 25116 30940 25284 30996
rect 25452 31276 25732 31332
rect 24892 30324 24948 30334
rect 24892 30230 24948 30268
rect 24780 30210 24836 30222
rect 24780 30158 24782 30210
rect 24834 30158 24836 30210
rect 24668 28868 24724 28878
rect 24780 28868 24836 30158
rect 25116 29876 25172 30940
rect 25340 30884 25396 30894
rect 25116 29810 25172 29820
rect 25228 30882 25396 30884
rect 25228 30830 25342 30882
rect 25394 30830 25396 30882
rect 25228 30828 25396 30830
rect 25228 29540 25284 30828
rect 25340 30818 25396 30828
rect 25452 30660 25508 31276
rect 25900 30994 25956 32508
rect 26124 32470 26180 32508
rect 27356 32564 27412 32574
rect 27356 32470 27412 32508
rect 26572 32452 26628 32462
rect 26236 31780 26292 31790
rect 25900 30942 25902 30994
rect 25954 30942 25956 30994
rect 25116 29484 25284 29540
rect 25340 30604 25508 30660
rect 25564 30884 25620 30894
rect 25116 29204 25172 29484
rect 24668 28866 24836 28868
rect 24668 28814 24670 28866
rect 24722 28814 24836 28866
rect 24668 28812 24836 28814
rect 25004 29148 25172 29204
rect 25228 29316 25284 29326
rect 24668 28802 24724 28812
rect 24892 28756 24948 28766
rect 24556 28588 24724 28644
rect 24332 28418 24388 28430
rect 24332 28366 24334 28418
rect 24386 28366 24388 28418
rect 24332 27972 24388 28366
rect 24556 28420 24612 28430
rect 24668 28420 24724 28588
rect 24892 28642 24948 28700
rect 24892 28590 24894 28642
rect 24946 28590 24948 28642
rect 24892 28578 24948 28590
rect 24668 28364 24948 28420
rect 24556 28326 24612 28364
rect 24556 28084 24612 28094
rect 24556 27990 24612 28028
rect 24332 27906 24388 27916
rect 24444 27970 24500 27982
rect 24444 27918 24446 27970
rect 24498 27918 24500 27970
rect 24444 27524 24500 27918
rect 24444 27458 24500 27468
rect 24668 27634 24724 27646
rect 24668 27582 24670 27634
rect 24722 27582 24724 27634
rect 24668 27300 24724 27582
rect 24780 27300 24836 27310
rect 24668 27298 24836 27300
rect 24668 27246 24782 27298
rect 24834 27246 24836 27298
rect 24668 27244 24836 27246
rect 24556 26964 24612 27002
rect 24556 26898 24612 26908
rect 24332 26292 24388 26302
rect 24108 25566 24110 25618
rect 24162 25566 24164 25618
rect 24108 23828 24164 25566
rect 24220 26290 24388 26292
rect 24220 26238 24334 26290
rect 24386 26238 24388 26290
rect 24220 26236 24388 26238
rect 24220 25620 24276 26236
rect 24332 26226 24388 26236
rect 24220 25506 24276 25564
rect 24220 25454 24222 25506
rect 24274 25454 24276 25506
rect 24220 25442 24276 25454
rect 24444 24724 24500 24734
rect 24500 24668 24612 24724
rect 24444 24658 24500 24668
rect 24108 23772 24500 23828
rect 23884 22540 24052 22596
rect 24108 23042 24164 23054
rect 24108 22990 24110 23042
rect 24162 22990 24164 23042
rect 23884 21924 23940 22540
rect 23884 21858 23940 21868
rect 23996 22370 24052 22382
rect 23996 22318 23998 22370
rect 24050 22318 24052 22370
rect 23996 21810 24052 22318
rect 24108 22036 24164 22990
rect 24108 21970 24164 21980
rect 24444 22370 24500 23772
rect 24556 23380 24612 24668
rect 24556 23378 24724 23380
rect 24556 23326 24558 23378
rect 24610 23326 24724 23378
rect 24556 23324 24724 23326
rect 24556 23314 24612 23324
rect 24444 22318 24446 22370
rect 24498 22318 24500 22370
rect 23996 21758 23998 21810
rect 24050 21758 24052 21810
rect 23996 21746 24052 21758
rect 24108 21812 24164 21822
rect 24108 21718 24164 21756
rect 24332 21700 24388 21710
rect 24220 21644 24332 21700
rect 23772 21588 23828 21598
rect 23772 20916 23828 21532
rect 23884 21586 23940 21598
rect 23884 21534 23886 21586
rect 23938 21534 23940 21586
rect 23884 21476 23940 21534
rect 23884 21410 23940 21420
rect 23772 20850 23828 20860
rect 24220 20914 24276 21644
rect 24332 21606 24388 21644
rect 24444 21026 24500 22318
rect 24444 20974 24446 21026
rect 24498 20974 24500 21026
rect 24444 20962 24500 20974
rect 24556 22258 24612 22270
rect 24556 22206 24558 22258
rect 24610 22206 24612 22258
rect 24220 20862 24222 20914
rect 24274 20862 24276 20914
rect 24220 20850 24276 20862
rect 23996 19908 24052 19918
rect 23996 19460 24052 19852
rect 24556 19572 24612 22206
rect 24668 21588 24724 23324
rect 24668 21522 24724 21532
rect 24668 21252 24724 21262
rect 24668 20914 24724 21196
rect 24668 20862 24670 20914
rect 24722 20862 24724 20914
rect 24668 20850 24724 20862
rect 23996 19394 24052 19404
rect 24332 19516 24612 19572
rect 24668 20356 24724 20366
rect 23772 19010 23828 19022
rect 23772 18958 23774 19010
rect 23826 18958 23828 19010
rect 23772 18676 23828 18958
rect 24220 19010 24276 19022
rect 24220 18958 24222 19010
rect 24274 18958 24276 19010
rect 24220 18900 24276 18958
rect 24220 18834 24276 18844
rect 23772 18610 23828 18620
rect 23884 18452 23940 18462
rect 23660 18450 23940 18452
rect 23660 18398 23886 18450
rect 23938 18398 23940 18450
rect 23660 18396 23940 18398
rect 23884 18386 23940 18396
rect 23996 18450 24052 18462
rect 23996 18398 23998 18450
rect 24050 18398 24052 18450
rect 23324 18274 23380 18284
rect 23996 18116 24052 18398
rect 23996 18050 24052 18060
rect 23324 17892 23380 17902
rect 23212 17890 23380 17892
rect 23212 17838 23326 17890
rect 23378 17838 23380 17890
rect 23212 17836 23380 17838
rect 23100 17780 23156 17818
rect 23100 17714 23156 17724
rect 23212 17556 23268 17836
rect 23324 17826 23380 17836
rect 22764 17554 23044 17556
rect 22764 17502 22766 17554
rect 22818 17502 23044 17554
rect 22764 17500 23044 17502
rect 23100 17500 23268 17556
rect 22764 17490 22820 17500
rect 23100 17220 23156 17500
rect 23772 17444 23828 17454
rect 23548 17442 23828 17444
rect 23548 17390 23774 17442
rect 23826 17390 23828 17442
rect 23548 17388 23828 17390
rect 23100 17106 23156 17164
rect 23100 17054 23102 17106
rect 23154 17054 23156 17106
rect 23100 17042 23156 17054
rect 23212 17332 23268 17342
rect 22428 14924 22708 14980
rect 22876 16996 22932 17006
rect 22876 15428 22932 16940
rect 22428 12290 22484 14924
rect 22764 13748 22820 13758
rect 22428 12238 22430 12290
rect 22482 12238 22484 12290
rect 22428 12226 22484 12238
rect 22652 13746 22820 13748
rect 22652 13694 22766 13746
rect 22818 13694 22820 13746
rect 22652 13692 22820 13694
rect 22652 12852 22708 13692
rect 22764 13682 22820 13692
rect 22876 13524 22932 15372
rect 23100 13860 23156 13870
rect 23100 13766 23156 13804
rect 22988 13746 23044 13758
rect 22988 13694 22990 13746
rect 23042 13694 23044 13746
rect 22988 13636 23044 13694
rect 23212 13636 23268 17276
rect 23324 16994 23380 17006
rect 23324 16942 23326 16994
rect 23378 16942 23380 16994
rect 23324 13860 23380 16942
rect 23548 15652 23604 17388
rect 23772 17378 23828 17388
rect 24108 17442 24164 17454
rect 24108 17390 24110 17442
rect 24162 17390 24164 17442
rect 24108 17332 24164 17390
rect 24108 17266 24164 17276
rect 24332 17108 24388 19516
rect 24668 18338 24724 20300
rect 24668 18286 24670 18338
rect 24722 18286 24724 18338
rect 24556 17444 24612 17454
rect 24556 17350 24612 17388
rect 24668 17332 24724 18286
rect 24668 17266 24724 17276
rect 23996 17052 24332 17108
rect 23660 16882 23716 16894
rect 23660 16830 23662 16882
rect 23714 16830 23716 16882
rect 23660 16660 23716 16830
rect 23660 16594 23716 16604
rect 23436 15540 23492 15550
rect 23548 15540 23604 15596
rect 23436 15538 23604 15540
rect 23436 15486 23438 15538
rect 23490 15486 23604 15538
rect 23436 15484 23604 15486
rect 23436 15474 23492 15484
rect 23996 15428 24052 17052
rect 24332 17014 24388 17052
rect 24444 16996 24500 17006
rect 24444 16902 24500 16940
rect 23996 15362 24052 15372
rect 24108 16882 24164 16894
rect 24108 16830 24110 16882
rect 24162 16830 24164 16882
rect 23324 13794 23380 13804
rect 23436 15316 23492 15326
rect 23436 13636 23492 15260
rect 23660 15316 23716 15354
rect 23660 15250 23716 15260
rect 24108 15314 24164 16830
rect 24332 16660 24388 16670
rect 24108 15262 24110 15314
rect 24162 15262 24164 15314
rect 24108 15250 24164 15262
rect 24220 15986 24276 15998
rect 24220 15934 24222 15986
rect 24274 15934 24276 15986
rect 23548 15202 23604 15214
rect 23548 15150 23550 15202
rect 23602 15150 23604 15202
rect 23548 15148 23604 15150
rect 24220 15148 24276 15934
rect 23548 15092 24276 15148
rect 23772 14980 23828 14990
rect 22988 13570 23044 13580
rect 23100 13580 23268 13636
rect 23324 13580 23492 13636
rect 23660 14924 23772 14980
rect 22876 13458 22932 13468
rect 22988 12964 23044 12974
rect 22540 11284 22596 11294
rect 22540 11190 22596 11228
rect 22316 11116 22484 11172
rect 22316 10948 22372 10958
rect 22204 10612 22260 10622
rect 22316 10612 22372 10892
rect 22260 10556 22372 10612
rect 22204 10518 22260 10556
rect 22092 9650 22148 9660
rect 21644 9100 21812 9156
rect 21644 8932 21700 8942
rect 21532 8930 21700 8932
rect 21532 8878 21646 8930
rect 21698 8878 21700 8930
rect 21532 8876 21700 8878
rect 21644 8866 21700 8876
rect 21420 8372 21476 8382
rect 20748 8370 21476 8372
rect 20748 8318 21422 8370
rect 21474 8318 21476 8370
rect 20748 8316 21476 8318
rect 20076 8260 20132 8270
rect 20076 7812 20132 8204
rect 20748 8258 20804 8316
rect 21420 8306 21476 8316
rect 20748 8206 20750 8258
rect 20802 8206 20804 8258
rect 20748 8194 20804 8206
rect 21756 8260 21812 9100
rect 21756 8194 21812 8204
rect 21980 8260 22036 8270
rect 20188 8148 20244 8158
rect 20412 8148 20468 8158
rect 20188 8146 20468 8148
rect 20188 8094 20190 8146
rect 20242 8094 20414 8146
rect 20466 8094 20468 8146
rect 20188 8092 20468 8094
rect 20188 8082 20244 8092
rect 20412 8082 20468 8092
rect 20636 8036 20692 8046
rect 20636 8034 20916 8036
rect 20636 7982 20638 8034
rect 20690 7982 20916 8034
rect 20636 7980 20916 7982
rect 20636 7970 20692 7980
rect 20532 7868 20796 7878
rect 20588 7812 20636 7868
rect 20692 7812 20740 7868
rect 20076 7756 20468 7812
rect 20532 7802 20796 7812
rect 20412 7700 20468 7756
rect 20524 7700 20580 7710
rect 20412 7698 20580 7700
rect 20412 7646 20526 7698
rect 20578 7646 20580 7698
rect 20412 7644 20580 7646
rect 20524 7634 20580 7644
rect 20188 7476 20244 7486
rect 20244 7420 20356 7476
rect 20188 7410 20244 7420
rect 20188 7028 20244 7038
rect 20076 6580 20132 6590
rect 19740 6132 19796 6524
rect 19740 6038 19796 6076
rect 19852 6578 20132 6580
rect 19852 6526 20078 6578
rect 20130 6526 20132 6578
rect 19852 6524 20132 6526
rect 19852 4338 19908 6524
rect 20076 6514 20132 6524
rect 19964 6020 20020 6030
rect 19964 5906 20020 5964
rect 19964 5854 19966 5906
rect 20018 5854 20020 5906
rect 19964 5842 20020 5854
rect 19852 4286 19854 4338
rect 19906 4286 19908 4338
rect 19852 4274 19908 4286
rect 20188 3668 20244 6972
rect 20300 6804 20356 7420
rect 20300 5796 20356 6748
rect 20412 6580 20468 6590
rect 20412 6486 20468 6524
rect 20532 6300 20796 6310
rect 20588 6244 20636 6300
rect 20692 6244 20740 6300
rect 20532 6234 20796 6244
rect 20412 6020 20468 6030
rect 20412 5926 20468 5964
rect 20636 5906 20692 5918
rect 20636 5854 20638 5906
rect 20690 5854 20692 5906
rect 20636 5796 20692 5854
rect 20300 5740 20692 5796
rect 20748 5684 20804 5694
rect 20748 5122 20804 5628
rect 20748 5070 20750 5122
rect 20802 5070 20804 5122
rect 20748 5058 20804 5070
rect 20412 4898 20468 4910
rect 20412 4846 20414 4898
rect 20466 4846 20468 4898
rect 20412 4452 20468 4846
rect 20532 4732 20796 4742
rect 20588 4676 20636 4732
rect 20692 4676 20740 4732
rect 20532 4666 20796 4676
rect 20636 4452 20692 4462
rect 20412 4450 20692 4452
rect 20412 4398 20638 4450
rect 20690 4398 20692 4450
rect 20412 4396 20692 4398
rect 20636 4386 20692 4396
rect 20188 3602 20244 3612
rect 19628 3266 19684 3276
rect 19740 3556 19796 3566
rect 19740 800 19796 3500
rect 20300 3556 20356 3566
rect 20300 3462 20356 3500
rect 20748 3444 20804 3454
rect 20860 3444 20916 7980
rect 21980 7588 22036 8204
rect 21532 7532 22036 7588
rect 21308 6804 21364 6814
rect 21308 6466 21364 6748
rect 21308 6414 21310 6466
rect 21362 6414 21364 6466
rect 21308 6130 21364 6414
rect 21308 6078 21310 6130
rect 21362 6078 21364 6130
rect 21308 6066 21364 6078
rect 21532 5122 21588 7532
rect 22428 7028 22484 11116
rect 22652 11060 22708 12796
rect 22876 12908 22988 12964
rect 22876 12178 22932 12908
rect 22988 12870 23044 12908
rect 22876 12126 22878 12178
rect 22930 12126 22932 12178
rect 22876 12114 22932 12126
rect 22764 11396 22820 11406
rect 22764 11302 22820 11340
rect 22876 11172 22932 11182
rect 22876 11078 22932 11116
rect 22988 11170 23044 11182
rect 22988 11118 22990 11170
rect 23042 11118 23044 11170
rect 22428 6962 22484 6972
rect 22540 11004 22708 11060
rect 21644 6580 21700 6590
rect 21644 6486 21700 6524
rect 21980 6020 22036 6030
rect 21980 6018 22260 6020
rect 21980 5966 21982 6018
rect 22034 5966 22260 6018
rect 21980 5964 22260 5966
rect 21980 5954 22036 5964
rect 21532 5070 21534 5122
rect 21586 5070 21588 5122
rect 21532 5058 21588 5070
rect 21756 5906 21812 5918
rect 21756 5854 21758 5906
rect 21810 5854 21812 5906
rect 21756 4564 21812 5854
rect 22204 5234 22260 5964
rect 22428 5684 22484 5694
rect 22540 5684 22596 11004
rect 22652 10724 22708 10734
rect 22652 10630 22708 10668
rect 22764 10500 22820 10510
rect 22764 9938 22820 10444
rect 22876 10164 22932 10174
rect 22988 10164 23044 11118
rect 22932 10108 23044 10164
rect 22876 10098 22932 10108
rect 22764 9886 22766 9938
rect 22818 9886 22820 9938
rect 22764 9874 22820 9886
rect 22988 9156 23044 9166
rect 22764 9154 23044 9156
rect 22764 9102 22990 9154
rect 23042 9102 23044 9154
rect 22764 9100 23044 9102
rect 22764 8370 22820 9100
rect 22988 9090 23044 9100
rect 22764 8318 22766 8370
rect 22818 8318 22820 8370
rect 22764 8306 22820 8318
rect 22764 5684 22820 5694
rect 22540 5682 22820 5684
rect 22540 5630 22766 5682
rect 22818 5630 22820 5682
rect 22540 5628 22820 5630
rect 22428 5590 22484 5628
rect 22204 5182 22206 5234
rect 22258 5182 22260 5234
rect 22204 5170 22260 5182
rect 21756 4498 21812 4508
rect 22764 4226 22820 5628
rect 23100 5012 23156 13580
rect 23212 12516 23268 12526
rect 23212 12402 23268 12460
rect 23212 12350 23214 12402
rect 23266 12350 23268 12402
rect 23212 11394 23268 12350
rect 23212 11342 23214 11394
rect 23266 11342 23268 11394
rect 23212 10834 23268 11342
rect 23212 10782 23214 10834
rect 23266 10782 23268 10834
rect 23212 10770 23268 10782
rect 23324 10164 23380 13580
rect 23548 13524 23604 13534
rect 23548 13430 23604 13468
rect 23660 12628 23716 14924
rect 23772 14914 23828 14924
rect 24220 14196 24276 14206
rect 23996 13860 24052 13870
rect 23996 13766 24052 13804
rect 24108 13636 24164 13646
rect 23996 13580 24108 13636
rect 23772 12740 23828 12750
rect 23772 12646 23828 12684
rect 23660 12562 23716 12572
rect 23884 12292 23940 12302
rect 23660 12066 23716 12078
rect 23660 12014 23662 12066
rect 23714 12014 23716 12066
rect 23660 11732 23716 12014
rect 23436 11676 23660 11732
rect 23436 11396 23492 11676
rect 23660 11666 23716 11676
rect 23884 11620 23940 12236
rect 23884 11554 23940 11564
rect 23996 12290 24052 13580
rect 24108 13570 24164 13580
rect 24220 13074 24276 14140
rect 24332 13970 24388 16604
rect 24332 13918 24334 13970
rect 24386 13918 24388 13970
rect 24332 13906 24388 13918
rect 24444 16212 24500 16222
rect 24444 15426 24500 16156
rect 24444 15374 24446 15426
rect 24498 15374 24500 15426
rect 24220 13022 24222 13074
rect 24274 13022 24276 13074
rect 24220 13010 24276 13022
rect 24332 13188 24388 13198
rect 24444 13188 24500 15374
rect 24556 15316 24612 15326
rect 24556 15222 24612 15260
rect 24780 14980 24836 27244
rect 24892 19460 24948 28364
rect 25004 27300 25060 29148
rect 25228 28196 25284 29260
rect 25228 28130 25284 28140
rect 25004 27234 25060 27244
rect 25228 27858 25284 27870
rect 25228 27806 25230 27858
rect 25282 27806 25284 27858
rect 25116 27188 25172 27198
rect 25228 27188 25284 27806
rect 25172 27132 25284 27188
rect 25116 27094 25172 27132
rect 25004 25508 25060 25518
rect 25004 25414 25060 25452
rect 25228 24276 25284 24286
rect 25228 24050 25284 24220
rect 25228 23998 25230 24050
rect 25282 23998 25284 24050
rect 25004 22370 25060 22382
rect 25004 22318 25006 22370
rect 25058 22318 25060 22370
rect 25004 22036 25060 22318
rect 25004 21970 25060 21980
rect 25228 21252 25284 23998
rect 25340 23378 25396 30604
rect 25452 30212 25508 30222
rect 25452 28866 25508 30156
rect 25564 29426 25620 30828
rect 25900 30436 25956 30942
rect 26124 31778 26292 31780
rect 26124 31726 26238 31778
rect 26290 31726 26292 31778
rect 26124 31724 26292 31726
rect 26012 30884 26068 30894
rect 26124 30884 26180 31724
rect 26236 31714 26292 31724
rect 26460 31778 26516 31790
rect 26460 31726 26462 31778
rect 26514 31726 26516 31778
rect 26460 31556 26516 31726
rect 26460 31490 26516 31500
rect 26236 31108 26292 31118
rect 26236 30994 26292 31052
rect 26236 30942 26238 30994
rect 26290 30942 26292 30994
rect 26236 30930 26292 30942
rect 26068 30828 26180 30884
rect 26012 30818 26068 30828
rect 26012 30436 26068 30446
rect 25900 30434 26068 30436
rect 25900 30382 26014 30434
rect 26066 30382 26068 30434
rect 25900 30380 26068 30382
rect 26012 30370 26068 30380
rect 25788 30322 25844 30334
rect 25788 30270 25790 30322
rect 25842 30270 25844 30322
rect 25564 29374 25566 29426
rect 25618 29374 25620 29426
rect 25564 29362 25620 29374
rect 25676 30210 25732 30222
rect 25676 30158 25678 30210
rect 25730 30158 25732 30210
rect 25452 28814 25454 28866
rect 25506 28814 25508 28866
rect 25452 28082 25508 28814
rect 25676 28644 25732 30158
rect 25788 28866 25844 30270
rect 26012 30212 26068 30222
rect 25788 28814 25790 28866
rect 25842 28814 25844 28866
rect 25788 28802 25844 28814
rect 25900 30156 26012 30212
rect 25452 28030 25454 28082
rect 25506 28030 25508 28082
rect 25452 28018 25508 28030
rect 25564 28588 25732 28644
rect 25788 28644 25844 28654
rect 25900 28644 25956 30156
rect 26012 30146 26068 30156
rect 26572 29988 26628 32396
rect 26684 31778 26740 31790
rect 26684 31726 26686 31778
rect 26738 31726 26740 31778
rect 26684 30436 26740 31726
rect 27356 31668 27412 31678
rect 27356 31574 27412 31612
rect 27132 31556 27188 31566
rect 27132 31462 27188 31500
rect 26684 30370 26740 30380
rect 26796 30100 26852 30110
rect 25788 28642 25956 28644
rect 25788 28590 25790 28642
rect 25842 28590 25956 28642
rect 25788 28588 25956 28590
rect 26012 29932 26628 29988
rect 26684 29986 26740 29998
rect 26684 29934 26686 29986
rect 26738 29934 26740 29986
rect 25564 28084 25620 28588
rect 25788 28578 25844 28588
rect 25564 28018 25620 28028
rect 25900 27970 25956 27982
rect 25900 27918 25902 27970
rect 25954 27918 25956 27970
rect 25900 27748 25956 27918
rect 25900 27682 25956 27692
rect 25900 27524 25956 27534
rect 25788 27188 25844 27198
rect 25788 27074 25844 27132
rect 25788 27022 25790 27074
rect 25842 27022 25844 27074
rect 25788 27010 25844 27022
rect 25564 26964 25620 26974
rect 25564 25956 25620 26908
rect 25900 26514 25956 27468
rect 26012 26908 26068 29932
rect 26124 29540 26180 29550
rect 26124 27188 26180 29484
rect 26460 29538 26516 29550
rect 26460 29486 26462 29538
rect 26514 29486 26516 29538
rect 26460 29428 26516 29486
rect 26460 29362 26516 29372
rect 26572 29426 26628 29438
rect 26572 29374 26574 29426
rect 26626 29374 26628 29426
rect 26236 28756 26292 28766
rect 26236 28642 26292 28700
rect 26236 28590 26238 28642
rect 26290 28590 26292 28642
rect 26236 28578 26292 28590
rect 26460 28532 26516 28542
rect 26460 28438 26516 28476
rect 26572 28530 26628 29374
rect 26684 29316 26740 29934
rect 26796 29540 26852 30044
rect 26796 29474 26852 29484
rect 27132 29538 27188 29550
rect 27132 29486 27134 29538
rect 27186 29486 27188 29538
rect 27132 29428 27188 29486
rect 27132 29362 27188 29372
rect 26684 29250 26740 29260
rect 26572 28478 26574 28530
rect 26626 28478 26628 28530
rect 26572 28308 26628 28478
rect 27132 28530 27188 28542
rect 27132 28478 27134 28530
rect 27186 28478 27188 28530
rect 26796 28420 26852 28430
rect 26572 28242 26628 28252
rect 26684 28418 26852 28420
rect 26684 28366 26798 28418
rect 26850 28366 26852 28418
rect 26684 28364 26852 28366
rect 26348 28084 26404 28094
rect 26348 27858 26404 28028
rect 26348 27806 26350 27858
rect 26402 27806 26404 27858
rect 26348 27794 26404 27806
rect 26684 27636 26740 28364
rect 26796 28354 26852 28364
rect 27020 28418 27076 28430
rect 27020 28366 27022 28418
rect 27074 28366 27076 28418
rect 26908 28308 26964 28318
rect 26796 27748 26852 27758
rect 26796 27654 26852 27692
rect 26348 27580 26740 27636
rect 26124 27132 26292 27188
rect 26236 26908 26292 27132
rect 26348 27074 26404 27580
rect 26684 27412 26740 27422
rect 26348 27022 26350 27074
rect 26402 27022 26404 27074
rect 26348 27010 26404 27022
rect 26572 27300 26628 27310
rect 26460 26962 26516 26974
rect 26460 26910 26462 26962
rect 26514 26910 26516 26962
rect 26460 26908 26516 26910
rect 26012 26852 26180 26908
rect 26236 26852 26516 26908
rect 25900 26462 25902 26514
rect 25954 26462 25956 26514
rect 25900 26450 25956 26462
rect 26124 26402 26180 26852
rect 26124 26350 26126 26402
rect 26178 26350 26180 26402
rect 25676 26180 25732 26190
rect 26124 26180 26180 26350
rect 26236 26404 26292 26414
rect 26572 26404 26628 27244
rect 26684 27074 26740 27356
rect 26684 27022 26686 27074
rect 26738 27022 26740 27074
rect 26684 27010 26740 27022
rect 26796 27188 26852 27198
rect 26796 26964 26852 27132
rect 26908 27076 26964 28252
rect 27020 27748 27076 28366
rect 27132 28084 27188 28478
rect 27468 28308 27524 32844
rect 27580 29426 27636 36204
rect 27692 36194 27748 36204
rect 28252 35922 28308 36428
rect 29148 36482 29204 36540
rect 29148 36430 29150 36482
rect 29202 36430 29204 36482
rect 29148 36418 29204 36430
rect 29596 37044 29652 37054
rect 28812 36372 28868 36382
rect 28700 36260 28756 36270
rect 28700 36166 28756 36204
rect 28812 36036 28868 36316
rect 28924 36260 28980 36270
rect 28924 36166 28980 36204
rect 29372 36260 29428 36270
rect 28812 35980 28980 36036
rect 28252 35870 28254 35922
rect 28306 35870 28308 35922
rect 28252 35858 28308 35870
rect 28812 35812 28868 35822
rect 28588 35810 28868 35812
rect 28588 35758 28814 35810
rect 28866 35758 28868 35810
rect 28588 35756 28868 35758
rect 27804 35028 27860 35038
rect 27692 34692 27748 34702
rect 27692 34354 27748 34636
rect 27692 34302 27694 34354
rect 27746 34302 27748 34354
rect 27692 34290 27748 34302
rect 27692 31554 27748 31566
rect 27692 31502 27694 31554
rect 27746 31502 27748 31554
rect 27692 30212 27748 31502
rect 27692 30146 27748 30156
rect 27580 29374 27582 29426
rect 27634 29374 27636 29426
rect 27580 28532 27636 29374
rect 27804 29092 27860 34972
rect 28364 34914 28420 34926
rect 28364 34862 28366 34914
rect 28418 34862 28420 34914
rect 28028 34690 28084 34702
rect 28028 34638 28030 34690
rect 28082 34638 28084 34690
rect 28028 34244 28084 34638
rect 28364 34692 28420 34862
rect 28364 34626 28420 34636
rect 28588 34690 28644 35756
rect 28812 35746 28868 35756
rect 28700 35588 28756 35598
rect 28924 35588 28980 35980
rect 29036 35700 29092 35710
rect 29036 35698 29204 35700
rect 29036 35646 29038 35698
rect 29090 35646 29204 35698
rect 29036 35644 29204 35646
rect 29036 35634 29092 35644
rect 28700 35586 28980 35588
rect 28700 35534 28702 35586
rect 28754 35534 28980 35586
rect 28700 35532 28980 35534
rect 28700 35476 28756 35532
rect 28700 35410 28756 35420
rect 29148 35476 29204 35644
rect 29148 35410 29204 35420
rect 29260 35588 29316 35598
rect 29036 35364 29092 35374
rect 28588 34638 28590 34690
rect 28642 34638 28644 34690
rect 28364 34356 28420 34366
rect 28364 34244 28420 34300
rect 28028 34188 28420 34244
rect 27916 34018 27972 34030
rect 27916 33966 27918 34018
rect 27970 33966 27972 34018
rect 27916 33236 27972 33966
rect 28028 34020 28084 34030
rect 28028 33926 28084 33964
rect 28252 33348 28308 33358
rect 28252 33254 28308 33292
rect 28140 33236 28196 33246
rect 27916 33180 28140 33236
rect 28140 32900 28196 33180
rect 28140 32844 28308 32900
rect 28252 32674 28308 32844
rect 28252 32622 28254 32674
rect 28306 32622 28308 32674
rect 28252 32610 28308 32622
rect 28140 32562 28196 32574
rect 28140 32510 28142 32562
rect 28194 32510 28196 32562
rect 27916 32452 27972 32462
rect 28140 32452 28196 32510
rect 27916 32450 28196 32452
rect 27916 32398 27918 32450
rect 27970 32398 28196 32450
rect 27916 32396 28196 32398
rect 27916 32004 27972 32396
rect 28364 32340 28420 34188
rect 28588 34244 28644 34638
rect 28588 34178 28644 34188
rect 28700 35252 28756 35262
rect 28700 34020 28756 35196
rect 28924 34916 28980 34926
rect 28812 34804 28868 34814
rect 28812 34242 28868 34748
rect 28812 34190 28814 34242
rect 28866 34190 28868 34242
rect 28812 34178 28868 34190
rect 28924 34130 28980 34860
rect 28924 34078 28926 34130
rect 28978 34078 28980 34130
rect 28924 34066 28980 34078
rect 28700 33964 28868 34020
rect 27916 31938 27972 31948
rect 28140 32284 28420 32340
rect 28588 33460 28644 33470
rect 28588 33122 28644 33404
rect 28588 33070 28590 33122
rect 28642 33070 28644 33122
rect 28140 30548 28196 32284
rect 28588 31668 28644 33070
rect 28588 31602 28644 31612
rect 28252 31444 28308 31454
rect 28252 30996 28308 31388
rect 28588 30996 28644 31006
rect 28252 30994 28420 30996
rect 28252 30942 28254 30994
rect 28306 30942 28420 30994
rect 28252 30940 28420 30942
rect 28252 30930 28308 30940
rect 28028 29316 28084 29326
rect 28028 29222 28084 29260
rect 27804 29036 28084 29092
rect 27580 28466 27636 28476
rect 27916 28642 27972 28654
rect 27916 28590 27918 28642
rect 27970 28590 27972 28642
rect 27468 28242 27524 28252
rect 27132 28018 27188 28028
rect 27804 28084 27860 28094
rect 27804 27990 27860 28028
rect 27020 27682 27076 27692
rect 27356 27746 27412 27758
rect 27356 27694 27358 27746
rect 27410 27694 27412 27746
rect 27132 27636 27188 27646
rect 27020 27076 27076 27114
rect 26908 27020 27020 27076
rect 27020 27010 27076 27020
rect 26796 26908 26964 26964
rect 27132 26908 27188 27580
rect 27356 27188 27412 27694
rect 27356 27122 27412 27132
rect 26908 26850 26964 26908
rect 26908 26798 26910 26850
rect 26962 26798 26964 26850
rect 26908 26786 26964 26798
rect 27020 26852 27188 26908
rect 27468 27076 27524 27086
rect 26236 26310 26292 26348
rect 26460 26348 26628 26404
rect 25676 26178 26180 26180
rect 25676 26126 25678 26178
rect 25730 26126 26180 26178
rect 25676 26124 26180 26126
rect 25676 26114 25732 26124
rect 25564 25900 26068 25956
rect 25900 25396 25956 25406
rect 25900 24948 25956 25340
rect 26012 25394 26068 25900
rect 26012 25342 26014 25394
rect 26066 25342 26068 25394
rect 26012 25330 26068 25342
rect 26012 24948 26068 24958
rect 25900 24946 26068 24948
rect 25900 24894 26014 24946
rect 26066 24894 26068 24946
rect 25900 24892 26068 24894
rect 26012 24882 26068 24892
rect 26012 24276 26068 24286
rect 26012 24050 26068 24220
rect 26012 23998 26014 24050
rect 26066 23998 26068 24050
rect 26012 23986 26068 23998
rect 25788 23714 25844 23726
rect 25788 23662 25790 23714
rect 25842 23662 25844 23714
rect 25340 23326 25342 23378
rect 25394 23326 25396 23378
rect 25340 23314 25396 23326
rect 25452 23604 25508 23614
rect 25228 21196 25396 21252
rect 25116 21026 25172 21038
rect 25116 20974 25118 21026
rect 25170 20974 25172 21026
rect 25116 20914 25172 20974
rect 25116 20862 25118 20914
rect 25170 20862 25172 20914
rect 25116 20850 25172 20862
rect 25228 21028 25284 21038
rect 24892 19394 24948 19404
rect 25004 20580 25060 20590
rect 24892 19124 24948 19134
rect 25004 19124 25060 20524
rect 25228 19908 25284 20972
rect 25340 21026 25396 21196
rect 25340 20974 25342 21026
rect 25394 20974 25396 21026
rect 25340 20962 25396 20974
rect 25228 19842 25284 19852
rect 24892 19122 25060 19124
rect 24892 19070 24894 19122
rect 24946 19070 25060 19122
rect 24892 19068 25060 19070
rect 24892 19058 24948 19068
rect 25228 19012 25284 19022
rect 25228 18918 25284 18956
rect 25004 17892 25060 17902
rect 25004 17778 25060 17836
rect 25004 17726 25006 17778
rect 25058 17726 25060 17778
rect 25004 16436 25060 17726
rect 25340 17108 25396 17118
rect 25340 17014 25396 17052
rect 25004 16370 25060 16380
rect 24780 14914 24836 14924
rect 25004 16098 25060 16110
rect 25004 16046 25006 16098
rect 25058 16046 25060 16098
rect 24892 13860 24948 13870
rect 24444 13132 24836 13188
rect 24332 12964 24388 13132
rect 24444 12964 24500 12974
rect 24332 12962 24500 12964
rect 24332 12910 24446 12962
rect 24498 12910 24500 12962
rect 24332 12908 24500 12910
rect 24444 12898 24500 12908
rect 24220 12852 24276 12862
rect 24220 12758 24276 12796
rect 24668 12852 24724 12862
rect 24780 12852 24836 13132
rect 24892 13076 24948 13804
rect 25004 13300 25060 16046
rect 25340 15316 25396 15326
rect 25340 15222 25396 15260
rect 25452 14308 25508 23548
rect 25676 23604 25732 23614
rect 25564 23492 25620 23502
rect 25564 21700 25620 23436
rect 25676 23156 25732 23548
rect 25676 23062 25732 23100
rect 25788 22484 25844 23662
rect 26124 23492 26180 26124
rect 26348 25620 26404 25630
rect 26348 25506 26404 25564
rect 26348 25454 26350 25506
rect 26402 25454 26404 25506
rect 26348 25442 26404 25454
rect 26348 23828 26404 23838
rect 26348 23734 26404 23772
rect 26124 23426 26180 23436
rect 26460 23380 26516 26348
rect 26684 26292 26740 26302
rect 26684 26178 26740 26236
rect 26684 26126 26686 26178
rect 26738 26126 26740 26178
rect 26684 26114 26740 26126
rect 26908 25620 26964 25630
rect 26908 25396 26964 25564
rect 26908 25302 26964 25340
rect 26796 24610 26852 24622
rect 26796 24558 26798 24610
rect 26850 24558 26852 24610
rect 26684 23714 26740 23726
rect 26684 23662 26686 23714
rect 26738 23662 26740 23714
rect 26684 23492 26740 23662
rect 26684 23426 26740 23436
rect 26236 23268 26292 23278
rect 26460 23268 26516 23324
rect 26236 23266 26516 23268
rect 26236 23214 26238 23266
rect 26290 23214 26516 23266
rect 26236 23212 26516 23214
rect 26236 23202 26292 23212
rect 26684 23156 26740 23166
rect 26796 23156 26852 24558
rect 27020 23940 27076 26852
rect 27132 26292 27188 26302
rect 27468 26292 27524 27020
rect 27580 27076 27636 27086
rect 27916 27076 27972 28590
rect 28028 28308 28084 29036
rect 28140 28530 28196 30492
rect 28364 30322 28420 30940
rect 28588 30902 28644 30940
rect 28364 30270 28366 30322
rect 28418 30270 28420 30322
rect 28364 30258 28420 30270
rect 28252 30212 28308 30222
rect 28252 30118 28308 30156
rect 28364 30098 28420 30110
rect 28364 30046 28366 30098
rect 28418 30046 28420 30098
rect 28364 29988 28420 30046
rect 28420 29932 28532 29988
rect 28364 29922 28420 29932
rect 28140 28478 28142 28530
rect 28194 28478 28196 28530
rect 28140 28466 28196 28478
rect 28028 28252 28308 28308
rect 28028 28084 28084 28094
rect 28028 27990 28084 28028
rect 27580 27074 27972 27076
rect 27580 27022 27582 27074
rect 27634 27022 27972 27074
rect 27580 27020 27972 27022
rect 27580 27010 27636 27020
rect 27132 26198 27188 26236
rect 27356 26290 27524 26292
rect 27356 26238 27470 26290
rect 27522 26238 27524 26290
rect 27356 26236 27524 26238
rect 27132 25396 27188 25406
rect 27356 25396 27412 26236
rect 27468 26226 27524 26236
rect 27692 26404 27748 26414
rect 27468 25508 27524 25518
rect 27468 25414 27524 25452
rect 27132 25394 27412 25396
rect 27132 25342 27134 25394
rect 27186 25342 27412 25394
rect 27132 25340 27412 25342
rect 27132 25330 27188 25340
rect 26348 23154 26852 23156
rect 26348 23102 26686 23154
rect 26738 23102 26852 23154
rect 26348 23100 26852 23102
rect 26908 23884 27076 23940
rect 27244 25172 27300 25182
rect 27244 24946 27300 25116
rect 27244 24894 27246 24946
rect 27298 24894 27300 24946
rect 26012 23044 26068 23054
rect 26012 22950 26068 22988
rect 26348 22596 26404 23100
rect 26684 23090 26740 23100
rect 26348 22502 26404 22540
rect 25788 22418 25844 22428
rect 26572 22484 26628 22494
rect 26460 22370 26516 22382
rect 26460 22318 26462 22370
rect 26514 22318 26516 22370
rect 25676 22258 25732 22270
rect 25676 22206 25678 22258
rect 25730 22206 25732 22258
rect 25676 21924 25732 22206
rect 25788 22148 25844 22158
rect 26012 22148 26068 22158
rect 25788 22146 25956 22148
rect 25788 22094 25790 22146
rect 25842 22094 25956 22146
rect 25788 22092 25956 22094
rect 25788 22082 25844 22092
rect 25676 21858 25732 21868
rect 25900 21812 25956 22092
rect 26012 22054 26068 22092
rect 25564 21644 25732 21700
rect 25564 21476 25620 21486
rect 25564 21382 25620 21420
rect 25564 21026 25620 21038
rect 25564 20974 25566 21026
rect 25618 20974 25620 21026
rect 25564 20692 25620 20974
rect 25676 20914 25732 21644
rect 25676 20862 25678 20914
rect 25730 20862 25732 20914
rect 25676 20850 25732 20862
rect 25788 21476 25844 21486
rect 25788 20804 25844 21420
rect 25900 21364 25956 21756
rect 26124 21588 26180 21598
rect 26124 21494 26180 21532
rect 26460 21588 26516 22318
rect 26572 22370 26628 22428
rect 26572 22318 26574 22370
rect 26626 22318 26628 22370
rect 26572 22260 26628 22318
rect 26628 22204 26740 22260
rect 26572 22194 26628 22204
rect 26460 21494 26516 21532
rect 26684 21698 26740 22204
rect 26684 21646 26686 21698
rect 26738 21646 26740 21698
rect 25900 21308 26292 21364
rect 25900 20804 25956 20814
rect 25788 20802 25956 20804
rect 25788 20750 25902 20802
rect 25954 20750 25956 20802
rect 25788 20748 25956 20750
rect 25564 20636 25844 20692
rect 25788 20356 25844 20636
rect 25900 20580 25956 20748
rect 26236 20804 26292 21308
rect 26236 20690 26292 20748
rect 26236 20638 26238 20690
rect 26290 20638 26292 20690
rect 26236 20626 26292 20638
rect 25900 20514 25956 20524
rect 26572 20578 26628 20590
rect 26572 20526 26574 20578
rect 26626 20526 26628 20578
rect 26572 20468 26628 20526
rect 26124 20412 26628 20468
rect 26124 20356 26180 20412
rect 25788 20300 26180 20356
rect 25788 20242 25844 20300
rect 25788 20190 25790 20242
rect 25842 20190 25844 20242
rect 25788 20178 25844 20190
rect 26236 20020 26292 20412
rect 26684 20356 26740 21646
rect 26348 20300 26740 20356
rect 26796 21924 26852 21934
rect 26348 20242 26404 20300
rect 26348 20190 26350 20242
rect 26402 20190 26404 20242
rect 26348 20178 26404 20190
rect 26236 19964 26628 20020
rect 26572 19684 26628 19964
rect 26684 19908 26740 19918
rect 26796 19908 26852 21868
rect 26908 20132 26964 23884
rect 27020 23714 27076 23726
rect 27020 23662 27022 23714
rect 27074 23662 27076 23714
rect 27020 21812 27076 23662
rect 27244 23604 27300 24894
rect 27244 23538 27300 23548
rect 27468 24836 27524 24846
rect 27468 24050 27524 24780
rect 27468 23998 27470 24050
rect 27522 23998 27524 24050
rect 27244 23380 27300 23390
rect 27244 23286 27300 23324
rect 27468 23156 27524 23998
rect 27468 23154 27636 23156
rect 27468 23102 27470 23154
rect 27522 23102 27636 23154
rect 27468 23100 27636 23102
rect 27468 23090 27524 23100
rect 27468 22370 27524 22382
rect 27468 22318 27470 22370
rect 27522 22318 27524 22370
rect 27020 21746 27076 21756
rect 27244 21812 27300 21822
rect 27244 21140 27300 21756
rect 26908 20066 26964 20076
rect 27020 21084 27300 21140
rect 27468 21586 27524 22318
rect 27580 21812 27636 23100
rect 27580 21746 27636 21756
rect 27468 21534 27470 21586
rect 27522 21534 27524 21586
rect 26684 19906 26852 19908
rect 26684 19854 26686 19906
rect 26738 19854 26852 19906
rect 26684 19852 26852 19854
rect 26684 19842 26740 19852
rect 27020 19684 27076 21084
rect 27132 20916 27188 20926
rect 27468 20916 27524 21534
rect 27692 21364 27748 26348
rect 27804 26292 27860 26302
rect 27804 25730 27860 26236
rect 27804 25678 27806 25730
rect 27858 25678 27860 25730
rect 27804 24836 27860 25678
rect 27916 25618 27972 27020
rect 28140 27860 28196 27870
rect 28028 26180 28084 26190
rect 28140 26180 28196 27804
rect 28252 26404 28308 28252
rect 28364 28196 28420 28206
rect 28364 27186 28420 28140
rect 28364 27134 28366 27186
rect 28418 27134 28420 27186
rect 28364 27122 28420 27134
rect 28476 26908 28532 29932
rect 28588 29316 28644 29326
rect 28588 29222 28644 29260
rect 28700 28084 28756 28094
rect 28700 27990 28756 28028
rect 28252 26338 28308 26348
rect 28364 26852 28532 26908
rect 28028 26178 28196 26180
rect 28028 26126 28030 26178
rect 28082 26126 28196 26178
rect 28028 26124 28196 26126
rect 28028 25956 28084 26124
rect 28028 25890 28084 25900
rect 28364 25620 28420 26852
rect 28588 26740 28644 26750
rect 28588 26178 28644 26684
rect 28588 26126 28590 26178
rect 28642 26126 28644 26178
rect 28588 25844 28644 26126
rect 28588 25778 28644 25788
rect 28700 25956 28756 25966
rect 27916 25566 27918 25618
rect 27970 25566 27972 25618
rect 27916 25554 27972 25566
rect 28252 25564 28420 25620
rect 28140 25506 28196 25518
rect 28140 25454 28142 25506
rect 28194 25454 28196 25506
rect 28140 25284 28196 25454
rect 28140 25218 28196 25228
rect 28252 25060 28308 25564
rect 28476 25508 28532 25518
rect 28700 25508 28756 25900
rect 27804 24770 27860 24780
rect 28028 25004 28308 25060
rect 28364 25452 28476 25508
rect 27916 24724 27972 24734
rect 27916 24630 27972 24668
rect 28028 23714 28084 25004
rect 28140 24836 28196 24846
rect 28140 24742 28196 24780
rect 28364 24162 28420 25452
rect 28476 25442 28532 25452
rect 28588 25452 28756 25508
rect 28588 25282 28644 25452
rect 28588 25230 28590 25282
rect 28642 25230 28644 25282
rect 28364 24110 28366 24162
rect 28418 24110 28420 24162
rect 28364 24098 28420 24110
rect 28476 24722 28532 24734
rect 28476 24670 28478 24722
rect 28530 24670 28532 24722
rect 28476 23940 28532 24670
rect 28588 24724 28644 25230
rect 28588 24658 28644 24668
rect 28700 25284 28756 25294
rect 28476 23874 28532 23884
rect 28252 23828 28308 23838
rect 28028 23662 28030 23714
rect 28082 23662 28084 23714
rect 27916 23492 27972 23502
rect 27804 22820 27860 22830
rect 27804 22484 27860 22764
rect 27804 22418 27860 22428
rect 27916 22370 27972 23436
rect 28028 22820 28084 23662
rect 28028 22754 28084 22764
rect 28140 23826 28308 23828
rect 28140 23774 28254 23826
rect 28306 23774 28308 23826
rect 28140 23772 28308 23774
rect 27916 22318 27918 22370
rect 27970 22318 27972 22370
rect 27916 22306 27972 22318
rect 28140 22148 28196 23772
rect 28252 23762 28308 23772
rect 28364 23714 28420 23726
rect 28364 23662 28366 23714
rect 28418 23662 28420 23714
rect 28364 23604 28420 23662
rect 28364 23268 28420 23548
rect 28364 23174 28420 23212
rect 28252 23156 28308 23166
rect 28252 22372 28308 23100
rect 28252 22370 28420 22372
rect 28252 22318 28254 22370
rect 28306 22318 28420 22370
rect 28252 22316 28420 22318
rect 28252 22306 28308 22316
rect 27804 21810 27860 21822
rect 27804 21758 27806 21810
rect 27858 21758 27860 21810
rect 27804 21588 27860 21758
rect 27804 21522 27860 21532
rect 27916 21588 27972 21598
rect 28140 21588 28196 22092
rect 27916 21586 28196 21588
rect 27916 21534 27918 21586
rect 27970 21534 28196 21586
rect 27916 21532 28196 21534
rect 28364 21924 28420 22316
rect 28700 22370 28756 25228
rect 28812 23044 28868 33964
rect 28924 28084 28980 28094
rect 29036 28084 29092 35308
rect 29260 33570 29316 35532
rect 29372 35364 29428 36204
rect 29484 35924 29540 35934
rect 29484 35700 29540 35868
rect 29484 35606 29540 35644
rect 29596 35476 29652 36988
rect 30192 36876 30456 36886
rect 30248 36820 30296 36876
rect 30352 36820 30400 36876
rect 30192 36810 30456 36820
rect 31164 36596 31220 36606
rect 31164 36502 31220 36540
rect 31612 36596 31668 37212
rect 33852 36708 33908 37212
rect 33852 36652 34916 36708
rect 31612 36502 31668 36540
rect 32844 36596 32900 36606
rect 30716 36482 30772 36494
rect 30716 36430 30718 36482
rect 30770 36430 30772 36482
rect 29820 36372 29876 36382
rect 29820 36278 29876 36316
rect 30380 36370 30436 36382
rect 30380 36318 30382 36370
rect 30434 36318 30436 36370
rect 30380 35922 30436 36318
rect 30380 35870 30382 35922
rect 30434 35870 30436 35922
rect 30380 35858 30436 35870
rect 30492 36258 30548 36270
rect 30492 36206 30494 36258
rect 30546 36206 30548 36258
rect 30156 35698 30212 35710
rect 30156 35646 30158 35698
rect 30210 35646 30212 35698
rect 30156 35588 30212 35646
rect 30492 35700 30548 36206
rect 30492 35644 30660 35700
rect 30156 35522 30212 35532
rect 29596 35410 29652 35420
rect 29708 35476 29764 35486
rect 30492 35476 30548 35514
rect 29708 35474 29876 35476
rect 29708 35422 29710 35474
rect 29762 35422 29876 35474
rect 29708 35420 29876 35422
rect 29708 35410 29764 35420
rect 29372 35298 29428 35308
rect 29484 34916 29540 34926
rect 29484 34822 29540 34860
rect 29708 34804 29764 34814
rect 29708 34710 29764 34748
rect 29596 34690 29652 34702
rect 29596 34638 29598 34690
rect 29650 34638 29652 34690
rect 29372 34354 29428 34366
rect 29372 34302 29374 34354
rect 29426 34302 29428 34354
rect 29372 33908 29428 34302
rect 29484 34132 29540 34142
rect 29596 34132 29652 34638
rect 29820 34580 29876 35420
rect 30492 35410 30548 35420
rect 30192 35308 30456 35318
rect 30248 35252 30296 35308
rect 30352 35252 30400 35308
rect 30192 35242 30456 35252
rect 29820 34468 29876 34524
rect 30044 34914 30100 34926
rect 30044 34862 30046 34914
rect 30098 34862 30100 34914
rect 29820 34412 29988 34468
rect 29932 34244 29988 34412
rect 30044 34356 30100 34862
rect 30604 34916 30660 35644
rect 30604 34850 30660 34860
rect 30716 34580 30772 36430
rect 32844 36482 32900 36540
rect 32844 36430 32846 36482
rect 32898 36430 32900 36482
rect 32844 36418 32900 36430
rect 33852 36482 33908 36652
rect 34860 36594 34916 36652
rect 34860 36542 34862 36594
rect 34914 36542 34916 36594
rect 34860 36530 34916 36542
rect 33852 36430 33854 36482
rect 33906 36430 33908 36482
rect 33852 36418 33908 36430
rect 34412 36482 34468 36494
rect 34412 36430 34414 36482
rect 34466 36430 34468 36482
rect 32508 36370 32564 36382
rect 32508 36318 32510 36370
rect 32562 36318 32564 36370
rect 32172 36258 32228 36270
rect 32172 36206 32174 36258
rect 32226 36206 32228 36258
rect 31276 35700 31332 35710
rect 31276 35606 31332 35644
rect 30828 35586 30884 35598
rect 30828 35534 30830 35586
rect 30882 35534 30884 35586
rect 30828 34916 30884 35534
rect 31948 35588 32004 35598
rect 31164 34916 31220 34926
rect 31948 34916 32004 35532
rect 30828 34914 31108 34916
rect 30828 34862 30830 34914
rect 30882 34862 31108 34914
rect 30828 34860 31108 34862
rect 30828 34804 30884 34860
rect 30828 34738 30884 34748
rect 30716 34514 30772 34524
rect 30044 34290 30100 34300
rect 29932 34178 29988 34188
rect 29484 34130 29652 34132
rect 29484 34078 29486 34130
rect 29538 34078 29652 34130
rect 29484 34076 29652 34078
rect 29820 34130 29876 34142
rect 29820 34078 29822 34130
rect 29874 34078 29876 34130
rect 29484 34066 29540 34076
rect 29708 34018 29764 34030
rect 29708 33966 29710 34018
rect 29762 33966 29764 34018
rect 29708 33908 29764 33966
rect 29372 33852 29764 33908
rect 29820 33572 29876 34078
rect 29260 33518 29262 33570
rect 29314 33518 29316 33570
rect 29260 33506 29316 33518
rect 29372 33516 29876 33572
rect 29932 34018 29988 34030
rect 29932 33966 29934 34018
rect 29986 33966 29988 34018
rect 29372 33346 29428 33516
rect 29372 33294 29374 33346
rect 29426 33294 29428 33346
rect 29372 33282 29428 33294
rect 29260 33236 29316 33246
rect 29260 33142 29316 33180
rect 29484 32004 29540 32014
rect 29708 32004 29764 33516
rect 29820 33124 29876 33134
rect 29820 33030 29876 33068
rect 29932 32562 29988 33966
rect 30192 33740 30456 33750
rect 30248 33684 30296 33740
rect 30352 33684 30400 33740
rect 30192 33674 30456 33684
rect 30380 33348 30436 33358
rect 29932 32510 29934 32562
rect 29986 32510 29988 32562
rect 29932 32498 29988 32510
rect 30044 33234 30100 33246
rect 30044 33182 30046 33234
rect 30098 33182 30100 33234
rect 29820 32004 29876 32014
rect 29708 32002 29876 32004
rect 29708 31950 29822 32002
rect 29874 31950 29876 32002
rect 29708 31948 29876 31950
rect 30044 32004 30100 33182
rect 30380 32340 30436 33292
rect 30828 32564 30884 32574
rect 30828 32470 30884 32508
rect 30716 32450 30772 32462
rect 30716 32398 30718 32450
rect 30770 32398 30772 32450
rect 30380 32284 30660 32340
rect 30192 32172 30456 32182
rect 30248 32116 30296 32172
rect 30352 32116 30400 32172
rect 30192 32106 30456 32116
rect 30604 32004 30660 32284
rect 30044 31948 30324 32004
rect 29484 31890 29540 31948
rect 29820 31938 29876 31948
rect 29484 31838 29486 31890
rect 29538 31838 29540 31890
rect 29484 31826 29540 31838
rect 30156 31780 30212 31790
rect 30156 31686 30212 31724
rect 30268 31668 30324 31948
rect 30604 31938 30660 31948
rect 30380 31668 30436 31678
rect 30268 31612 30380 31668
rect 30380 31574 30436 31612
rect 29596 31556 29652 31566
rect 29596 30660 29652 31500
rect 30492 31556 30548 31566
rect 30156 31108 30212 31118
rect 30044 31052 30156 31108
rect 29484 30604 29652 30660
rect 29932 30994 29988 31006
rect 29932 30942 29934 30994
rect 29986 30942 29988 30994
rect 28980 28028 29092 28084
rect 29148 30212 29204 30222
rect 28924 28018 28980 28028
rect 29036 27860 29092 27870
rect 29036 27766 29092 27804
rect 28924 26290 28980 26302
rect 28924 26238 28926 26290
rect 28978 26238 28980 26290
rect 28924 25284 28980 26238
rect 28924 25218 28980 25228
rect 29036 25282 29092 25294
rect 29036 25230 29038 25282
rect 29090 25230 29092 25282
rect 28924 25060 28980 25070
rect 28924 24946 28980 25004
rect 28924 24894 28926 24946
rect 28978 24894 28980 24946
rect 28924 24882 28980 24894
rect 29036 24948 29092 25230
rect 29036 24882 29092 24892
rect 29036 24724 29092 24734
rect 28924 24500 28980 24510
rect 28924 24406 28980 24444
rect 28812 22978 28868 22988
rect 29036 22932 29092 24668
rect 29148 23042 29204 30156
rect 29372 30212 29428 30222
rect 29260 29988 29316 29998
rect 29260 29894 29316 29932
rect 29372 29652 29428 30156
rect 29372 29586 29428 29596
rect 29484 29428 29540 30604
rect 29596 30324 29652 30334
rect 29596 30210 29652 30268
rect 29932 30212 29988 30942
rect 30044 30436 30100 31052
rect 30156 31014 30212 31052
rect 30492 30994 30548 31500
rect 30492 30942 30494 30994
rect 30546 30942 30548 30994
rect 30492 30930 30548 30942
rect 30716 30660 30772 32398
rect 30940 31666 30996 31678
rect 30940 31614 30942 31666
rect 30994 31614 30996 31666
rect 30940 31444 30996 31614
rect 31052 31556 31108 34860
rect 31164 34914 32004 34916
rect 31164 34862 31166 34914
rect 31218 34862 32004 34914
rect 31164 34860 32004 34862
rect 31164 34850 31220 34860
rect 31164 33236 31220 33246
rect 31164 33142 31220 33180
rect 31276 31778 31332 34860
rect 31500 34580 31556 34590
rect 31500 34132 31556 34524
rect 31948 34356 32004 34860
rect 31948 34290 32004 34300
rect 32172 35476 32228 36206
rect 31500 33570 31556 34076
rect 32060 34132 32116 34142
rect 32060 34038 32116 34076
rect 31948 34020 32004 34030
rect 31948 33926 32004 33964
rect 31500 33518 31502 33570
rect 31554 33518 31556 33570
rect 31500 33506 31556 33518
rect 31388 33460 31444 33470
rect 31388 32116 31444 33404
rect 31836 33460 31892 33470
rect 31836 33234 31892 33404
rect 31836 33182 31838 33234
rect 31890 33182 31892 33234
rect 31836 33170 31892 33182
rect 32060 33236 32116 33246
rect 32060 33142 32116 33180
rect 31388 32050 31444 32060
rect 31836 32562 31892 32574
rect 31836 32510 31838 32562
rect 31890 32510 31892 32562
rect 31836 32452 31892 32510
rect 31836 32004 31892 32396
rect 31836 31938 31892 31948
rect 31388 31892 31444 31902
rect 31388 31798 31444 31836
rect 31276 31726 31278 31778
rect 31330 31726 31332 31778
rect 31276 31714 31332 31726
rect 31500 31780 31556 31790
rect 31836 31780 31892 31790
rect 31500 31686 31556 31724
rect 31612 31778 31892 31780
rect 31612 31726 31838 31778
rect 31890 31726 31892 31778
rect 31612 31724 31892 31726
rect 31052 31490 31108 31500
rect 31388 31668 31444 31678
rect 30940 31378 30996 31388
rect 31276 31332 31332 31342
rect 30192 30604 30456 30614
rect 30248 30548 30296 30604
rect 30352 30548 30400 30604
rect 30192 30538 30456 30548
rect 30044 30380 30212 30436
rect 29596 30158 29598 30210
rect 29650 30158 29652 30210
rect 29596 30146 29652 30158
rect 29820 30156 29932 30212
rect 29708 30100 29764 30110
rect 29708 30006 29764 30044
rect 29708 29540 29764 29550
rect 29596 29428 29652 29438
rect 29484 29426 29652 29428
rect 29484 29374 29598 29426
rect 29650 29374 29652 29426
rect 29484 29372 29652 29374
rect 29596 29362 29652 29372
rect 29708 26628 29764 29484
rect 29820 28868 29876 30156
rect 29932 30146 29988 30156
rect 29932 29652 29988 29662
rect 29932 29558 29988 29596
rect 30156 29652 30212 30380
rect 30716 29988 30772 30604
rect 30156 29558 30212 29596
rect 30604 29932 30772 29988
rect 30828 31106 30884 31118
rect 30828 31054 30830 31106
rect 30882 31054 30884 31106
rect 30044 29540 30100 29550
rect 30044 29314 30100 29484
rect 30044 29262 30046 29314
rect 30098 29262 30100 29314
rect 30044 29250 30100 29262
rect 30192 29036 30456 29046
rect 30248 28980 30296 29036
rect 30352 28980 30400 29036
rect 30192 28970 30456 28980
rect 30380 28868 30436 28878
rect 29820 28812 30212 28868
rect 30156 28756 30212 28812
rect 30268 28756 30324 28766
rect 30156 28754 30324 28756
rect 30156 28702 30270 28754
rect 30322 28702 30324 28754
rect 30156 28700 30324 28702
rect 30268 28690 30324 28700
rect 29820 28642 29876 28654
rect 29820 28590 29822 28642
rect 29874 28590 29876 28642
rect 29820 27076 29876 28590
rect 30044 28642 30100 28654
rect 30044 28590 30046 28642
rect 30098 28590 30100 28642
rect 30044 27300 30100 28590
rect 30380 27858 30436 28812
rect 30380 27806 30382 27858
rect 30434 27806 30436 27858
rect 30380 27794 30436 27806
rect 30492 27860 30548 27898
rect 30492 27794 30548 27804
rect 30492 27636 30548 27646
rect 30604 27636 30660 29932
rect 30828 29764 30884 31054
rect 30828 29426 30884 29708
rect 31164 29986 31220 29998
rect 31164 29934 31166 29986
rect 31218 29934 31220 29986
rect 30828 29374 30830 29426
rect 30882 29374 30884 29426
rect 30828 29362 30884 29374
rect 31052 29652 31108 29662
rect 31052 29426 31108 29596
rect 31052 29374 31054 29426
rect 31106 29374 31108 29426
rect 31052 29362 31108 29374
rect 31164 28642 31220 29934
rect 31276 28754 31332 31276
rect 31276 28702 31278 28754
rect 31330 28702 31332 28754
rect 31276 28690 31332 28702
rect 31164 28590 31166 28642
rect 31218 28590 31220 28642
rect 31164 28578 31220 28590
rect 30940 28532 30996 28542
rect 30940 28438 30996 28476
rect 31164 28308 31220 28318
rect 30716 27972 30772 27982
rect 30716 27858 30772 27916
rect 30716 27806 30718 27858
rect 30770 27806 30772 27858
rect 30716 27794 30772 27806
rect 30548 27580 30660 27636
rect 30828 27636 30884 27646
rect 30492 27570 30548 27580
rect 30828 27542 30884 27580
rect 30192 27468 30456 27478
rect 30248 27412 30296 27468
rect 30352 27412 30400 27468
rect 30192 27402 30456 27412
rect 30380 27300 30436 27310
rect 30044 27298 30436 27300
rect 30044 27246 30382 27298
rect 30434 27246 30436 27298
rect 30044 27244 30436 27246
rect 30380 27234 30436 27244
rect 31164 27300 31220 28252
rect 29820 27010 29876 27020
rect 30828 27074 30884 27086
rect 30828 27022 30830 27074
rect 30882 27022 30884 27074
rect 30380 26964 30436 27002
rect 30380 26898 30436 26908
rect 30492 26964 30548 26974
rect 30828 26964 30884 27022
rect 30492 26962 30884 26964
rect 30492 26910 30494 26962
rect 30546 26910 30884 26962
rect 30492 26908 30884 26910
rect 30492 26898 30548 26908
rect 29708 26562 29764 26572
rect 30716 26404 30772 26414
rect 29372 26292 29428 26302
rect 29372 26198 29428 26236
rect 29820 26178 29876 26190
rect 29820 26126 29822 26178
rect 29874 26126 29876 26178
rect 29260 25620 29316 25630
rect 29260 25394 29316 25564
rect 29260 25342 29262 25394
rect 29314 25342 29316 25394
rect 29260 25330 29316 25342
rect 29372 25394 29428 25406
rect 29372 25342 29374 25394
rect 29426 25342 29428 25394
rect 29372 24724 29428 25342
rect 29596 25396 29652 25406
rect 29596 24948 29652 25340
rect 29820 25396 29876 26126
rect 30716 26178 30772 26348
rect 30716 26126 30718 26178
rect 30770 26126 30772 26178
rect 30192 25900 30456 25910
rect 30248 25844 30296 25900
rect 30352 25844 30400 25900
rect 30192 25834 30456 25844
rect 30268 25620 30324 25630
rect 30268 25526 30324 25564
rect 29820 25330 29876 25340
rect 29596 24882 29652 24892
rect 29708 25284 29764 25294
rect 29708 24946 29764 25228
rect 29932 25282 29988 25294
rect 29932 25230 29934 25282
rect 29986 25230 29988 25282
rect 29932 25060 29988 25230
rect 29932 24994 29988 25004
rect 30156 25284 30212 25294
rect 29708 24894 29710 24946
rect 29762 24894 29764 24946
rect 29708 24882 29764 24894
rect 30044 24948 30100 24958
rect 29372 24658 29428 24668
rect 29820 24052 29876 24062
rect 29708 23940 29764 23978
rect 29820 23958 29876 23996
rect 29708 23874 29764 23884
rect 29484 23828 29540 23838
rect 29484 23826 29652 23828
rect 29484 23774 29486 23826
rect 29538 23774 29652 23826
rect 29484 23772 29652 23774
rect 29484 23762 29540 23772
rect 29148 22990 29150 23042
rect 29202 22990 29204 23042
rect 29148 22978 29204 22990
rect 29260 23268 29316 23278
rect 29036 22866 29092 22876
rect 28700 22318 28702 22370
rect 28754 22318 28756 22370
rect 28700 22306 28756 22318
rect 29148 22820 29204 22830
rect 29148 22370 29204 22764
rect 29148 22318 29150 22370
rect 29202 22318 29204 22370
rect 27916 21522 27972 21532
rect 27692 21308 27972 21364
rect 27132 20914 27524 20916
rect 27132 20862 27134 20914
rect 27186 20862 27524 20914
rect 27132 20860 27524 20862
rect 27132 20850 27188 20860
rect 27468 20804 27524 20860
rect 27468 20802 27748 20804
rect 27468 20750 27470 20802
rect 27522 20750 27748 20802
rect 27468 20748 27748 20750
rect 27468 20738 27524 20748
rect 27356 20580 27412 20590
rect 27412 20524 27524 20580
rect 27356 20514 27412 20524
rect 27468 20244 27524 20524
rect 27468 20188 27636 20244
rect 27132 20020 27188 20030
rect 27132 19926 27188 19964
rect 27468 20020 27524 20030
rect 27244 19796 27300 19806
rect 26572 19628 26852 19684
rect 27020 19628 27188 19684
rect 26796 19572 26852 19628
rect 26796 19516 27076 19572
rect 26236 19460 26292 19470
rect 26124 19236 26180 19246
rect 26124 19142 26180 19180
rect 25676 19012 25732 19022
rect 25676 17892 25732 18956
rect 26124 18676 26180 18686
rect 25676 17826 25732 17836
rect 26012 18562 26068 18574
rect 26012 18510 26014 18562
rect 26066 18510 26068 18562
rect 25564 17444 25620 17454
rect 25564 16658 25620 17388
rect 25564 16606 25566 16658
rect 25618 16606 25620 16658
rect 25564 16594 25620 16606
rect 25676 17220 25732 17230
rect 25564 16436 25620 16446
rect 25564 15314 25620 16380
rect 25564 15262 25566 15314
rect 25618 15262 25620 15314
rect 25564 15250 25620 15262
rect 25676 15316 25732 17164
rect 25788 16996 25844 17006
rect 26012 16996 26068 18510
rect 25844 16940 26068 16996
rect 25788 16902 25844 16940
rect 25788 16658 25844 16670
rect 25788 16606 25790 16658
rect 25842 16606 25844 16658
rect 25788 15988 25844 16606
rect 25788 15922 25844 15932
rect 25788 15316 25844 15326
rect 25676 15260 25788 15316
rect 25788 15222 25844 15260
rect 26012 15090 26068 15102
rect 26012 15038 26014 15090
rect 26066 15038 26068 15090
rect 25452 14252 25732 14308
rect 25452 13972 25508 13982
rect 25452 13970 25620 13972
rect 25452 13918 25454 13970
rect 25506 13918 25620 13970
rect 25452 13916 25620 13918
rect 25452 13906 25508 13916
rect 25564 13860 25620 13916
rect 25564 13794 25620 13804
rect 25004 13234 25060 13244
rect 25228 13748 25284 13758
rect 24892 12962 24948 13020
rect 25116 13076 25172 13114
rect 25116 13010 25172 13020
rect 24892 12910 24894 12962
rect 24946 12910 24948 12962
rect 24892 12898 24948 12910
rect 25228 12964 25284 13692
rect 25452 13748 25508 13758
rect 25340 13636 25396 13646
rect 25340 13542 25396 13580
rect 25452 13412 25508 13692
rect 25452 13346 25508 13356
rect 25228 12870 25284 12908
rect 25340 13300 25396 13310
rect 24668 12850 24836 12852
rect 24668 12798 24670 12850
rect 24722 12798 24836 12850
rect 24668 12796 24836 12798
rect 24668 12786 24724 12796
rect 23996 12238 23998 12290
rect 24050 12238 24052 12290
rect 23436 10500 23492 11340
rect 23548 11394 23604 11406
rect 23548 11342 23550 11394
rect 23602 11342 23604 11394
rect 23548 10948 23604 11342
rect 23772 11394 23828 11406
rect 23772 11342 23774 11394
rect 23826 11342 23828 11394
rect 23548 10882 23604 10892
rect 23660 11284 23716 11294
rect 23660 10724 23716 11228
rect 23660 10658 23716 10668
rect 23660 10500 23716 10510
rect 23436 10498 23716 10500
rect 23436 10446 23662 10498
rect 23714 10446 23716 10498
rect 23436 10444 23716 10446
rect 23660 10434 23716 10444
rect 23772 10276 23828 11342
rect 23996 11396 24052 12238
rect 24108 12740 24164 12750
rect 24108 11956 24164 12684
rect 24444 12740 24500 12750
rect 25340 12740 25396 13244
rect 24108 11890 24164 11900
rect 24220 12178 24276 12190
rect 24220 12126 24222 12178
rect 24274 12126 24276 12178
rect 24220 11732 24276 12126
rect 24332 12180 24388 12190
rect 24332 12086 24388 12124
rect 24444 12178 24500 12684
rect 25116 12684 25396 12740
rect 25452 12740 25508 12750
rect 24780 12628 24836 12638
rect 24444 12126 24446 12178
rect 24498 12126 24500 12178
rect 24444 11788 24500 12126
rect 24668 12516 24724 12526
rect 24668 12178 24724 12460
rect 24668 12126 24670 12178
rect 24722 12126 24724 12178
rect 24668 12114 24724 12126
rect 24220 11666 24276 11676
rect 24332 11732 24500 11788
rect 23996 11330 24052 11340
rect 24108 11284 24164 11294
rect 24108 11190 24164 11228
rect 23996 11170 24052 11182
rect 23996 11118 23998 11170
rect 24050 11118 24052 11170
rect 23996 10948 24052 11118
rect 23996 10882 24052 10892
rect 24220 11172 24276 11182
rect 24332 11172 24388 11732
rect 24444 11620 24500 11630
rect 24444 11394 24500 11564
rect 24444 11342 24446 11394
rect 24498 11342 24500 11394
rect 24444 11330 24500 11342
rect 24556 11284 24612 11294
rect 24556 11190 24612 11228
rect 24332 11116 24500 11172
rect 24220 10666 24276 11116
rect 23884 10610 23940 10622
rect 23884 10558 23886 10610
rect 23938 10558 23940 10610
rect 23884 10388 23940 10558
rect 24108 10612 24164 10650
rect 24220 10614 24222 10666
rect 24274 10614 24276 10666
rect 24220 10602 24276 10614
rect 24444 10612 24500 11116
rect 24668 11170 24724 11182
rect 24668 11118 24670 11170
rect 24722 11118 24724 11170
rect 24668 11060 24724 11118
rect 24556 11004 24724 11060
rect 24556 10836 24612 11004
rect 24556 10770 24612 10780
rect 24668 10836 24724 10846
rect 24780 10836 24836 12572
rect 25116 11508 25172 12684
rect 25452 12646 25508 12684
rect 25676 12516 25732 14252
rect 25900 14196 25956 14206
rect 25228 12460 25732 12516
rect 25788 13972 25844 13982
rect 25228 12402 25284 12460
rect 25228 12350 25230 12402
rect 25282 12350 25284 12402
rect 25228 12338 25284 12350
rect 25788 12404 25844 13916
rect 25900 12516 25956 14140
rect 26012 13860 26068 15038
rect 26012 13794 26068 13804
rect 26012 13634 26068 13646
rect 26012 13582 26014 13634
rect 26066 13582 26068 13634
rect 26012 13300 26068 13582
rect 26124 13636 26180 18620
rect 26236 14868 26292 19404
rect 27020 19460 27076 19516
rect 27020 19346 27076 19404
rect 27020 19294 27022 19346
rect 27074 19294 27076 19346
rect 27020 19282 27076 19294
rect 26572 19236 26628 19246
rect 26572 19142 26628 19180
rect 27132 19236 27188 19628
rect 27132 19170 27188 19180
rect 27244 19012 27300 19740
rect 27468 19458 27524 19964
rect 27468 19406 27470 19458
rect 27522 19406 27524 19458
rect 27468 19394 27524 19406
rect 27356 19236 27412 19246
rect 27356 19142 27412 19180
rect 27132 18956 27300 19012
rect 27132 18564 27188 18956
rect 27020 18508 27188 18564
rect 27244 18788 27300 18798
rect 27580 18788 27636 20188
rect 27692 19236 27748 20748
rect 27916 20132 27972 21308
rect 28252 20914 28308 20926
rect 28252 20862 28254 20914
rect 28306 20862 28308 20914
rect 28140 20692 28196 20702
rect 28140 20132 28196 20636
rect 27916 20066 27972 20076
rect 28028 20076 28196 20132
rect 27804 20020 27860 20030
rect 27804 19926 27860 19964
rect 27804 19236 27860 19246
rect 27692 19234 27860 19236
rect 27692 19182 27806 19234
rect 27858 19182 27860 19234
rect 27692 19180 27860 19182
rect 27804 19170 27860 19180
rect 27916 19236 27972 19246
rect 27916 19122 27972 19180
rect 27916 19070 27918 19122
rect 27970 19070 27972 19122
rect 27916 19058 27972 19070
rect 28028 19124 28084 20076
rect 28140 19908 28196 19918
rect 28140 19234 28196 19852
rect 28140 19182 28142 19234
rect 28194 19182 28196 19234
rect 28140 19170 28196 19182
rect 28028 19058 28084 19068
rect 28028 18900 28084 18910
rect 27580 18732 27972 18788
rect 26348 18452 26404 18462
rect 26348 18450 26628 18452
rect 26348 18398 26350 18450
rect 26402 18398 26628 18450
rect 26348 18396 26628 18398
rect 26348 18386 26404 18396
rect 26572 18226 26628 18396
rect 26572 18174 26574 18226
rect 26626 18174 26628 18226
rect 26572 18162 26628 18174
rect 26908 18338 26964 18350
rect 26908 18286 26910 18338
rect 26962 18286 26964 18338
rect 26908 18226 26964 18286
rect 26908 18174 26910 18226
rect 26962 18174 26964 18226
rect 26908 18162 26964 18174
rect 26796 17556 26852 17566
rect 26796 17462 26852 17500
rect 26684 16884 26740 16894
rect 27020 16884 27076 18508
rect 27132 17442 27188 17454
rect 27132 17390 27134 17442
rect 27186 17390 27188 17442
rect 27132 17108 27188 17390
rect 27132 17042 27188 17052
rect 27244 17108 27300 18732
rect 27692 18450 27748 18462
rect 27692 18398 27694 18450
rect 27746 18398 27748 18450
rect 27356 18340 27412 18350
rect 27692 18340 27748 18398
rect 27356 18338 27748 18340
rect 27356 18286 27358 18338
rect 27410 18286 27748 18338
rect 27356 18284 27748 18286
rect 27356 18226 27412 18284
rect 27356 18174 27358 18226
rect 27410 18174 27412 18226
rect 27356 18162 27412 18174
rect 27692 18228 27748 18284
rect 27692 18162 27748 18172
rect 27916 17554 27972 18732
rect 28028 18338 28084 18844
rect 28252 18452 28308 20862
rect 28364 20802 28420 21868
rect 29036 21586 29092 21598
rect 29036 21534 29038 21586
rect 29090 21534 29092 21586
rect 28588 21476 28644 21486
rect 28588 21382 28644 21420
rect 28364 20750 28366 20802
rect 28418 20750 28420 20802
rect 28364 20738 28420 20750
rect 28700 20468 28756 20478
rect 28364 20132 28420 20142
rect 28364 20130 28644 20132
rect 28364 20078 28366 20130
rect 28418 20078 28644 20130
rect 28364 20076 28644 20078
rect 28364 20066 28420 20076
rect 28588 19460 28644 20076
rect 28588 19346 28644 19404
rect 28588 19294 28590 19346
rect 28642 19294 28644 19346
rect 28588 19236 28644 19294
rect 28588 19170 28644 19180
rect 28700 19012 28756 20412
rect 29036 19908 29092 21534
rect 29148 21476 29204 22318
rect 29260 21586 29316 23212
rect 29596 23154 29652 23772
rect 29596 23102 29598 23154
rect 29650 23102 29652 23154
rect 29596 22370 29652 23102
rect 29596 22318 29598 22370
rect 29650 22318 29652 22370
rect 29596 22148 29652 22318
rect 29932 22258 29988 22270
rect 29932 22206 29934 22258
rect 29986 22206 29988 22258
rect 29932 22148 29988 22206
rect 29596 22092 29764 22148
rect 29596 21812 29652 21822
rect 29260 21534 29262 21586
rect 29314 21534 29316 21586
rect 29260 21522 29316 21534
rect 29372 21588 29428 21598
rect 29148 20580 29204 21420
rect 29372 20804 29428 21532
rect 29596 21588 29652 21756
rect 29596 21522 29652 21532
rect 29596 21364 29652 21374
rect 29708 21364 29764 22092
rect 29932 22082 29988 22092
rect 29932 21812 29988 21822
rect 29932 21718 29988 21756
rect 29652 21308 29764 21364
rect 29820 21698 29876 21710
rect 29820 21646 29822 21698
rect 29874 21646 29876 21698
rect 29820 21588 29876 21646
rect 29484 20804 29540 20814
rect 29372 20802 29540 20804
rect 29372 20750 29486 20802
rect 29538 20750 29540 20802
rect 29372 20748 29540 20750
rect 29484 20738 29540 20748
rect 29260 20580 29316 20590
rect 29148 20524 29260 20580
rect 29260 20514 29316 20524
rect 29036 19842 29092 19852
rect 29372 20020 29428 20030
rect 29036 19236 29092 19246
rect 29036 19142 29092 19180
rect 29372 19234 29428 19964
rect 29596 20018 29652 21308
rect 29820 21028 29876 21532
rect 29708 20972 29876 21028
rect 29708 20468 29764 20972
rect 29820 20804 29876 20814
rect 29820 20690 29876 20748
rect 29820 20638 29822 20690
rect 29874 20638 29876 20690
rect 29820 20626 29876 20638
rect 29708 20402 29764 20412
rect 29596 19966 29598 20018
rect 29650 19966 29652 20018
rect 29596 19954 29652 19966
rect 29820 20244 29876 20254
rect 29372 19182 29374 19234
rect 29426 19182 29428 19234
rect 29372 19170 29428 19182
rect 29708 19236 29764 19246
rect 29708 19142 29764 19180
rect 29596 19012 29652 19022
rect 28700 19010 29652 19012
rect 28700 18958 29598 19010
rect 29650 18958 29652 19010
rect 28700 18956 29652 18958
rect 28700 18674 28756 18956
rect 29596 18946 29652 18956
rect 29708 19012 29764 19022
rect 28700 18622 28702 18674
rect 28754 18622 28756 18674
rect 28700 18610 28756 18622
rect 28252 18386 28308 18396
rect 29036 18452 29092 18462
rect 29092 18396 29316 18452
rect 29036 18358 29092 18396
rect 28028 18286 28030 18338
rect 28082 18286 28084 18338
rect 28028 18274 28084 18286
rect 27916 17502 27918 17554
rect 27970 17502 27972 17554
rect 27916 17490 27972 17502
rect 29260 17666 29316 18396
rect 29484 18340 29540 18350
rect 29484 18116 29540 18284
rect 29484 18050 29540 18060
rect 29260 17614 29262 17666
rect 29314 17614 29316 17666
rect 27692 17442 27748 17454
rect 27692 17390 27694 17442
rect 27746 17390 27748 17442
rect 27580 17108 27636 17118
rect 27244 17106 27636 17108
rect 27244 17054 27246 17106
rect 27298 17054 27582 17106
rect 27634 17054 27636 17106
rect 27244 17052 27636 17054
rect 27244 17042 27300 17052
rect 27580 17042 27636 17052
rect 27692 16996 27748 17390
rect 28252 17442 28308 17454
rect 28252 17390 28254 17442
rect 28306 17390 28308 17442
rect 27692 16930 27748 16940
rect 27804 17332 27860 17342
rect 27020 16828 27188 16884
rect 26684 16790 26740 16828
rect 26348 16212 26404 16222
rect 26348 15652 26404 16156
rect 26460 16100 26516 16110
rect 26460 16098 26628 16100
rect 26460 16046 26462 16098
rect 26514 16046 26628 16098
rect 26460 16044 26628 16046
rect 26460 16034 26516 16044
rect 26348 15596 26516 15652
rect 26348 15314 26404 15326
rect 26348 15262 26350 15314
rect 26402 15262 26404 15314
rect 26348 15092 26404 15262
rect 26460 15314 26516 15596
rect 26460 15262 26462 15314
rect 26514 15262 26516 15314
rect 26460 15250 26516 15262
rect 26348 15026 26404 15036
rect 26236 14812 26404 14868
rect 26124 13570 26180 13580
rect 26236 13748 26292 13758
rect 26012 12628 26068 13244
rect 26236 13076 26292 13692
rect 26124 12964 26180 12974
rect 26236 12964 26292 13020
rect 26124 12962 26292 12964
rect 26124 12910 26126 12962
rect 26178 12910 26292 12962
rect 26124 12908 26292 12910
rect 26124 12898 26180 12908
rect 26348 12628 26404 14812
rect 26572 14084 26628 16044
rect 27020 15988 27076 15998
rect 27020 15894 27076 15932
rect 27132 15876 27188 16828
rect 27468 15988 27524 15998
rect 27468 15894 27524 15932
rect 27132 15820 27300 15876
rect 26460 14028 26628 14084
rect 26684 15538 26740 15550
rect 26684 15486 26686 15538
rect 26738 15486 26740 15538
rect 26684 14084 26740 15486
rect 27132 15316 27188 15326
rect 27132 15202 27188 15260
rect 27132 15150 27134 15202
rect 27186 15150 27188 15202
rect 26908 14754 26964 14766
rect 26908 14702 26910 14754
rect 26962 14702 26964 14754
rect 26908 14642 26964 14702
rect 26908 14590 26910 14642
rect 26962 14590 26964 14642
rect 26908 14578 26964 14590
rect 27132 14308 27188 15150
rect 27132 14242 27188 14252
rect 26684 14028 27188 14084
rect 26460 13860 26516 14028
rect 26460 13804 26628 13860
rect 26460 13636 26516 13646
rect 26460 13300 26516 13580
rect 26572 13412 26628 13804
rect 27132 13746 27188 14028
rect 27132 13694 27134 13746
rect 27186 13694 27188 13746
rect 27132 13682 27188 13694
rect 26684 13636 26740 13646
rect 26684 13542 26740 13580
rect 26908 13524 26964 13534
rect 26908 13430 26964 13468
rect 26572 13356 26740 13412
rect 26460 13244 26628 13300
rect 26460 13076 26516 13086
rect 26460 12962 26516 13020
rect 26460 12910 26462 12962
rect 26514 12910 26516 12962
rect 26460 12898 26516 12910
rect 26572 12740 26628 13244
rect 26012 12572 26180 12628
rect 25900 12460 26068 12516
rect 25788 12348 25956 12404
rect 25676 12180 25732 12190
rect 25676 12086 25732 12124
rect 25788 12178 25844 12190
rect 25788 12126 25790 12178
rect 25842 12126 25844 12178
rect 25452 12068 25508 12078
rect 25340 11620 25396 11630
rect 25004 11452 25172 11508
rect 25228 11564 25340 11620
rect 24668 10834 24836 10836
rect 24668 10782 24670 10834
rect 24722 10782 24836 10834
rect 24668 10780 24836 10782
rect 24892 11396 24948 11406
rect 24668 10770 24724 10780
rect 24892 10612 24948 11340
rect 24444 10556 24612 10612
rect 24108 10546 24164 10556
rect 23996 10388 24052 10398
rect 23884 10332 23996 10388
rect 23996 10322 24052 10332
rect 23772 10210 23828 10220
rect 23324 10098 23380 10108
rect 24108 10164 24164 10174
rect 24556 10108 24612 10556
rect 23324 9044 23380 9054
rect 23324 9042 23492 9044
rect 23324 8990 23326 9042
rect 23378 8990 23492 9042
rect 23324 8988 23492 8990
rect 23324 8978 23380 8988
rect 23436 7698 23492 8988
rect 23884 8148 23940 8158
rect 23436 7646 23438 7698
rect 23490 7646 23492 7698
rect 23436 7634 23492 7646
rect 23772 8092 23884 8148
rect 23772 7474 23828 8092
rect 23884 8082 23940 8092
rect 24108 7812 24164 10108
rect 24332 10052 24612 10108
rect 24668 10556 24948 10612
rect 24332 7812 24388 10052
rect 24668 8484 24724 10556
rect 25004 10500 25060 11452
rect 24780 10444 25060 10500
rect 25116 11282 25172 11294
rect 25116 11230 25118 11282
rect 25170 11230 25172 11282
rect 24780 8596 24836 10444
rect 24892 10164 24948 10174
rect 24892 9938 24948 10108
rect 25116 10052 25172 11230
rect 25116 9986 25172 9996
rect 24892 9886 24894 9938
rect 24946 9886 24948 9938
rect 24892 9874 24948 9886
rect 25228 9940 25284 11564
rect 25340 11554 25396 11564
rect 25340 11396 25396 11406
rect 25452 11396 25508 12012
rect 25676 11956 25732 11966
rect 25340 11394 25508 11396
rect 25340 11342 25342 11394
rect 25394 11342 25508 11394
rect 25340 11340 25508 11342
rect 25564 11508 25620 11518
rect 25564 11394 25620 11452
rect 25564 11342 25566 11394
rect 25618 11342 25620 11394
rect 25340 11330 25396 11340
rect 25452 11172 25508 11182
rect 25340 11170 25508 11172
rect 25340 11118 25454 11170
rect 25506 11118 25508 11170
rect 25340 11116 25508 11118
rect 25340 10388 25396 11116
rect 25452 11106 25508 11116
rect 25452 10948 25508 10958
rect 25452 10834 25508 10892
rect 25452 10782 25454 10834
rect 25506 10782 25508 10834
rect 25452 10770 25508 10782
rect 25340 10322 25396 10332
rect 25564 10164 25620 11342
rect 25676 11394 25732 11900
rect 25788 11508 25844 12126
rect 25788 11442 25844 11452
rect 25676 11342 25678 11394
rect 25730 11342 25732 11394
rect 25676 11330 25732 11342
rect 25788 11284 25844 11294
rect 25788 10948 25844 11228
rect 25788 10882 25844 10892
rect 25564 10098 25620 10108
rect 25788 10276 25844 10286
rect 25340 9940 25396 9950
rect 25228 9938 25396 9940
rect 25228 9886 25342 9938
rect 25394 9886 25396 9938
rect 25228 9884 25396 9886
rect 25340 9874 25396 9884
rect 25788 9938 25844 10220
rect 25788 9886 25790 9938
rect 25842 9886 25844 9938
rect 25788 9874 25844 9886
rect 24780 8540 25172 8596
rect 24668 8428 24948 8484
rect 24668 8148 24724 8428
rect 24892 8370 24948 8428
rect 24892 8318 24894 8370
rect 24946 8318 24948 8370
rect 24892 8306 24948 8318
rect 24668 8082 24724 8092
rect 24108 7756 24276 7812
rect 24332 7756 24500 7812
rect 24220 7700 24276 7756
rect 23996 7588 24052 7598
rect 24220 7588 24276 7644
rect 24332 7588 24388 7598
rect 24220 7586 24388 7588
rect 24220 7534 24334 7586
rect 24386 7534 24388 7586
rect 24220 7532 24388 7534
rect 23996 7494 24052 7532
rect 24332 7522 24388 7532
rect 23772 7422 23774 7474
rect 23826 7422 23828 7474
rect 23772 7410 23828 7422
rect 23436 6018 23492 6030
rect 23436 5966 23438 6018
rect 23490 5966 23492 6018
rect 23212 5012 23268 5022
rect 23100 4956 23212 5012
rect 23436 5012 23492 5966
rect 23548 5906 23604 5918
rect 23548 5854 23550 5906
rect 23602 5854 23604 5906
rect 23548 5796 23604 5854
rect 23548 5730 23604 5740
rect 24220 5796 24276 5806
rect 24220 5702 24276 5740
rect 24332 5236 24388 5246
rect 24444 5236 24500 7756
rect 25004 7700 25060 7710
rect 25004 6802 25060 7644
rect 25004 6750 25006 6802
rect 25058 6750 25060 6802
rect 25004 6738 25060 6750
rect 25116 6132 25172 8540
rect 25340 8036 25396 8046
rect 25340 7700 25396 7980
rect 25900 7924 25956 12348
rect 26012 12178 26068 12460
rect 26124 12292 26180 12572
rect 26236 12572 26404 12628
rect 26460 12684 26628 12740
rect 26684 12962 26740 13356
rect 26684 12910 26686 12962
rect 26738 12910 26740 12962
rect 26236 12404 26292 12572
rect 26236 12348 26404 12404
rect 26124 12236 26292 12292
rect 26012 12126 26014 12178
rect 26066 12126 26068 12178
rect 26012 12114 26068 12126
rect 26236 12068 26292 12236
rect 26236 12002 26292 12012
rect 26124 11956 26180 11966
rect 26124 10834 26180 11900
rect 26348 11732 26404 12348
rect 26124 10782 26126 10834
rect 26178 10782 26180 10834
rect 26124 10770 26180 10782
rect 26236 11676 26404 11732
rect 26124 9042 26180 9054
rect 26124 8990 26126 9042
rect 26178 8990 26180 9042
rect 26124 8260 26180 8990
rect 26012 8036 26068 8046
rect 26012 7942 26068 7980
rect 25900 7858 25956 7868
rect 26124 7700 26180 8204
rect 25396 7644 25620 7700
rect 25340 7606 25396 7644
rect 25564 6690 25620 7644
rect 26124 7634 26180 7644
rect 25900 7588 25956 7598
rect 25900 7494 25956 7532
rect 25564 6638 25566 6690
rect 25618 6638 25620 6690
rect 25564 6626 25620 6638
rect 25340 6468 25396 6478
rect 25340 6374 25396 6412
rect 25116 6066 25172 6076
rect 25676 6132 25732 6142
rect 23660 5234 24500 5236
rect 23660 5182 24334 5234
rect 24386 5182 24500 5234
rect 23660 5180 24500 5182
rect 25004 5796 25060 5806
rect 23436 4956 23604 5012
rect 23212 4946 23268 4956
rect 23548 4676 23604 4956
rect 23548 4610 23604 4620
rect 23324 4564 23380 4574
rect 23324 4470 23380 4508
rect 23660 4338 23716 5180
rect 24332 5170 24388 5180
rect 24556 5012 24612 5022
rect 24444 4676 24500 4686
rect 23660 4286 23662 4338
rect 23714 4286 23716 4338
rect 23660 4274 23716 4286
rect 23884 4450 23940 4462
rect 23884 4398 23886 4450
rect 23938 4398 23940 4450
rect 23884 4340 23940 4398
rect 24444 4450 24500 4620
rect 24444 4398 24446 4450
rect 24498 4398 24500 4450
rect 24444 4386 24500 4398
rect 23884 4274 23940 4284
rect 22764 4174 22766 4226
rect 22818 4174 22820 4226
rect 22764 4162 22820 4174
rect 20972 3556 21028 3566
rect 20972 3462 21028 3500
rect 20748 3442 20916 3444
rect 20748 3390 20750 3442
rect 20802 3390 20916 3442
rect 20748 3388 20916 3390
rect 24108 3442 24164 3454
rect 24108 3390 24110 3442
rect 24162 3390 24164 3442
rect 20748 3378 20804 3388
rect 20532 3164 20796 3174
rect 20588 3108 20636 3164
rect 20692 3108 20740 3164
rect 20532 3098 20796 3108
rect 24108 3108 24164 3390
rect 24556 3330 24612 4956
rect 24556 3278 24558 3330
rect 24610 3278 24612 3330
rect 24556 3266 24612 3278
rect 24780 3554 24836 3566
rect 24780 3502 24782 3554
rect 24834 3502 24836 3554
rect 24780 3108 24836 3502
rect 24108 3052 24836 3108
rect 24108 2212 24164 3052
rect 25004 2548 25060 5740
rect 25676 5122 25732 6076
rect 26012 6132 26068 6142
rect 26012 6038 26068 6076
rect 26236 5572 26292 11676
rect 26348 11172 26404 11182
rect 26348 11078 26404 11116
rect 26460 9492 26516 12684
rect 26684 12292 26740 12910
rect 26572 12236 26740 12292
rect 26796 13188 26852 13198
rect 26796 12290 26852 13132
rect 27244 12850 27300 15820
rect 27356 15316 27412 15326
rect 27356 15148 27412 15260
rect 27580 15202 27636 15214
rect 27580 15150 27582 15202
rect 27634 15150 27636 15202
rect 27580 15148 27636 15150
rect 27356 15092 27636 15148
rect 27356 14754 27412 15092
rect 27356 14702 27358 14754
rect 27410 14702 27412 14754
rect 27356 13188 27412 14702
rect 27580 14308 27636 14318
rect 27356 13122 27412 13132
rect 27468 14306 27636 14308
rect 27468 14254 27582 14306
rect 27634 14254 27636 14306
rect 27468 14252 27636 14254
rect 27468 12964 27524 14252
rect 27580 14242 27636 14252
rect 27804 13860 27860 17276
rect 28028 17220 28084 17230
rect 28028 16770 28084 17164
rect 28252 16996 28308 17390
rect 28812 17108 28868 17118
rect 28812 17014 28868 17052
rect 28252 16930 28308 16940
rect 28476 16994 28532 17006
rect 28476 16942 28478 16994
rect 28530 16942 28532 16994
rect 28028 16718 28030 16770
rect 28082 16718 28084 16770
rect 28028 16706 28084 16718
rect 28476 16660 28532 16942
rect 29260 16884 29316 17614
rect 29260 16818 29316 16828
rect 29372 17780 29428 17790
rect 29708 17780 29764 18956
rect 28476 15876 28532 16604
rect 29372 16210 29428 17724
rect 29372 16158 29374 16210
rect 29426 16158 29428 16210
rect 29372 15876 29428 16158
rect 28476 15810 28532 15820
rect 28700 15820 29428 15876
rect 29484 17778 29764 17780
rect 29484 17726 29710 17778
rect 29762 17726 29764 17778
rect 29484 17724 29764 17726
rect 28140 15314 28196 15326
rect 28140 15262 28142 15314
rect 28194 15262 28196 15314
rect 28140 15204 28196 15262
rect 27916 15092 28196 15148
rect 28364 15316 28420 15326
rect 27916 14530 27972 15092
rect 27916 14478 27918 14530
rect 27970 14478 27972 14530
rect 27916 14466 27972 14478
rect 27804 13804 28196 13860
rect 27804 13636 27860 13646
rect 27804 13542 27860 13580
rect 27580 13522 27636 13534
rect 27580 13470 27582 13522
rect 27634 13470 27636 13522
rect 27580 13076 27636 13470
rect 27580 12982 27636 13020
rect 27468 12898 27524 12908
rect 27916 12962 27972 12974
rect 27916 12910 27918 12962
rect 27970 12910 27972 12962
rect 27244 12798 27246 12850
rect 27298 12798 27300 12850
rect 27244 12786 27300 12798
rect 26796 12238 26798 12290
rect 26850 12238 26852 12290
rect 26572 11844 26628 12236
rect 26796 12226 26852 12238
rect 26908 12738 26964 12750
rect 26908 12686 26910 12738
rect 26962 12686 26964 12738
rect 26572 11778 26628 11788
rect 26796 12068 26852 12078
rect 26796 11506 26852 12012
rect 26908 11732 26964 12686
rect 27020 12738 27076 12750
rect 27020 12686 27022 12738
rect 27074 12686 27076 12738
rect 27020 12178 27076 12686
rect 27916 12404 27972 12910
rect 28140 12516 28196 13804
rect 28364 13858 28420 15260
rect 28588 15090 28644 15102
rect 28588 15038 28590 15090
rect 28642 15038 28644 15090
rect 28588 14756 28644 15038
rect 28588 14690 28644 14700
rect 28588 14532 28644 14542
rect 28700 14532 28756 15820
rect 29484 15148 29540 17724
rect 29708 17714 29764 17724
rect 29820 17668 29876 20188
rect 29932 19908 29988 19918
rect 29932 19458 29988 19852
rect 29932 19406 29934 19458
rect 29986 19406 29988 19458
rect 29932 19394 29988 19406
rect 30044 19236 30100 24892
rect 30156 24610 30212 25228
rect 30156 24558 30158 24610
rect 30210 24558 30212 24610
rect 30156 24546 30212 24558
rect 30716 24610 30772 26126
rect 30716 24558 30718 24610
rect 30770 24558 30772 24610
rect 30192 24332 30456 24342
rect 30248 24276 30296 24332
rect 30352 24276 30400 24332
rect 30192 24266 30456 24276
rect 30492 23940 30548 23950
rect 30492 23378 30548 23884
rect 30604 23828 30660 23838
rect 30716 23828 30772 24558
rect 30660 23772 30772 23828
rect 30604 23734 30660 23772
rect 30492 23326 30494 23378
rect 30546 23326 30548 23378
rect 30492 23314 30548 23326
rect 30380 23268 30436 23278
rect 30380 23174 30436 23212
rect 30716 23156 30772 23166
rect 30716 23062 30772 23100
rect 30192 22764 30456 22774
rect 30248 22708 30296 22764
rect 30352 22708 30400 22764
rect 30828 22708 30884 26908
rect 31164 26404 31220 27244
rect 31164 26310 31220 26348
rect 31276 26964 31332 27002
rect 31052 26290 31108 26302
rect 31052 26238 31054 26290
rect 31106 26238 31108 26290
rect 31052 25508 31108 26238
rect 31276 26178 31332 26908
rect 31276 26126 31278 26178
rect 31330 26126 31332 26178
rect 31276 26114 31332 26126
rect 30940 24052 30996 24062
rect 31052 24052 31108 25452
rect 31388 24164 31444 31612
rect 31500 31218 31556 31230
rect 31500 31166 31502 31218
rect 31554 31166 31556 31218
rect 31500 29652 31556 31166
rect 31612 31108 31668 31724
rect 31836 31714 31892 31724
rect 32172 31780 32228 35420
rect 32396 35698 32452 35710
rect 32396 35646 32398 35698
rect 32450 35646 32452 35698
rect 32396 34244 32452 35646
rect 32508 35588 32564 36318
rect 33180 36258 33236 36270
rect 33180 36206 33182 36258
rect 33234 36206 33236 36258
rect 33068 35588 33124 35598
rect 32508 35586 33124 35588
rect 32508 35534 33070 35586
rect 33122 35534 33124 35586
rect 32508 35532 33124 35534
rect 32844 34916 32900 34926
rect 32956 34916 33012 35532
rect 33068 35522 33124 35532
rect 32844 34914 33012 34916
rect 32844 34862 32846 34914
rect 32898 34862 33012 34914
rect 32844 34860 33012 34862
rect 33068 35364 33124 35374
rect 32396 34188 32564 34244
rect 32396 34020 32452 34030
rect 32396 33906 32452 33964
rect 32396 33854 32398 33906
rect 32450 33854 32452 33906
rect 32396 33842 32452 33854
rect 32508 33796 32564 34188
rect 32396 33458 32452 33470
rect 32396 33406 32398 33458
rect 32450 33406 32452 33458
rect 32284 33234 32340 33246
rect 32284 33182 32286 33234
rect 32338 33182 32340 33234
rect 32284 32004 32340 33182
rect 32396 33124 32452 33406
rect 32396 33058 32452 33068
rect 32284 31938 32340 31948
rect 32172 31686 32228 31724
rect 32396 31778 32452 31790
rect 32396 31726 32398 31778
rect 32450 31726 32452 31778
rect 31612 30994 31668 31052
rect 31612 30942 31614 30994
rect 31666 30942 31668 30994
rect 31612 30930 31668 30942
rect 32060 31666 32116 31678
rect 32060 31614 32062 31666
rect 32114 31614 32116 31666
rect 31724 30212 31780 30222
rect 31724 30118 31780 30156
rect 32060 29764 32116 31614
rect 32284 31668 32340 31678
rect 32060 29708 32228 29764
rect 31500 29596 31668 29652
rect 31612 29540 31668 29596
rect 32060 29540 32116 29550
rect 31612 29538 32116 29540
rect 31612 29486 32062 29538
rect 32114 29486 32116 29538
rect 31612 29484 32116 29486
rect 31500 29428 31556 29438
rect 31500 29314 31556 29372
rect 31500 29262 31502 29314
rect 31554 29262 31556 29314
rect 31500 29250 31556 29262
rect 31612 29202 31668 29214
rect 31612 29150 31614 29202
rect 31666 29150 31668 29202
rect 31500 28868 31556 28878
rect 31500 27858 31556 28812
rect 31612 28644 31668 29150
rect 31612 28578 31668 28588
rect 31500 27806 31502 27858
rect 31554 27806 31556 27858
rect 31500 27794 31556 27806
rect 31724 27860 31780 29484
rect 32060 29474 32116 29484
rect 32172 29428 32228 29708
rect 32172 29362 32228 29372
rect 32284 29650 32340 31612
rect 32396 31556 32452 31726
rect 32396 31490 32452 31500
rect 32396 31332 32452 31342
rect 32508 31332 32564 33740
rect 32844 33234 32900 34860
rect 33068 34354 33124 35308
rect 33180 34580 33236 36206
rect 33292 35700 33348 35710
rect 33292 35606 33348 35644
rect 33516 35476 33572 35486
rect 33516 35382 33572 35420
rect 33964 35474 34020 35486
rect 33964 35422 33966 35474
rect 34018 35422 34020 35474
rect 33628 35364 33684 35374
rect 33516 35026 33572 35038
rect 33516 34974 33518 35026
rect 33570 34974 33572 35026
rect 33180 34524 33460 34580
rect 33068 34302 33070 34354
rect 33122 34302 33124 34354
rect 33068 34290 33124 34302
rect 33292 34356 33348 34366
rect 33292 34262 33348 34300
rect 33180 34130 33236 34142
rect 33180 34078 33182 34130
rect 33234 34078 33236 34130
rect 33180 33460 33236 34078
rect 33180 33394 33236 33404
rect 32844 33182 32846 33234
rect 32898 33182 32900 33234
rect 32844 33170 32900 33182
rect 33180 33124 33236 33134
rect 33236 33068 33348 33124
rect 33180 33058 33236 33068
rect 33292 32786 33348 33068
rect 33292 32734 33294 32786
rect 33346 32734 33348 32786
rect 33292 32722 33348 32734
rect 33404 32564 33460 34524
rect 33516 33460 33572 34974
rect 33516 33394 33572 33404
rect 33292 32508 33460 32564
rect 33180 31890 33236 31902
rect 33180 31838 33182 31890
rect 33234 31838 33236 31890
rect 33180 31668 33236 31838
rect 33180 31602 33236 31612
rect 32452 31276 32564 31332
rect 32844 31554 32900 31566
rect 32844 31502 32846 31554
rect 32898 31502 32900 31554
rect 32396 31266 32452 31276
rect 32284 29598 32286 29650
rect 32338 29598 32340 29650
rect 32060 28756 32116 28766
rect 31724 27746 31780 27804
rect 31724 27694 31726 27746
rect 31778 27694 31780 27746
rect 31724 27682 31780 27694
rect 31836 27972 31892 27982
rect 31724 27076 31780 27086
rect 31724 26982 31780 27020
rect 31836 26850 31892 27916
rect 31836 26798 31838 26850
rect 31890 26798 31892 26850
rect 31836 26786 31892 26798
rect 31836 26404 31892 26414
rect 31836 24836 31892 26348
rect 31724 24834 31892 24836
rect 31724 24782 31838 24834
rect 31890 24782 31892 24834
rect 31724 24780 31892 24782
rect 31500 24164 31556 24174
rect 31388 24162 31556 24164
rect 31388 24110 31502 24162
rect 31554 24110 31556 24162
rect 31388 24108 31556 24110
rect 31500 24098 31556 24108
rect 31724 24164 31780 24780
rect 31836 24770 31892 24780
rect 31948 24612 32004 24622
rect 32060 24612 32116 28700
rect 32284 28420 32340 29598
rect 32620 30772 32676 30782
rect 32396 29202 32452 29214
rect 32396 29150 32398 29202
rect 32450 29150 32452 29202
rect 32396 29092 32452 29150
rect 32396 29026 32452 29036
rect 32396 28644 32452 28654
rect 32396 28550 32452 28588
rect 32284 28364 32452 28420
rect 32172 27972 32228 27982
rect 32172 27858 32228 27916
rect 32172 27806 32174 27858
rect 32226 27806 32228 27858
rect 32172 27794 32228 27806
rect 32284 27970 32340 27982
rect 32284 27918 32286 27970
rect 32338 27918 32340 27970
rect 32172 27636 32228 27646
rect 32172 26402 32228 27580
rect 32284 26962 32340 27918
rect 32284 26910 32286 26962
rect 32338 26910 32340 26962
rect 32284 26898 32340 26910
rect 32396 26514 32452 28364
rect 32396 26462 32398 26514
rect 32450 26462 32452 26514
rect 32396 26450 32452 26462
rect 32508 27074 32564 27086
rect 32508 27022 32510 27074
rect 32562 27022 32564 27074
rect 32172 26350 32174 26402
rect 32226 26350 32228 26402
rect 32172 26338 32228 26350
rect 32508 26178 32564 27022
rect 32620 26404 32676 30716
rect 32844 29652 32900 31502
rect 33292 30324 33348 32508
rect 33628 32340 33684 35308
rect 33852 34914 33908 34926
rect 33852 34862 33854 34914
rect 33906 34862 33908 34914
rect 33628 32274 33684 32284
rect 33740 34130 33796 34142
rect 33740 34078 33742 34130
rect 33794 34078 33796 34130
rect 33404 32116 33460 32126
rect 33404 31780 33460 32060
rect 33740 31892 33796 34078
rect 33852 34020 33908 34862
rect 33964 34130 34020 35422
rect 34412 35308 34468 36430
rect 34412 35252 34692 35308
rect 34524 34914 34580 34926
rect 34524 34862 34526 34914
rect 34578 34862 34580 34914
rect 34300 34804 34356 34814
rect 34188 34802 34356 34804
rect 34188 34750 34302 34802
rect 34354 34750 34356 34802
rect 34188 34748 34356 34750
rect 33964 34078 33966 34130
rect 34018 34078 34020 34130
rect 33964 34066 34020 34078
rect 34076 34132 34132 34142
rect 34188 34132 34244 34748
rect 34300 34738 34356 34748
rect 34132 34076 34244 34132
rect 34300 34130 34356 34142
rect 34300 34078 34302 34130
rect 34354 34078 34356 34130
rect 34076 34066 34132 34076
rect 33852 33954 33908 33964
rect 34300 33796 34356 34078
rect 34300 33730 34356 33740
rect 33964 33684 34020 33694
rect 33964 33458 34020 33628
rect 34524 33684 34580 34862
rect 34524 33618 34580 33628
rect 33964 33406 33966 33458
rect 34018 33406 34020 33458
rect 33852 33346 33908 33358
rect 33852 33294 33854 33346
rect 33906 33294 33908 33346
rect 33852 33236 33908 33294
rect 33852 33170 33908 33180
rect 33740 31826 33796 31836
rect 33852 32450 33908 32462
rect 33852 32398 33854 32450
rect 33906 32398 33908 32450
rect 33404 31220 33460 31724
rect 33516 31778 33572 31790
rect 33516 31726 33518 31778
rect 33570 31726 33572 31778
rect 33516 31556 33572 31726
rect 33516 31490 33572 31500
rect 33740 31220 33796 31230
rect 33852 31220 33908 32398
rect 33404 31218 33572 31220
rect 33404 31166 33406 31218
rect 33458 31166 33572 31218
rect 33404 31164 33572 31166
rect 33404 31154 33460 31164
rect 33516 30324 33572 31164
rect 33796 31164 33908 31220
rect 33740 31154 33796 31164
rect 33964 30996 34020 33406
rect 34188 32452 34244 32462
rect 34300 32452 34356 32462
rect 34244 32450 34356 32452
rect 34244 32398 34302 32450
rect 34354 32398 34356 32450
rect 34244 32396 34356 32398
rect 33292 30268 33460 30324
rect 32844 29586 32900 29596
rect 33292 30098 33348 30110
rect 33292 30046 33294 30098
rect 33346 30046 33348 30098
rect 33180 29540 33236 29550
rect 33180 29446 33236 29484
rect 33068 29426 33124 29438
rect 33068 29374 33070 29426
rect 33122 29374 33124 29426
rect 33068 29092 33124 29374
rect 33292 29428 33348 30046
rect 33068 29026 33124 29036
rect 33180 29314 33236 29326
rect 33180 29262 33182 29314
rect 33234 29262 33236 29314
rect 33180 28756 33236 29262
rect 33180 28690 33236 28700
rect 33292 28644 33348 29372
rect 33404 29316 33460 30268
rect 33516 30258 33572 30268
rect 33740 30940 34020 30996
rect 34076 32004 34132 32014
rect 33404 29250 33460 29260
rect 33292 28082 33348 28588
rect 33740 28532 33796 30940
rect 34076 30210 34132 31948
rect 34076 30158 34078 30210
rect 34130 30158 34132 30210
rect 34076 30100 34132 30158
rect 34076 30034 34132 30044
rect 33740 28466 33796 28476
rect 33852 29986 33908 29998
rect 33852 29934 33854 29986
rect 33906 29934 33908 29986
rect 33292 28030 33294 28082
rect 33346 28030 33348 28082
rect 33292 28018 33348 28030
rect 33628 28420 33684 28430
rect 33628 27970 33684 28364
rect 33852 28196 33908 29934
rect 33964 29986 34020 29998
rect 33964 29934 33966 29986
rect 34018 29934 34020 29986
rect 33964 29426 34020 29934
rect 34188 29764 34244 32396
rect 34300 32386 34356 32396
rect 34636 31108 34692 35252
rect 34748 34916 34804 34926
rect 34748 33236 34804 34860
rect 34748 33122 34804 33180
rect 34748 33070 34750 33122
rect 34802 33070 34804 33122
rect 34748 32116 34804 33070
rect 34748 32050 34804 32060
rect 34524 31052 34692 31108
rect 34524 30548 34580 31052
rect 34636 30884 34692 30894
rect 34636 30882 34916 30884
rect 34636 30830 34638 30882
rect 34690 30830 34916 30882
rect 34636 30828 34916 30830
rect 34636 30818 34692 30828
rect 34524 30492 34692 30548
rect 34524 30324 34580 30334
rect 34524 30230 34580 30268
rect 34188 29698 34244 29708
rect 34300 30210 34356 30222
rect 34300 30158 34302 30210
rect 34354 30158 34356 30210
rect 33964 29374 33966 29426
rect 34018 29374 34020 29426
rect 33964 29362 34020 29374
rect 34300 29316 34356 30158
rect 34300 29250 34356 29260
rect 33964 28700 34580 28756
rect 33964 28642 34020 28700
rect 33964 28590 33966 28642
rect 34018 28590 34020 28642
rect 33964 28578 34020 28590
rect 34524 28642 34580 28700
rect 34524 28590 34526 28642
rect 34578 28590 34580 28642
rect 34524 28578 34580 28590
rect 34412 28308 34468 28318
rect 34636 28308 34692 30492
rect 34860 30210 34916 30828
rect 34860 30158 34862 30210
rect 34914 30158 34916 30210
rect 34860 29988 34916 30158
rect 34860 29922 34916 29932
rect 34972 29428 35028 37212
rect 35532 36596 35588 39228
rect 35868 39060 35924 39228
rect 36064 39200 36176 40000
rect 38528 39200 38640 40000
rect 40992 39200 41104 40000
rect 43456 39200 43568 40000
rect 45920 39200 46032 40000
rect 46172 39228 47012 39284
rect 36092 39060 36148 39200
rect 35868 39004 36148 39060
rect 38444 36596 38500 36606
rect 38556 36596 38612 39200
rect 39564 37604 39620 37614
rect 35532 36594 36596 36596
rect 35532 36542 35534 36594
rect 35586 36542 36596 36594
rect 35532 36540 36596 36542
rect 35532 36530 35588 36540
rect 36540 36482 36596 36540
rect 38444 36594 38724 36596
rect 38444 36542 38446 36594
rect 38498 36542 38724 36594
rect 38444 36540 38724 36542
rect 38444 36530 38500 36540
rect 36540 36430 36542 36482
rect 36594 36430 36596 36482
rect 36540 36418 36596 36430
rect 38668 36482 38724 36540
rect 38668 36430 38670 36482
rect 38722 36430 38724 36482
rect 38668 36418 38724 36430
rect 39228 36482 39284 36494
rect 39228 36430 39230 36482
rect 39282 36430 39284 36482
rect 36316 36258 36372 36270
rect 36316 36206 36318 36258
rect 36370 36206 36372 36258
rect 35420 35586 35476 35598
rect 35420 35534 35422 35586
rect 35474 35534 35476 35586
rect 35420 34916 35476 35534
rect 35420 34850 35476 34860
rect 35868 34914 35924 34926
rect 35868 34862 35870 34914
rect 35922 34862 35924 34914
rect 35756 34690 35812 34702
rect 35756 34638 35758 34690
rect 35810 34638 35812 34690
rect 35644 34468 35700 34478
rect 35756 34468 35812 34638
rect 35700 34412 35812 34468
rect 35644 31220 35700 34412
rect 35868 33570 35924 34862
rect 36204 34916 36260 34926
rect 36204 34822 36260 34860
rect 35868 33518 35870 33570
rect 35922 33518 35924 33570
rect 35868 33506 35924 33518
rect 36092 34018 36148 34030
rect 36092 33966 36094 34018
rect 36146 33966 36148 34018
rect 35756 32450 35812 32462
rect 35756 32398 35758 32450
rect 35810 32398 35812 32450
rect 35756 31780 35812 32398
rect 35756 31714 35812 31724
rect 36092 31220 36148 33966
rect 36204 33460 36260 33470
rect 36204 33366 36260 33404
rect 36316 32676 36372 36206
rect 37212 35812 37268 35822
rect 38220 35812 38276 35822
rect 37212 35810 38276 35812
rect 37212 35758 37214 35810
rect 37266 35758 38222 35810
rect 38274 35758 38276 35810
rect 37212 35756 38276 35758
rect 37212 35746 37268 35756
rect 36876 35698 36932 35710
rect 36876 35646 36878 35698
rect 36930 35646 36932 35698
rect 36540 35586 36596 35598
rect 36540 35534 36542 35586
rect 36594 35534 36596 35586
rect 36540 35476 36596 35534
rect 36540 35410 36596 35420
rect 36764 35252 36820 35262
rect 36428 34690 36484 34702
rect 36428 34638 36430 34690
rect 36482 34638 36484 34690
rect 36428 34468 36484 34638
rect 36428 34402 36484 34412
rect 36540 34690 36596 34702
rect 36540 34638 36542 34690
rect 36594 34638 36596 34690
rect 36540 34356 36596 34638
rect 36540 34290 36596 34300
rect 36540 34132 36596 34142
rect 36540 34038 36596 34076
rect 36652 33348 36708 33358
rect 36428 33236 36484 33246
rect 36428 33142 36484 33180
rect 35644 31126 35700 31164
rect 35868 31164 36148 31220
rect 35868 30322 35924 31164
rect 36092 31106 36148 31164
rect 36092 31054 36094 31106
rect 36146 31054 36148 31106
rect 36092 31042 36148 31054
rect 36204 32620 36372 32676
rect 36428 32900 36484 32910
rect 35980 30994 36036 31006
rect 35980 30942 35982 30994
rect 36034 30942 36036 30994
rect 35980 30436 36036 30942
rect 36092 30436 36148 30446
rect 35980 30380 36092 30436
rect 36092 30342 36148 30380
rect 35868 30270 35870 30322
rect 35922 30270 35924 30322
rect 35084 30100 35140 30110
rect 35140 30044 35252 30100
rect 35084 30034 35140 30044
rect 35196 29988 35252 30044
rect 35196 29986 35700 29988
rect 35196 29934 35198 29986
rect 35250 29934 35700 29986
rect 35196 29932 35700 29934
rect 35196 29922 35252 29932
rect 35644 29650 35700 29932
rect 35644 29598 35646 29650
rect 35698 29598 35700 29650
rect 35644 29586 35700 29598
rect 35868 29652 35924 30270
rect 36204 29652 36260 32620
rect 36316 32452 36372 32462
rect 36428 32452 36484 32844
rect 36652 32562 36708 33292
rect 36652 32510 36654 32562
rect 36706 32510 36708 32562
rect 36652 32498 36708 32510
rect 36316 32450 36484 32452
rect 36316 32398 36318 32450
rect 36370 32398 36484 32450
rect 36316 32396 36484 32398
rect 36316 32386 36372 32396
rect 36540 32338 36596 32350
rect 36540 32286 36542 32338
rect 36594 32286 36596 32338
rect 36540 31780 36596 32286
rect 36540 31714 36596 31724
rect 36540 30996 36596 31006
rect 36428 30436 36484 30446
rect 36540 30436 36596 30940
rect 36652 30884 36708 30894
rect 36652 30790 36708 30828
rect 36428 30434 36596 30436
rect 36428 30382 36430 30434
rect 36482 30382 36596 30434
rect 36428 30380 36596 30382
rect 36652 30436 36708 30446
rect 36428 30370 36484 30380
rect 35868 29586 35924 29596
rect 36092 29596 36260 29652
rect 36428 30212 36484 30222
rect 35420 29538 35476 29550
rect 35420 29486 35422 29538
rect 35474 29486 35476 29538
rect 34972 29372 35140 29428
rect 34860 29316 34916 29326
rect 34916 29260 35028 29316
rect 34860 29250 34916 29260
rect 34860 28530 34916 28542
rect 34860 28478 34862 28530
rect 34914 28478 34916 28530
rect 34748 28420 34804 28430
rect 34748 28326 34804 28364
rect 33852 28140 34356 28196
rect 33628 27918 33630 27970
rect 33682 27918 33684 27970
rect 33628 27906 33684 27918
rect 33740 27860 33796 27870
rect 33852 27860 33908 27870
rect 33740 27858 33852 27860
rect 33740 27806 33742 27858
rect 33794 27806 33852 27858
rect 33740 27804 33852 27806
rect 33740 27794 33796 27804
rect 32620 26338 32676 26348
rect 32732 26852 32788 26862
rect 32508 26126 32510 26178
rect 32562 26126 32564 26178
rect 32508 26114 32564 26126
rect 32732 25508 32788 26796
rect 33740 26402 33796 26414
rect 33740 26350 33742 26402
rect 33794 26350 33796 26402
rect 33068 26292 33124 26302
rect 33068 26198 33124 26236
rect 33292 26292 33348 26302
rect 32732 25442 32788 25452
rect 33068 25282 33124 25294
rect 33068 25230 33070 25282
rect 33122 25230 33124 25282
rect 32172 24612 32228 24622
rect 32060 24610 32228 24612
rect 32060 24558 32174 24610
rect 32226 24558 32228 24610
rect 32060 24556 32228 24558
rect 31724 24098 31780 24108
rect 31836 24164 31892 24174
rect 31948 24164 32004 24556
rect 31836 24162 32004 24164
rect 31836 24110 31838 24162
rect 31890 24110 32004 24162
rect 31836 24108 32004 24110
rect 31836 24098 31892 24108
rect 31052 23996 31332 24052
rect 30940 23828 30996 23996
rect 31052 23828 31108 23838
rect 30940 23826 31108 23828
rect 30940 23774 31054 23826
rect 31106 23774 31108 23826
rect 30940 23772 31108 23774
rect 31052 23762 31108 23772
rect 31164 23828 31220 23838
rect 31052 23156 31108 23166
rect 31164 23156 31220 23772
rect 31052 23154 31220 23156
rect 31052 23102 31054 23154
rect 31106 23102 31220 23154
rect 31052 23100 31220 23102
rect 31276 23154 31332 23996
rect 31276 23102 31278 23154
rect 31330 23102 31332 23154
rect 31052 23090 31108 23100
rect 31276 23090 31332 23102
rect 31500 23492 31556 23502
rect 30192 22698 30456 22708
rect 30604 22652 30884 22708
rect 30604 22484 30660 22652
rect 30492 22428 30660 22484
rect 30828 22484 30884 22494
rect 30828 22482 31444 22484
rect 30828 22430 30830 22482
rect 30882 22430 31444 22482
rect 30828 22428 31444 22430
rect 30380 21588 30436 21598
rect 30380 21494 30436 21532
rect 30268 21474 30324 21486
rect 30268 21422 30270 21474
rect 30322 21422 30324 21474
rect 30268 21364 30324 21422
rect 30492 21476 30548 22428
rect 30828 22418 30884 22428
rect 31388 22370 31444 22428
rect 31388 22318 31390 22370
rect 31442 22318 31444 22370
rect 31388 22306 31444 22318
rect 30604 22260 30660 22270
rect 30604 22166 30660 22204
rect 31052 22260 31108 22270
rect 30716 22146 30772 22158
rect 30716 22094 30718 22146
rect 30770 22094 30772 22146
rect 30716 21588 30772 22094
rect 30940 22146 30996 22158
rect 30940 22094 30942 22146
rect 30994 22094 30996 22146
rect 30940 21924 30996 22094
rect 30940 21858 30996 21868
rect 31052 21810 31108 22204
rect 31052 21758 31054 21810
rect 31106 21758 31108 21810
rect 31052 21746 31108 21758
rect 31164 22258 31220 22270
rect 31164 22206 31166 22258
rect 31218 22206 31220 22258
rect 31164 21700 31220 22206
rect 30716 21532 30996 21588
rect 30492 21420 30772 21476
rect 30268 21298 30324 21308
rect 30192 21196 30456 21206
rect 30248 21140 30296 21196
rect 30352 21140 30400 21196
rect 30192 21130 30456 21140
rect 30268 20580 30324 20590
rect 30716 20580 30772 21420
rect 30828 20804 30884 20814
rect 30828 20710 30884 20748
rect 30940 20580 30996 21532
rect 31164 21364 31220 21644
rect 31164 21298 31220 21308
rect 31276 22036 31332 22046
rect 31164 20916 31220 20926
rect 31276 20916 31332 21980
rect 31220 20860 31332 20916
rect 31388 21586 31444 21598
rect 31388 21534 31390 21586
rect 31442 21534 31444 21586
rect 31164 20822 31220 20860
rect 31388 20804 31444 21534
rect 31388 20738 31444 20748
rect 31164 20580 31220 20590
rect 30716 20524 30884 20580
rect 30940 20524 31164 20580
rect 30268 20486 30324 20524
rect 30156 20356 30212 20366
rect 30156 20242 30212 20300
rect 30156 20190 30158 20242
rect 30210 20190 30212 20242
rect 30156 20178 30212 20190
rect 30192 19628 30456 19638
rect 30248 19572 30296 19628
rect 30352 19572 30400 19628
rect 30192 19562 30456 19572
rect 30716 19572 30772 19582
rect 29932 19180 30100 19236
rect 30268 19234 30324 19246
rect 30268 19182 30270 19234
rect 30322 19182 30324 19234
rect 29932 18450 29988 19180
rect 30268 19124 30324 19182
rect 30268 19058 30324 19068
rect 29932 18398 29934 18450
rect 29986 18398 29988 18450
rect 29932 18386 29988 18398
rect 30044 19010 30100 19022
rect 30044 18958 30046 19010
rect 30098 18958 30100 19010
rect 30044 18452 30100 18958
rect 30716 19012 30772 19516
rect 30716 18946 30772 18956
rect 30044 18386 30100 18396
rect 30492 18452 30548 18462
rect 30492 18358 30548 18396
rect 30192 18060 30456 18070
rect 30248 18004 30296 18060
rect 30352 18004 30400 18060
rect 30192 17994 30456 18004
rect 30828 17668 30884 20524
rect 30940 20132 30996 20142
rect 30940 19124 30996 20076
rect 30940 19058 30996 19068
rect 31052 20018 31108 20030
rect 31052 19966 31054 20018
rect 31106 19966 31108 20018
rect 31052 18340 31108 19966
rect 31052 18274 31108 18284
rect 30828 17612 30996 17668
rect 29820 17602 29876 17612
rect 30380 17556 30436 17566
rect 30380 17106 30436 17500
rect 30380 17054 30382 17106
rect 30434 17054 30436 17106
rect 30380 17042 30436 17054
rect 30716 17554 30772 17566
rect 30716 17502 30718 17554
rect 30770 17502 30772 17554
rect 30604 16884 30660 16894
rect 30604 16790 30660 16828
rect 29932 16772 29988 16782
rect 29932 16770 30100 16772
rect 29932 16718 29934 16770
rect 29986 16718 30100 16770
rect 29932 16716 30100 16718
rect 29932 16706 29988 16716
rect 29932 16098 29988 16110
rect 29932 16046 29934 16098
rect 29986 16046 29988 16098
rect 29708 15652 29764 15662
rect 29708 15426 29764 15596
rect 29708 15374 29710 15426
rect 29762 15374 29764 15426
rect 29708 15362 29764 15374
rect 29260 15092 29540 15148
rect 29596 15314 29652 15326
rect 29596 15262 29598 15314
rect 29650 15262 29652 15314
rect 29596 15204 29652 15262
rect 29932 15316 29988 16046
rect 29932 15250 29988 15260
rect 30044 16100 30100 16716
rect 30192 16492 30456 16502
rect 30248 16436 30296 16492
rect 30352 16436 30400 16492
rect 30192 16426 30456 16436
rect 30716 16324 30772 17502
rect 30828 16660 30884 16670
rect 30940 16660 30996 17612
rect 30828 16658 30996 16660
rect 30828 16606 30830 16658
rect 30882 16606 30996 16658
rect 30828 16604 30996 16606
rect 30828 16594 30884 16604
rect 31164 16548 31220 20524
rect 31500 19906 31556 23436
rect 31612 23380 31668 23390
rect 31612 23286 31668 23324
rect 32060 23380 32116 23390
rect 31948 23268 32004 23278
rect 31948 21924 32004 23212
rect 32060 23154 32116 23324
rect 32060 23102 32062 23154
rect 32114 23102 32116 23154
rect 32060 23090 32116 23102
rect 32172 22370 32228 24556
rect 33068 24612 33124 25230
rect 33068 24546 33124 24556
rect 33180 24722 33236 24734
rect 33180 24670 33182 24722
rect 33234 24670 33236 24722
rect 32620 23938 32676 23950
rect 32620 23886 32622 23938
rect 32674 23886 32676 23938
rect 32396 23828 32452 23838
rect 32396 23734 32452 23772
rect 32620 23492 32676 23886
rect 32620 23426 32676 23436
rect 33180 23380 33236 24670
rect 33180 23314 33236 23324
rect 33292 23268 33348 26236
rect 33404 25506 33460 25518
rect 33404 25454 33406 25506
rect 33458 25454 33460 25506
rect 33404 25396 33460 25454
rect 33404 25330 33460 25340
rect 33628 25506 33684 25518
rect 33628 25454 33630 25506
rect 33682 25454 33684 25506
rect 33628 24836 33684 25454
rect 33628 24770 33684 24780
rect 33740 24724 33796 26350
rect 33852 25508 33908 27804
rect 34188 27858 34244 27870
rect 34188 27806 34190 27858
rect 34242 27806 34244 27858
rect 34188 27748 34244 27806
rect 34188 27682 34244 27692
rect 33964 27074 34020 27086
rect 33964 27022 33966 27074
rect 34018 27022 34020 27074
rect 33964 25730 34020 27022
rect 33964 25678 33966 25730
rect 34018 25678 34020 25730
rect 33964 25666 34020 25678
rect 34300 27076 34356 28140
rect 33852 25452 34020 25508
rect 33740 24658 33796 24668
rect 33628 24610 33684 24622
rect 33628 24558 33630 24610
rect 33682 24558 33684 24610
rect 33628 24500 33684 24558
rect 33628 24434 33684 24444
rect 33852 24052 33908 24062
rect 33852 23958 33908 23996
rect 33404 23940 33460 23950
rect 33404 23604 33460 23884
rect 33404 23538 33460 23548
rect 33628 23548 33684 23558
rect 33964 23548 34020 25452
rect 34076 24836 34132 24846
rect 34076 24724 34132 24780
rect 34076 24722 34244 24724
rect 34076 24670 34078 24722
rect 34130 24670 34244 24722
rect 34076 24668 34244 24670
rect 34076 24658 34132 24668
rect 34188 24164 34244 24668
rect 33516 23380 33572 23390
rect 33628 23380 33684 23492
rect 33292 23202 33348 23212
rect 33404 23378 33684 23380
rect 33404 23326 33518 23378
rect 33570 23326 33684 23378
rect 33404 23324 33684 23326
rect 33740 23492 34020 23548
rect 34076 23938 34132 23950
rect 34076 23886 34078 23938
rect 34130 23886 34132 23938
rect 33740 23378 33796 23492
rect 33740 23326 33742 23378
rect 33794 23326 33796 23378
rect 32508 23156 32564 23166
rect 32508 23062 32564 23100
rect 32172 22318 32174 22370
rect 32226 22318 32228 22370
rect 32172 22306 32228 22318
rect 32732 22370 32788 22382
rect 32732 22318 32734 22370
rect 32786 22318 32788 22370
rect 31948 21810 32004 21868
rect 31948 21758 31950 21810
rect 32002 21758 32004 21810
rect 31948 21746 32004 21758
rect 32284 22258 32340 22270
rect 32284 22206 32286 22258
rect 32338 22206 32340 22258
rect 32284 21700 32340 22206
rect 32060 21644 32340 21700
rect 32732 21700 32788 22318
rect 31612 21588 31668 21598
rect 31612 20914 31668 21532
rect 31612 20862 31614 20914
rect 31666 20862 31668 20914
rect 31612 20850 31668 20862
rect 31500 19854 31502 19906
rect 31554 19854 31556 19906
rect 31500 19842 31556 19854
rect 31500 18452 31556 18462
rect 31276 17556 31332 17566
rect 31276 17462 31332 17500
rect 30940 16492 31220 16548
rect 30828 16324 30884 16334
rect 30716 16268 30828 16324
rect 30044 16044 30324 16100
rect 30044 15148 30100 16044
rect 30268 15986 30324 16044
rect 30268 15934 30270 15986
rect 30322 15934 30324 15986
rect 30268 15922 30324 15934
rect 30828 15538 30884 16268
rect 30828 15486 30830 15538
rect 30882 15486 30884 15538
rect 30828 15474 30884 15486
rect 29596 15138 29652 15148
rect 29708 15092 30100 15148
rect 28644 14476 28756 14532
rect 28812 14756 28868 14766
rect 28588 14438 28644 14476
rect 28812 14420 28868 14700
rect 29148 14532 29204 14542
rect 28812 14354 28868 14364
rect 29036 14530 29204 14532
rect 29036 14478 29150 14530
rect 29202 14478 29204 14530
rect 29036 14476 29204 14478
rect 28364 13806 28366 13858
rect 28418 13806 28420 13858
rect 28364 13794 28420 13806
rect 28252 13748 28308 13758
rect 28252 13654 28308 13692
rect 28476 13746 28532 13758
rect 28476 13694 28478 13746
rect 28530 13694 28532 13746
rect 28140 12460 28308 12516
rect 27916 12348 28084 12404
rect 28028 12292 28084 12348
rect 28140 12292 28196 12302
rect 28028 12236 28140 12292
rect 28140 12198 28196 12236
rect 27020 12126 27022 12178
rect 27074 12126 27076 12178
rect 27020 12114 27076 12126
rect 27916 12178 27972 12190
rect 27916 12126 27918 12178
rect 27970 12126 27972 12178
rect 27692 12068 27748 12078
rect 27692 12066 27860 12068
rect 27692 12014 27694 12066
rect 27746 12014 27860 12066
rect 27692 12012 27860 12014
rect 27692 12002 27748 12012
rect 26908 11676 27748 11732
rect 26796 11454 26798 11506
rect 26850 11454 26852 11506
rect 26796 11442 26852 11454
rect 27020 10276 27076 11676
rect 27244 11508 27300 11518
rect 27244 11414 27300 11452
rect 27468 11506 27524 11518
rect 27468 11454 27470 11506
rect 27522 11454 27524 11506
rect 27132 11394 27188 11406
rect 27132 11342 27134 11394
rect 27186 11342 27188 11394
rect 27132 10500 27188 11342
rect 27468 10724 27524 11454
rect 27692 11394 27748 11676
rect 27692 11342 27694 11394
rect 27746 11342 27748 11394
rect 27692 11330 27748 11342
rect 27804 11172 27860 12012
rect 27804 11106 27860 11116
rect 27804 10836 27860 10846
rect 27916 10836 27972 12126
rect 28028 11620 28084 11630
rect 28028 11394 28084 11564
rect 28028 11342 28030 11394
rect 28082 11342 28084 11394
rect 28028 11060 28084 11342
rect 28140 11396 28196 11406
rect 28140 11302 28196 11340
rect 28028 10994 28084 11004
rect 27804 10834 27972 10836
rect 27804 10782 27806 10834
rect 27858 10782 27972 10834
rect 27804 10780 27972 10782
rect 27804 10770 27860 10780
rect 27468 10658 27524 10668
rect 27692 10500 27748 10510
rect 27132 10498 27748 10500
rect 27132 10446 27694 10498
rect 27746 10446 27748 10498
rect 27132 10444 27748 10446
rect 27020 10220 27412 10276
rect 26460 9426 26516 9436
rect 26572 9714 26628 9726
rect 26572 9662 26574 9714
rect 26626 9662 26628 9714
rect 26460 8484 26516 8494
rect 26572 8484 26628 9662
rect 26908 9602 26964 9614
rect 26908 9550 26910 9602
rect 26962 9550 26964 9602
rect 26908 9154 26964 9550
rect 26908 9102 26910 9154
rect 26962 9102 26964 9154
rect 26908 9090 26964 9102
rect 26460 8482 26628 8484
rect 26460 8430 26462 8482
rect 26514 8430 26628 8482
rect 26460 8428 26628 8430
rect 27356 8932 27412 10220
rect 26460 8418 26516 8428
rect 26796 8260 26852 8270
rect 26796 8166 26852 8204
rect 27356 8146 27412 8876
rect 27356 8094 27358 8146
rect 27410 8094 27412 8146
rect 27356 8082 27412 8094
rect 27468 8260 27524 8270
rect 26908 7700 26964 7710
rect 26908 6804 26964 7644
rect 27468 7140 27524 8204
rect 27468 7074 27524 7084
rect 27692 6804 27748 10444
rect 28252 10164 28308 12460
rect 28252 10098 28308 10108
rect 28364 11396 28420 11406
rect 28476 11396 28532 13694
rect 29036 13748 29092 14476
rect 29148 14466 29204 14476
rect 29036 13654 29092 13692
rect 28924 13076 28980 13086
rect 28700 12964 28756 12974
rect 28700 12870 28756 12908
rect 28700 12292 28756 12302
rect 28700 12198 28756 12236
rect 28364 11394 28532 11396
rect 28364 11342 28366 11394
rect 28418 11342 28532 11394
rect 28364 11340 28532 11342
rect 28588 12180 28644 12190
rect 28140 8260 28196 8270
rect 28140 8166 28196 8204
rect 28140 6804 28196 6814
rect 27692 6802 28196 6804
rect 27692 6750 28142 6802
rect 28194 6750 28196 6802
rect 27692 6748 28196 6750
rect 26572 6578 26628 6590
rect 26572 6526 26574 6578
rect 26626 6526 26628 6578
rect 26572 6132 26628 6526
rect 26908 6578 26964 6748
rect 26908 6526 26910 6578
rect 26962 6526 26964 6578
rect 26908 6514 26964 6526
rect 27468 6578 27524 6590
rect 27468 6526 27470 6578
rect 27522 6526 27524 6578
rect 26572 6066 26628 6076
rect 27020 6468 27076 6478
rect 26348 5908 26404 5918
rect 26348 5814 26404 5852
rect 26684 5796 26740 5806
rect 26684 5702 26740 5740
rect 26236 5506 26292 5516
rect 25676 5070 25678 5122
rect 25730 5070 25732 5122
rect 25676 5058 25732 5070
rect 26348 5012 26404 5022
rect 26124 5010 26404 5012
rect 26124 4958 26350 5010
rect 26402 4958 26404 5010
rect 26124 4956 26404 4958
rect 26124 4562 26180 4956
rect 26348 4946 26404 4956
rect 27020 4676 27076 6412
rect 27468 6468 27524 6526
rect 27468 6402 27524 6412
rect 27916 6578 27972 6590
rect 27916 6526 27918 6578
rect 27970 6526 27972 6578
rect 27916 6468 27972 6526
rect 27916 5460 27972 6412
rect 28140 5796 28196 6748
rect 28140 5730 28196 5740
rect 27916 5394 27972 5404
rect 28364 5236 28420 11340
rect 28476 11172 28532 11182
rect 28476 9716 28532 11116
rect 28588 10836 28644 12124
rect 28924 12178 28980 13020
rect 29260 13074 29316 15092
rect 29708 14530 29764 15092
rect 29708 14478 29710 14530
rect 29762 14478 29764 14530
rect 29708 14466 29764 14478
rect 29932 14756 29988 14766
rect 30044 14756 30100 15092
rect 30192 14924 30456 14934
rect 30248 14868 30296 14924
rect 30352 14868 30400 14924
rect 30192 14858 30456 14868
rect 30268 14756 30324 14766
rect 30044 14700 30268 14756
rect 29484 14308 29540 14318
rect 29484 13636 29540 14252
rect 29932 13972 29988 14700
rect 30268 14690 30324 14700
rect 30828 14644 30884 14654
rect 30268 14532 30324 14542
rect 30268 14438 30324 14476
rect 30044 13972 30100 13982
rect 29932 13916 30044 13972
rect 30044 13878 30100 13916
rect 30492 13860 30548 13870
rect 30492 13858 30660 13860
rect 30492 13806 30494 13858
rect 30546 13806 30660 13858
rect 30492 13804 30660 13806
rect 30492 13794 30548 13804
rect 29484 13542 29540 13580
rect 30192 13356 30456 13366
rect 30248 13300 30296 13356
rect 30352 13300 30400 13356
rect 30192 13290 30456 13300
rect 29260 13022 29262 13074
rect 29314 13022 29316 13074
rect 29260 12964 29316 13022
rect 29260 12898 29316 12908
rect 28924 12126 28926 12178
rect 28978 12126 28980 12178
rect 28924 12114 28980 12126
rect 29036 12852 29092 12862
rect 29036 11956 29092 12796
rect 29036 11890 29092 11900
rect 29260 11954 29316 11966
rect 29260 11902 29262 11954
rect 29314 11902 29316 11954
rect 29260 11620 29316 11902
rect 30192 11788 30456 11798
rect 30248 11732 30296 11788
rect 30352 11732 30400 11788
rect 30192 11722 30456 11732
rect 29260 11554 29316 11564
rect 29260 11396 29316 11406
rect 30604 11396 30660 13804
rect 30716 13636 30772 13646
rect 30716 13522 30772 13580
rect 30716 13470 30718 13522
rect 30770 13470 30772 13522
rect 30716 13458 30772 13470
rect 30828 12404 30884 14588
rect 30828 12338 30884 12348
rect 30716 11396 30772 11406
rect 30604 11394 30772 11396
rect 30604 11342 30718 11394
rect 30770 11342 30772 11394
rect 30604 11340 30772 11342
rect 29260 11302 29316 11340
rect 30716 11284 30772 11340
rect 30716 11218 30772 11228
rect 29708 11170 29764 11182
rect 29708 11118 29710 11170
rect 29762 11118 29764 11170
rect 29708 11060 29764 11118
rect 30156 11172 30212 11182
rect 30492 11172 30548 11182
rect 30212 11170 30548 11172
rect 30212 11118 30494 11170
rect 30546 11118 30548 11170
rect 30212 11116 30548 11118
rect 30156 11078 30212 11116
rect 30492 11106 30548 11116
rect 30604 11170 30660 11182
rect 30604 11118 30606 11170
rect 30658 11118 30660 11170
rect 29708 10994 29764 11004
rect 28588 10770 28644 10780
rect 30380 10724 30436 10734
rect 30604 10724 30660 11118
rect 30380 10722 30660 10724
rect 30380 10670 30382 10722
rect 30434 10670 30660 10722
rect 30380 10668 30660 10670
rect 30380 10658 30436 10668
rect 28588 10612 28644 10622
rect 28588 10518 28644 10556
rect 29708 10610 29764 10622
rect 29708 10558 29710 10610
rect 29762 10558 29764 10610
rect 28476 9650 28532 9660
rect 29036 8932 29092 8942
rect 29036 8838 29092 8876
rect 29708 8258 29764 10558
rect 30192 10220 30456 10230
rect 30248 10164 30296 10220
rect 30352 10164 30400 10220
rect 30192 10154 30456 10164
rect 30492 10052 30548 10062
rect 30492 9716 30548 9996
rect 30492 9650 30548 9660
rect 30940 9268 30996 16492
rect 31052 16324 31108 16334
rect 31052 16098 31108 16268
rect 31052 16046 31054 16098
rect 31106 16046 31108 16098
rect 31052 16034 31108 16046
rect 31388 16100 31444 16110
rect 31164 15988 31220 15998
rect 31164 15876 31220 15932
rect 31388 15986 31444 16044
rect 31388 15934 31390 15986
rect 31442 15934 31444 15986
rect 31388 15922 31444 15934
rect 31052 15820 31220 15876
rect 31052 13748 31108 15820
rect 31500 15764 31556 18396
rect 31612 17666 31668 17678
rect 31612 17614 31614 17666
rect 31666 17614 31668 17666
rect 31612 15988 31668 17614
rect 32060 17108 32116 21644
rect 32284 21474 32340 21486
rect 32284 21422 32286 21474
rect 32338 21422 32340 21474
rect 32284 21364 32340 21422
rect 32284 21298 32340 21308
rect 32732 20916 32788 21644
rect 33180 21476 33236 21486
rect 33180 21382 33236 21420
rect 32732 20850 32788 20860
rect 32396 20802 32452 20814
rect 32396 20750 32398 20802
rect 32450 20750 32452 20802
rect 32172 20132 32228 20142
rect 32172 20038 32228 20076
rect 32396 19236 32452 20750
rect 33292 20692 33348 20702
rect 33292 20598 33348 20636
rect 32844 20244 32900 20254
rect 32508 20132 32564 20142
rect 32508 20038 32564 20076
rect 32396 19170 32452 19180
rect 32620 17668 32676 17678
rect 31948 17052 32116 17108
rect 32172 17442 32228 17454
rect 32172 17390 32174 17442
rect 32226 17390 32228 17442
rect 31836 16996 31892 17006
rect 31836 16212 31892 16940
rect 31948 16324 32004 17052
rect 32060 16884 32116 16894
rect 32060 16770 32116 16828
rect 32060 16718 32062 16770
rect 32114 16718 32116 16770
rect 32060 16706 32116 16718
rect 32172 16772 32228 17390
rect 32172 16706 32228 16716
rect 32508 16882 32564 16894
rect 32508 16830 32510 16882
rect 32562 16830 32564 16882
rect 32284 16658 32340 16670
rect 32284 16606 32286 16658
rect 32338 16606 32340 16658
rect 32284 16324 32340 16606
rect 31948 16268 32228 16324
rect 31836 16156 32004 16212
rect 31612 15922 31668 15932
rect 31724 15986 31780 15998
rect 31724 15934 31726 15986
rect 31778 15934 31780 15986
rect 31388 15708 31556 15764
rect 31724 15764 31780 15934
rect 31276 15652 31332 15662
rect 31276 15538 31332 15596
rect 31276 15486 31278 15538
rect 31330 15486 31332 15538
rect 31276 15474 31332 15486
rect 31276 14530 31332 14542
rect 31276 14478 31278 14530
rect 31330 14478 31332 14530
rect 31052 13682 31108 13692
rect 31164 14084 31220 14094
rect 31164 13636 31220 14028
rect 31164 13570 31220 13580
rect 31276 13186 31332 14478
rect 31388 13860 31444 15708
rect 31724 15698 31780 15708
rect 31836 15988 31892 15998
rect 31724 15316 31780 15326
rect 31724 15222 31780 15260
rect 31388 13794 31444 13804
rect 31836 13858 31892 15932
rect 31836 13806 31838 13858
rect 31890 13806 31892 13858
rect 31836 13794 31892 13806
rect 31276 13134 31278 13186
rect 31330 13134 31332 13186
rect 31276 13122 31332 13134
rect 31500 13748 31556 13758
rect 31388 12850 31444 12862
rect 31388 12798 31390 12850
rect 31442 12798 31444 12850
rect 31388 12292 31444 12798
rect 31500 12404 31556 13692
rect 31836 13524 31892 13534
rect 31612 13188 31668 13198
rect 31612 12852 31668 13132
rect 31836 13186 31892 13468
rect 31836 13134 31838 13186
rect 31890 13134 31892 13186
rect 31836 13122 31892 13134
rect 31724 12852 31780 12862
rect 31612 12850 31780 12852
rect 31612 12798 31726 12850
rect 31778 12798 31780 12850
rect 31612 12796 31780 12798
rect 31724 12628 31780 12796
rect 31948 12740 32004 16156
rect 32060 15876 32116 15886
rect 32060 15426 32116 15820
rect 32060 15374 32062 15426
rect 32114 15374 32116 15426
rect 32060 15362 32116 15374
rect 32172 15316 32228 16268
rect 32284 16258 32340 16268
rect 32508 16098 32564 16830
rect 32508 16046 32510 16098
rect 32562 16046 32564 16098
rect 32284 15988 32340 15998
rect 32508 15988 32564 16046
rect 32284 15986 32452 15988
rect 32284 15934 32286 15986
rect 32338 15934 32452 15986
rect 32284 15932 32452 15934
rect 32284 15922 32340 15932
rect 32284 15540 32340 15550
rect 32284 15446 32340 15484
rect 32172 15260 32340 15316
rect 32172 15092 32228 15102
rect 32060 15090 32228 15092
rect 32060 15038 32174 15090
rect 32226 15038 32228 15090
rect 32060 15036 32228 15038
rect 32060 13746 32116 15036
rect 32172 15026 32228 15036
rect 32060 13694 32062 13746
rect 32114 13694 32116 13746
rect 32060 13682 32116 13694
rect 32284 13300 32340 15260
rect 32396 14530 32452 15932
rect 32508 15922 32564 15932
rect 32396 14478 32398 14530
rect 32450 14478 32452 14530
rect 32396 14466 32452 14478
rect 32508 15426 32564 15438
rect 32508 15374 32510 15426
rect 32562 15374 32564 15426
rect 31948 12674 32004 12684
rect 32060 13244 32340 13300
rect 32396 14196 32452 14206
rect 32060 12628 32116 13244
rect 32284 12964 32340 12974
rect 32396 12964 32452 14140
rect 32508 13748 32564 15374
rect 32508 13682 32564 13692
rect 32620 12964 32676 17612
rect 32732 16884 32788 16894
rect 32732 16322 32788 16828
rect 32732 16270 32734 16322
rect 32786 16270 32788 16322
rect 32732 14642 32788 16270
rect 32732 14590 32734 14642
rect 32786 14590 32788 14642
rect 32732 14578 32788 14590
rect 32844 13188 32900 20188
rect 33404 20132 33460 23324
rect 33516 23314 33572 23324
rect 33740 23314 33796 23326
rect 33628 22370 33684 22382
rect 33628 22318 33630 22370
rect 33682 22318 33684 22370
rect 33404 20066 33460 20076
rect 33516 21812 33572 21822
rect 33628 21812 33684 22318
rect 33572 21756 33684 21812
rect 33516 20130 33572 21756
rect 33516 20078 33518 20130
rect 33570 20078 33572 20130
rect 33516 20066 33572 20078
rect 33740 20802 33796 20814
rect 33740 20750 33742 20802
rect 33794 20750 33796 20802
rect 33740 20130 33796 20750
rect 34076 20244 34132 23886
rect 34188 23154 34244 24108
rect 34300 24162 34356 27020
rect 34412 28082 34468 28252
rect 34412 28030 34414 28082
rect 34466 28030 34468 28082
rect 34412 25620 34468 28030
rect 34524 28252 34692 28308
rect 34524 27860 34580 28252
rect 34860 28196 34916 28478
rect 34636 28140 34916 28196
rect 34636 28082 34692 28140
rect 34972 28084 35028 29260
rect 35084 28308 35140 29372
rect 35196 28868 35252 28878
rect 35196 28774 35252 28812
rect 35420 28868 35476 29486
rect 35532 29540 35588 29550
rect 35532 29446 35588 29484
rect 35868 29426 35924 29438
rect 35868 29374 35870 29426
rect 35922 29374 35924 29426
rect 35756 29316 35812 29326
rect 35756 29222 35812 29260
rect 35420 28802 35476 28812
rect 35308 28644 35364 28654
rect 35308 28550 35364 28588
rect 35868 28642 35924 29374
rect 36092 29092 36148 29596
rect 36428 29538 36484 30156
rect 36428 29486 36430 29538
rect 36482 29486 36484 29538
rect 36428 29474 36484 29486
rect 36204 29428 36260 29438
rect 36204 29334 36260 29372
rect 35868 28590 35870 28642
rect 35922 28590 35924 28642
rect 35084 28242 35140 28252
rect 35644 28532 35700 28542
rect 34636 28030 34638 28082
rect 34690 28030 34692 28082
rect 34636 28018 34692 28030
rect 34860 28028 35028 28084
rect 35420 28084 35476 28094
rect 34860 27972 34916 28028
rect 34860 27878 34916 27916
rect 34972 27860 35028 27870
rect 34524 27804 34804 27860
rect 34748 27748 34804 27804
rect 34972 27766 35028 27804
rect 35420 27748 35476 28028
rect 34748 27692 34916 27748
rect 34412 25554 34468 25564
rect 34524 27636 34580 27646
rect 34300 24110 34302 24162
rect 34354 24110 34356 24162
rect 34300 24098 34356 24110
rect 34412 24724 34468 24734
rect 34412 23156 34468 24668
rect 34524 23940 34580 27580
rect 34524 23874 34580 23884
rect 34748 27076 34804 27086
rect 34188 23102 34190 23154
rect 34242 23102 34244 23154
rect 34188 23090 34244 23102
rect 34300 23100 34468 23156
rect 34636 23156 34692 23166
rect 34188 22932 34244 22942
rect 34188 21140 34244 22876
rect 34300 21476 34356 23100
rect 34636 23062 34692 23100
rect 34412 22932 34468 22942
rect 34412 22838 34468 22876
rect 34300 21382 34356 21420
rect 34636 22260 34692 22270
rect 34636 21588 34692 22204
rect 34748 21812 34804 27020
rect 34860 25506 34916 27692
rect 35420 27682 35476 27692
rect 35084 27188 35140 27198
rect 35084 26908 35140 27132
rect 35532 26962 35588 26974
rect 35532 26910 35534 26962
rect 35586 26910 35588 26962
rect 35084 26852 35252 26908
rect 35196 25732 35252 26852
rect 35532 26740 35588 26910
rect 35532 26674 35588 26684
rect 35308 26628 35364 26638
rect 35308 26290 35364 26572
rect 35308 26238 35310 26290
rect 35362 26238 35364 26290
rect 35308 26226 35364 26238
rect 35196 25618 35252 25676
rect 35196 25566 35198 25618
rect 35250 25566 35252 25618
rect 35196 25554 35252 25566
rect 35532 25620 35588 25630
rect 34860 25454 34862 25506
rect 34914 25454 34916 25506
rect 34860 23492 34916 25454
rect 35308 25060 35364 25070
rect 35308 23828 35364 25004
rect 35532 24052 35588 25564
rect 35644 24500 35700 28476
rect 35868 27412 35924 28590
rect 35868 27346 35924 27356
rect 35980 29036 36148 29092
rect 36540 29202 36596 29214
rect 36540 29150 36542 29202
rect 36594 29150 36596 29202
rect 35756 27300 35812 27310
rect 35756 26964 35812 27244
rect 35756 26898 35812 26908
rect 35756 25620 35812 25630
rect 35756 25526 35812 25564
rect 35644 24444 35812 24500
rect 35532 23938 35588 23996
rect 35532 23886 35534 23938
rect 35586 23886 35588 23938
rect 35532 23874 35588 23886
rect 35308 23826 35476 23828
rect 35308 23774 35310 23826
rect 35362 23774 35476 23826
rect 35308 23772 35476 23774
rect 35308 23762 35364 23772
rect 35420 23716 35476 23772
rect 35420 23660 35588 23716
rect 34860 23426 34916 23436
rect 35420 23156 35476 23166
rect 35308 23042 35364 23054
rect 35308 22990 35310 23042
rect 35362 22990 35364 23042
rect 35308 21812 35364 22990
rect 35420 22370 35476 23100
rect 35532 23154 35588 23660
rect 35532 23102 35534 23154
rect 35586 23102 35588 23154
rect 35532 23090 35588 23102
rect 35756 22482 35812 24444
rect 35980 24164 36036 29036
rect 36092 28868 36148 28878
rect 36092 28642 36148 28812
rect 36092 28590 36094 28642
rect 36146 28590 36148 28642
rect 36092 28578 36148 28590
rect 36428 28530 36484 28542
rect 36428 28478 36430 28530
rect 36482 28478 36484 28530
rect 36092 28420 36148 28430
rect 36316 28420 36372 28430
rect 36092 27074 36148 28364
rect 36092 27022 36094 27074
rect 36146 27022 36148 27074
rect 36092 24498 36148 27022
rect 36204 28418 36372 28420
rect 36204 28366 36318 28418
rect 36370 28366 36372 28418
rect 36204 28364 36372 28366
rect 36204 26908 36260 28364
rect 36316 28354 36372 28364
rect 36428 28420 36484 28478
rect 36428 28354 36484 28364
rect 36540 26908 36596 29150
rect 36652 28644 36708 30380
rect 36652 28578 36708 28588
rect 36764 28084 36820 35196
rect 36876 35140 36932 35646
rect 37548 35588 37604 35598
rect 36876 35074 36932 35084
rect 36988 35476 37044 35486
rect 36876 34356 36932 34366
rect 36876 33684 36932 34300
rect 36988 34130 37044 35420
rect 36988 34078 36990 34130
rect 37042 34078 37044 34130
rect 36988 34066 37044 34078
rect 37100 34916 37156 34926
rect 37324 34916 37380 34926
rect 36876 33628 37044 33684
rect 36876 33012 36932 33022
rect 36876 32564 36932 32956
rect 36988 32786 37044 33628
rect 37100 33570 37156 34860
rect 37212 34914 37380 34916
rect 37212 34862 37326 34914
rect 37378 34862 37380 34914
rect 37212 34860 37380 34862
rect 37212 33684 37268 34860
rect 37324 34850 37380 34860
rect 37436 34020 37492 34030
rect 37436 33926 37492 33964
rect 37212 33628 37380 33684
rect 37100 33518 37102 33570
rect 37154 33518 37156 33570
rect 37100 33506 37156 33518
rect 37212 33460 37268 33470
rect 37212 33346 37268 33404
rect 37212 33294 37214 33346
rect 37266 33294 37268 33346
rect 37212 33282 37268 33294
rect 37324 33236 37380 33628
rect 37548 33348 37604 35532
rect 37660 34916 37716 35756
rect 38220 35746 38276 35756
rect 38780 35698 38836 35710
rect 38780 35646 38782 35698
rect 38834 35646 38836 35698
rect 37772 35588 37828 35598
rect 37772 35494 37828 35532
rect 37884 35474 37940 35486
rect 37884 35422 37886 35474
rect 37938 35422 37940 35474
rect 37884 35252 37940 35422
rect 37884 35186 37940 35196
rect 38444 35252 38500 35262
rect 38780 35252 38836 35646
rect 38500 35196 38612 35252
rect 38444 35186 38500 35196
rect 37772 34916 37828 34926
rect 37660 34914 37828 34916
rect 37660 34862 37774 34914
rect 37826 34862 37828 34914
rect 37660 34860 37828 34862
rect 37772 34850 37828 34860
rect 38444 34916 38500 34926
rect 38444 34822 38500 34860
rect 38556 34802 38612 35196
rect 38556 34750 38558 34802
rect 38610 34750 38612 34802
rect 38556 34738 38612 34750
rect 38780 34356 38836 35196
rect 39116 35586 39172 35598
rect 39116 35534 39118 35586
rect 39170 35534 39172 35586
rect 38556 34300 38836 34356
rect 38892 35140 38948 35150
rect 37548 33282 37604 33292
rect 37772 33460 37828 33470
rect 37772 33346 37828 33404
rect 37772 33294 37774 33346
rect 37826 33294 37828 33346
rect 37772 33282 37828 33294
rect 38332 33458 38388 33470
rect 38332 33406 38334 33458
rect 38386 33406 38388 33458
rect 36988 32734 36990 32786
rect 37042 32734 37044 32786
rect 36988 32722 37044 32734
rect 37100 33124 37156 33134
rect 37324 33124 37380 33180
rect 37996 33236 38052 33246
rect 37996 33142 38052 33180
rect 37100 33122 37380 33124
rect 37100 33070 37102 33122
rect 37154 33070 37380 33122
rect 37100 33068 37380 33070
rect 36876 32508 37044 32564
rect 36988 31780 37044 32508
rect 37100 32002 37156 33068
rect 37212 32900 37268 32910
rect 37212 32674 37268 32844
rect 37212 32622 37214 32674
rect 37266 32622 37268 32674
rect 37212 32610 37268 32622
rect 37324 32564 37380 32574
rect 37100 31950 37102 32002
rect 37154 31950 37156 32002
rect 37100 31938 37156 31950
rect 37212 32452 37268 32462
rect 37212 31780 37268 32396
rect 37324 31890 37380 32508
rect 37436 32562 37492 32574
rect 37436 32510 37438 32562
rect 37490 32510 37492 32562
rect 37436 32004 37492 32510
rect 37884 32562 37940 32574
rect 37884 32510 37886 32562
rect 37938 32510 37940 32562
rect 37548 32452 37604 32462
rect 37884 32452 37940 32510
rect 37548 32450 37940 32452
rect 37548 32398 37550 32450
rect 37602 32398 37940 32450
rect 37548 32396 37940 32398
rect 37548 32386 37604 32396
rect 37436 31938 37492 31948
rect 37324 31838 37326 31890
rect 37378 31838 37380 31890
rect 37324 31826 37380 31838
rect 36988 31714 37044 31724
rect 37100 31724 37268 31780
rect 37548 31780 37604 31790
rect 37548 31778 37716 31780
rect 37548 31726 37550 31778
rect 37602 31726 37716 31778
rect 37548 31724 37716 31726
rect 36988 31220 37044 31230
rect 36988 31126 37044 31164
rect 36988 30882 37044 30894
rect 36988 30830 36990 30882
rect 37042 30830 37044 30882
rect 36988 29540 37044 30830
rect 37100 30324 37156 31724
rect 37548 31714 37604 31724
rect 37436 31556 37492 31566
rect 37436 31554 37604 31556
rect 37436 31502 37438 31554
rect 37490 31502 37604 31554
rect 37436 31500 37604 31502
rect 37436 31490 37492 31500
rect 37212 30994 37268 31006
rect 37212 30942 37214 30994
rect 37266 30942 37268 30994
rect 37212 30884 37268 30942
rect 37436 30996 37492 31006
rect 37436 30902 37492 30940
rect 37212 30818 37268 30828
rect 37100 30268 37268 30324
rect 36988 29474 37044 29484
rect 36764 28018 36820 28028
rect 36876 29426 36932 29438
rect 36876 29374 36878 29426
rect 36930 29374 36932 29426
rect 36204 26852 36372 26908
rect 36540 26852 36820 26908
rect 36316 26740 36372 26852
rect 36316 26674 36372 26684
rect 36652 26516 36708 26526
rect 36652 26422 36708 26460
rect 36764 26402 36820 26852
rect 36764 26350 36766 26402
rect 36818 26350 36820 26402
rect 36764 26338 36820 26350
rect 36876 25172 36932 29374
rect 36988 29316 37044 29326
rect 36988 28642 37044 29260
rect 36988 28590 36990 28642
rect 37042 28590 37044 28642
rect 36988 28578 37044 28590
rect 37100 28980 37156 28990
rect 37100 27972 37156 28924
rect 37100 27906 37156 27916
rect 37100 27746 37156 27758
rect 37100 27694 37102 27746
rect 37154 27694 37156 27746
rect 37100 27412 37156 27694
rect 37100 27346 37156 27356
rect 37212 26908 37268 30268
rect 37436 30212 37492 30222
rect 37548 30212 37604 31500
rect 37660 30436 37716 31724
rect 38332 31778 38388 33406
rect 38444 33124 38500 33134
rect 38444 32452 38500 33068
rect 38556 32900 38612 34300
rect 38556 32834 38612 32844
rect 38892 33906 38948 35084
rect 39116 35140 39172 35534
rect 39228 35364 39284 36430
rect 39228 35298 39284 35308
rect 39116 35074 39172 35084
rect 39340 34916 39396 34926
rect 38892 33854 38894 33906
rect 38946 33854 38948 33906
rect 38892 33348 38948 33854
rect 38892 32674 38948 33292
rect 39004 34914 39396 34916
rect 39004 34862 39342 34914
rect 39394 34862 39396 34914
rect 39004 34860 39396 34862
rect 39004 32786 39060 34860
rect 39340 34850 39396 34860
rect 39340 34692 39396 34702
rect 39004 32734 39006 32786
rect 39058 32734 39060 32786
rect 39004 32722 39060 32734
rect 39228 34690 39396 34692
rect 39228 34638 39342 34690
rect 39394 34638 39396 34690
rect 39228 34636 39396 34638
rect 38892 32622 38894 32674
rect 38946 32622 38948 32674
rect 38892 32564 38948 32622
rect 38892 32498 38948 32508
rect 38444 32358 38500 32396
rect 39228 31890 39284 34636
rect 39340 34626 39396 34636
rect 39340 34132 39396 34142
rect 39340 32786 39396 34076
rect 39452 33348 39508 33358
rect 39452 33254 39508 33292
rect 39340 32734 39342 32786
rect 39394 32734 39396 32786
rect 39340 32722 39396 32734
rect 39452 32788 39508 32798
rect 39452 32452 39508 32732
rect 39452 32386 39508 32396
rect 39228 31838 39230 31890
rect 39282 31838 39284 31890
rect 39228 31826 39284 31838
rect 39452 31892 39508 31902
rect 38332 31726 38334 31778
rect 38386 31726 38388 31778
rect 38332 31714 38388 31726
rect 39004 31778 39060 31790
rect 39004 31726 39006 31778
rect 39058 31726 39060 31778
rect 39004 31668 39060 31726
rect 38108 31556 38164 31566
rect 38108 31554 38276 31556
rect 38108 31502 38110 31554
rect 38162 31502 38276 31554
rect 38108 31500 38276 31502
rect 38108 31490 38164 31500
rect 37660 30370 37716 30380
rect 37772 30994 37828 31006
rect 37772 30942 37774 30994
rect 37826 30942 37828 30994
rect 37492 30156 37604 30212
rect 37660 30212 37716 30222
rect 37436 30146 37492 30156
rect 37324 30100 37380 30110
rect 37324 28420 37380 30044
rect 37660 29876 37716 30156
rect 37772 30100 37828 30942
rect 37996 30994 38052 31006
rect 37996 30942 37998 30994
rect 38050 30942 38052 30994
rect 37996 30884 38052 30942
rect 37772 30034 37828 30044
rect 37884 30548 37940 30558
rect 37324 28354 37380 28364
rect 37436 29820 37716 29876
rect 37436 27860 37492 29820
rect 37884 29764 37940 30492
rect 37996 30212 38052 30828
rect 37996 30146 38052 30156
rect 38108 30994 38164 31006
rect 38108 30942 38110 30994
rect 38162 30942 38164 30994
rect 38108 30212 38164 30942
rect 38220 30996 38276 31500
rect 38220 30930 38276 30940
rect 38892 30996 38948 31006
rect 38556 30772 38612 30782
rect 38556 30770 38724 30772
rect 38556 30718 38558 30770
rect 38610 30718 38724 30770
rect 38556 30716 38724 30718
rect 38556 30706 38612 30716
rect 38108 30210 38276 30212
rect 38108 30158 38110 30210
rect 38162 30158 38276 30210
rect 38108 30156 38276 30158
rect 38108 30146 38164 30156
rect 38108 29988 38164 29998
rect 38108 29894 38164 29932
rect 37548 29708 37940 29764
rect 37548 28756 37604 29708
rect 38220 29652 38276 30156
rect 38668 30210 38724 30716
rect 38668 30158 38670 30210
rect 38722 30158 38724 30210
rect 38668 30146 38724 30158
rect 37996 29650 38276 29652
rect 37996 29598 38222 29650
rect 38274 29598 38276 29650
rect 37996 29596 38276 29598
rect 37996 29540 38052 29596
rect 38220 29586 38276 29596
rect 37660 29484 38052 29540
rect 38444 29540 38500 29550
rect 37660 29426 37716 29484
rect 38444 29446 38500 29484
rect 37660 29374 37662 29426
rect 37714 29374 37716 29426
rect 37660 29362 37716 29374
rect 38556 29428 38612 29438
rect 38668 29428 38724 29438
rect 38556 29426 38668 29428
rect 38556 29374 38558 29426
rect 38610 29374 38668 29426
rect 38556 29372 38668 29374
rect 38556 29362 38612 29372
rect 38668 29362 38724 29372
rect 38892 29426 38948 30940
rect 39004 29876 39060 31612
rect 39116 31556 39172 31566
rect 39116 30210 39172 31500
rect 39116 30158 39118 30210
rect 39170 30158 39172 30210
rect 39116 30146 39172 30158
rect 39340 31106 39396 31118
rect 39340 31054 39342 31106
rect 39394 31054 39396 31106
rect 39340 29988 39396 31054
rect 39452 30994 39508 31836
rect 39452 30942 39454 30994
rect 39506 30942 39508 30994
rect 39452 30660 39508 30942
rect 39452 30594 39508 30604
rect 39452 30322 39508 30334
rect 39452 30270 39454 30322
rect 39506 30270 39508 30322
rect 39452 30212 39508 30270
rect 39452 30146 39508 30156
rect 39340 29922 39396 29932
rect 39004 29820 39172 29876
rect 38892 29374 38894 29426
rect 38946 29374 38948 29426
rect 38444 29316 38500 29326
rect 37660 28756 37716 28766
rect 37548 28754 37716 28756
rect 37548 28702 37662 28754
rect 37714 28702 37716 28754
rect 37548 28700 37716 28702
rect 38444 28756 38500 29260
rect 38556 28756 38612 28766
rect 38444 28754 38612 28756
rect 38444 28702 38558 28754
rect 38610 28702 38612 28754
rect 38444 28700 38612 28702
rect 37436 27794 37492 27804
rect 37548 28196 37604 28206
rect 37436 27524 37492 27534
rect 37212 26852 37380 26908
rect 37212 25282 37268 25294
rect 37212 25230 37214 25282
rect 37266 25230 37268 25282
rect 36876 25116 37156 25172
rect 37100 24946 37156 25116
rect 37100 24894 37102 24946
rect 37154 24894 37156 24946
rect 37100 24882 37156 24894
rect 37212 25060 37268 25230
rect 36092 24446 36094 24498
rect 36146 24446 36148 24498
rect 36092 24434 36148 24446
rect 36316 24722 36372 24734
rect 36316 24670 36318 24722
rect 36370 24670 36372 24722
rect 36316 24500 36372 24670
rect 36316 24434 36372 24444
rect 36764 24610 36820 24622
rect 36764 24558 36766 24610
rect 36818 24558 36820 24610
rect 36316 24164 36372 24174
rect 35980 24108 36148 24164
rect 35980 23938 36036 23950
rect 35980 23886 35982 23938
rect 36034 23886 36036 23938
rect 35980 23604 36036 23886
rect 35980 23538 36036 23548
rect 35756 22430 35758 22482
rect 35810 22430 35812 22482
rect 35756 22418 35812 22430
rect 36092 23378 36148 24108
rect 36316 24070 36372 24108
rect 36540 23492 36596 23502
rect 36092 23326 36094 23378
rect 36146 23326 36148 23378
rect 35420 22318 35422 22370
rect 35474 22318 35476 22370
rect 35420 22306 35476 22318
rect 34748 21756 35140 21812
rect 34748 21588 34804 21598
rect 34636 21586 34804 21588
rect 34636 21534 34750 21586
rect 34802 21534 34804 21586
rect 34636 21532 34804 21534
rect 34188 21084 34356 21140
rect 34076 20178 34132 20188
rect 33740 20078 33742 20130
rect 33794 20078 33796 20130
rect 33180 19796 33236 19806
rect 33180 19794 33348 19796
rect 33180 19742 33182 19794
rect 33234 19742 33348 19794
rect 33180 19740 33348 19742
rect 33180 19730 33236 19740
rect 33180 19236 33236 19246
rect 33180 19142 33236 19180
rect 33292 17666 33348 19740
rect 33628 19460 33684 19470
rect 33628 19124 33684 19404
rect 33740 19346 33796 20078
rect 33964 20132 34020 20142
rect 33964 20038 34020 20076
rect 33740 19294 33742 19346
rect 33794 19294 33796 19346
rect 33740 19236 33796 19294
rect 34076 19236 34132 19246
rect 33740 19234 34244 19236
rect 33740 19182 34078 19234
rect 34130 19182 34244 19234
rect 33740 19180 34244 19182
rect 34076 19170 34132 19180
rect 33628 19068 33796 19124
rect 33516 18676 33572 18686
rect 33404 17780 33460 17790
rect 33404 17686 33460 17724
rect 33292 17614 33294 17666
rect 33346 17614 33348 17666
rect 33068 16882 33124 16894
rect 33068 16830 33070 16882
rect 33122 16830 33124 16882
rect 32956 16324 33012 16334
rect 32956 15538 33012 16268
rect 33068 16100 33124 16830
rect 33292 16884 33348 17614
rect 33516 17220 33572 18620
rect 33628 17556 33684 17566
rect 33628 17462 33684 17500
rect 33292 16818 33348 16828
rect 33404 17164 33572 17220
rect 33404 16322 33460 17164
rect 33516 16882 33572 16894
rect 33516 16830 33518 16882
rect 33570 16830 33572 16882
rect 33516 16772 33572 16830
rect 33516 16706 33572 16716
rect 33404 16270 33406 16322
rect 33458 16270 33460 16322
rect 33404 16258 33460 16270
rect 33628 16324 33684 16334
rect 33068 16034 33124 16044
rect 32956 15486 32958 15538
rect 33010 15486 33012 15538
rect 32956 15474 33012 15486
rect 33068 15764 33124 15774
rect 33068 14196 33124 15708
rect 33628 15652 33684 16268
rect 33068 14130 33124 14140
rect 33180 15426 33236 15438
rect 33180 15374 33182 15426
rect 33234 15374 33236 15426
rect 33068 13860 33124 13870
rect 33068 13766 33124 13804
rect 33180 13636 33236 15374
rect 33628 15426 33684 15596
rect 33628 15374 33630 15426
rect 33682 15374 33684 15426
rect 33628 15362 33684 15374
rect 33292 15314 33348 15326
rect 33292 15262 33294 15314
rect 33346 15262 33348 15314
rect 33292 15148 33348 15262
rect 33740 15316 33796 19068
rect 34188 18228 34244 19180
rect 34300 18452 34356 21084
rect 34636 20690 34692 21532
rect 34748 21522 34804 21532
rect 34636 20638 34638 20690
rect 34690 20638 34692 20690
rect 34524 20132 34580 20142
rect 34524 20018 34580 20076
rect 34524 19966 34526 20018
rect 34578 19966 34580 20018
rect 34524 19954 34580 19966
rect 34636 19796 34692 20638
rect 34636 19730 34692 19740
rect 34748 20914 34804 20926
rect 34748 20862 34750 20914
rect 34802 20862 34804 20914
rect 34300 18358 34356 18396
rect 34636 18450 34692 18462
rect 34636 18398 34638 18450
rect 34690 18398 34692 18450
rect 34636 18228 34692 18398
rect 34188 18172 34692 18228
rect 34748 18004 34804 20862
rect 34972 18564 35028 18574
rect 34972 18470 35028 18508
rect 34748 17892 34804 17948
rect 34300 17836 34804 17892
rect 34972 17892 35028 17902
rect 34300 17666 34356 17836
rect 34636 17668 34692 17678
rect 34300 17614 34302 17666
rect 34354 17614 34356 17666
rect 34300 17602 34356 17614
rect 34524 17612 34636 17668
rect 34188 17554 34244 17566
rect 34188 17502 34190 17554
rect 34242 17502 34244 17554
rect 34188 17220 34244 17502
rect 34188 17154 34244 17164
rect 34524 17106 34580 17612
rect 34636 17574 34692 17612
rect 34524 17054 34526 17106
rect 34578 17054 34580 17106
rect 34524 17042 34580 17054
rect 34748 17444 34804 17454
rect 34748 16994 34804 17388
rect 34748 16942 34750 16994
rect 34802 16942 34804 16994
rect 34748 16930 34804 16942
rect 34412 16772 34468 16782
rect 34412 16678 34468 16716
rect 33852 16660 33908 16670
rect 33852 15652 33908 16604
rect 34300 16324 34356 16334
rect 34300 16210 34356 16268
rect 34300 16158 34302 16210
rect 34354 16158 34356 16210
rect 34300 16146 34356 16158
rect 33852 15538 33908 15596
rect 33852 15486 33854 15538
rect 33906 15486 33908 15538
rect 33852 15474 33908 15486
rect 33964 15876 34020 15886
rect 33740 15260 33908 15316
rect 33292 15092 33796 15148
rect 33740 15090 33796 15092
rect 33740 15038 33742 15090
rect 33794 15038 33796 15090
rect 33740 15026 33796 15038
rect 33628 14530 33684 14542
rect 33628 14478 33630 14530
rect 33682 14478 33684 14530
rect 33404 14196 33460 14206
rect 33404 13970 33460 14140
rect 33404 13918 33406 13970
rect 33458 13918 33460 13970
rect 33404 13906 33460 13918
rect 33628 13972 33684 14478
rect 33628 13906 33684 13916
rect 33852 13972 33908 15260
rect 33180 13570 33236 13580
rect 33292 13746 33348 13758
rect 33292 13694 33294 13746
rect 33346 13694 33348 13746
rect 33068 13188 33124 13198
rect 32844 13186 33124 13188
rect 32844 13134 33070 13186
rect 33122 13134 33124 13186
rect 32844 13132 33124 13134
rect 33068 13122 33124 13132
rect 33292 13188 33348 13694
rect 33628 13748 33684 13758
rect 33852 13748 33908 13916
rect 33964 13858 34020 15820
rect 34524 15652 34580 15662
rect 34524 15540 34580 15596
rect 34860 15540 34916 15550
rect 34524 15538 34916 15540
rect 34524 15486 34526 15538
rect 34578 15486 34862 15538
rect 34914 15486 34916 15538
rect 34524 15484 34916 15486
rect 34524 15474 34580 15484
rect 34860 15474 34916 15484
rect 33964 13806 33966 13858
rect 34018 13806 34020 13858
rect 33964 13794 34020 13806
rect 34076 15426 34132 15438
rect 34076 15374 34078 15426
rect 34130 15374 34132 15426
rect 34076 13860 34132 15374
rect 34188 15092 34244 15102
rect 34188 14532 34244 15036
rect 34188 13970 34244 14476
rect 34636 14530 34692 14542
rect 34636 14478 34638 14530
rect 34690 14478 34692 14530
rect 34188 13918 34190 13970
rect 34242 13918 34244 13970
rect 34188 13906 34244 13918
rect 34524 14196 34580 14206
rect 34076 13794 34132 13804
rect 34412 13858 34468 13870
rect 34412 13806 34414 13858
rect 34466 13806 34468 13858
rect 33628 13746 33908 13748
rect 33628 13694 33630 13746
rect 33682 13694 33908 13746
rect 33628 13692 33908 13694
rect 33628 13682 33684 13692
rect 34076 13636 34132 13646
rect 34076 13542 34132 13580
rect 33292 13122 33348 13132
rect 32284 12962 32452 12964
rect 32284 12910 32286 12962
rect 32338 12910 32452 12962
rect 32284 12908 32452 12910
rect 32508 12908 32676 12964
rect 32732 13074 32788 13086
rect 32732 13022 32734 13074
rect 32786 13022 32788 13074
rect 32732 12964 32788 13022
rect 32060 12572 32228 12628
rect 31724 12562 31780 12572
rect 32060 12404 32116 12414
rect 31500 12402 32116 12404
rect 31500 12350 32062 12402
rect 32114 12350 32116 12402
rect 31500 12348 32116 12350
rect 32060 12338 32116 12348
rect 31388 12226 31444 12236
rect 31948 11954 32004 11966
rect 31948 11902 31950 11954
rect 32002 11902 32004 11954
rect 31948 11506 32004 11902
rect 31948 11454 31950 11506
rect 32002 11454 32004 11506
rect 31948 11442 32004 11454
rect 31164 11394 31220 11406
rect 31164 11342 31166 11394
rect 31218 11342 31220 11394
rect 31164 9826 31220 11342
rect 31836 11394 31892 11406
rect 31836 11342 31838 11394
rect 31890 11342 31892 11394
rect 31724 11284 31780 11294
rect 31836 11284 31892 11342
rect 31780 11228 31892 11284
rect 31724 11218 31780 11228
rect 32172 10052 32228 12572
rect 31948 9996 32228 10052
rect 31948 9940 32004 9996
rect 31164 9774 31166 9826
rect 31218 9774 31220 9826
rect 31164 9762 31220 9774
rect 31388 9938 32004 9940
rect 31388 9886 31950 9938
rect 32002 9886 32004 9938
rect 31388 9884 32004 9886
rect 30716 9212 30996 9268
rect 31388 9714 31444 9884
rect 31948 9874 32004 9884
rect 31388 9662 31390 9714
rect 31442 9662 31444 9714
rect 30492 9156 30548 9166
rect 30492 9154 30660 9156
rect 30492 9102 30494 9154
rect 30546 9102 30660 9154
rect 30492 9100 30660 9102
rect 30492 9090 30548 9100
rect 30192 8652 30456 8662
rect 30248 8596 30296 8652
rect 30352 8596 30400 8652
rect 30192 8586 30456 8596
rect 30380 8372 30436 8382
rect 30604 8372 30660 9100
rect 30380 8370 30660 8372
rect 30380 8318 30382 8370
rect 30434 8318 30660 8370
rect 30380 8316 30660 8318
rect 30380 8306 30436 8316
rect 29708 8206 29710 8258
rect 29762 8206 29764 8258
rect 29484 6804 29540 6814
rect 28476 6466 28532 6478
rect 28476 6414 28478 6466
rect 28530 6414 28532 6466
rect 28476 5684 28532 6414
rect 29372 6468 29428 6478
rect 28812 5796 28868 5806
rect 28812 5794 29204 5796
rect 28812 5742 28814 5794
rect 28866 5742 29204 5794
rect 28812 5740 29204 5742
rect 28812 5730 28868 5740
rect 28476 5618 28532 5628
rect 28476 5236 28532 5246
rect 27020 4610 27076 4620
rect 27244 5234 28532 5236
rect 27244 5182 28478 5234
rect 28530 5182 28532 5234
rect 27244 5180 28532 5182
rect 26124 4510 26126 4562
rect 26178 4510 26180 4562
rect 26124 4498 26180 4510
rect 25788 4452 25844 4462
rect 25452 4340 25508 4350
rect 25452 4246 25508 4284
rect 25788 4228 25844 4396
rect 26460 4340 26516 4350
rect 26908 4340 26964 4350
rect 26460 4338 26964 4340
rect 26460 4286 26462 4338
rect 26514 4286 26910 4338
rect 26962 4286 26964 4338
rect 26460 4284 26964 4286
rect 26460 4274 26516 4284
rect 26908 4274 26964 4284
rect 27244 4338 27300 5180
rect 28476 5170 28532 5180
rect 28700 5012 28756 5022
rect 27804 4676 27860 4686
rect 27804 4450 27860 4620
rect 27804 4398 27806 4450
rect 27858 4398 27860 4450
rect 27804 4386 27860 4398
rect 27244 4286 27246 4338
rect 27298 4286 27300 4338
rect 27244 4274 27300 4286
rect 28028 4340 28084 4350
rect 28028 4246 28084 4284
rect 25788 4162 25844 4172
rect 27916 3444 27972 3454
rect 28364 3444 28420 3454
rect 25004 2482 25060 2492
rect 27804 3442 28420 3444
rect 27804 3390 27918 3442
rect 27970 3390 28366 3442
rect 28418 3390 28420 3442
rect 27804 3388 28420 3390
rect 23772 2156 24164 2212
rect 23772 800 23828 2156
rect 27804 800 27860 3388
rect 27916 3378 27972 3388
rect 28364 3378 28420 3388
rect 28700 3442 28756 4956
rect 29148 5010 29204 5740
rect 29148 4958 29150 5010
rect 29202 4958 29204 5010
rect 29148 4946 29204 4958
rect 28700 3390 28702 3442
rect 28754 3390 28756 3442
rect 28700 3378 28756 3390
rect 29372 2660 29428 6412
rect 29484 5906 29540 6748
rect 29484 5854 29486 5906
rect 29538 5854 29540 5906
rect 29484 5842 29540 5854
rect 29484 5684 29540 5694
rect 29484 5122 29540 5628
rect 29484 5070 29486 5122
rect 29538 5070 29540 5122
rect 29484 5058 29540 5070
rect 29708 5124 29764 8206
rect 30192 7084 30456 7094
rect 30248 7028 30296 7084
rect 30352 7028 30400 7084
rect 30192 7018 30456 7028
rect 30192 5516 30456 5526
rect 30248 5460 30296 5516
rect 30352 5460 30400 5516
rect 30192 5450 30456 5460
rect 29708 4338 29764 5068
rect 30268 5012 30324 5022
rect 30716 5012 30772 9212
rect 30828 9044 30884 9054
rect 30828 9042 31108 9044
rect 30828 8990 30830 9042
rect 30882 8990 31108 9042
rect 30828 8988 31108 8990
rect 30828 8978 30884 8988
rect 31052 7698 31108 8988
rect 31052 7646 31054 7698
rect 31106 7646 31108 7698
rect 31052 7634 31108 7646
rect 31388 8596 31444 9662
rect 31500 9716 31556 9726
rect 31500 9622 31556 9660
rect 31388 7474 31444 8540
rect 32284 8428 32340 12908
rect 32396 12740 32452 12750
rect 32508 12740 32564 12908
rect 32732 12898 32788 12908
rect 32844 12964 32900 12974
rect 32844 12962 33012 12964
rect 32844 12910 32846 12962
rect 32898 12910 33012 12962
rect 32844 12908 33012 12910
rect 32844 12898 32900 12908
rect 32396 12738 32564 12740
rect 32396 12686 32398 12738
rect 32450 12686 32564 12738
rect 32396 12684 32564 12686
rect 32620 12738 32676 12750
rect 32620 12686 32622 12738
rect 32674 12686 32676 12738
rect 32396 12068 32452 12684
rect 32508 12068 32564 12078
rect 32396 12066 32564 12068
rect 32396 12014 32510 12066
rect 32562 12014 32564 12066
rect 32396 12012 32564 12014
rect 32508 11172 32564 12012
rect 32508 11106 32564 11116
rect 32620 11954 32676 12686
rect 32956 12740 33012 12908
rect 32620 11902 32622 11954
rect 32674 11902 32676 11954
rect 32508 10500 32564 10510
rect 32620 10500 32676 11902
rect 32508 10498 32676 10500
rect 32508 10446 32510 10498
rect 32562 10446 32676 10498
rect 32508 10444 32676 10446
rect 32732 12628 32788 12638
rect 32508 10434 32564 10444
rect 32396 10052 32452 10062
rect 32396 9716 32452 9996
rect 32396 9622 32452 9660
rect 32508 8428 32564 8438
rect 32284 8426 32564 8428
rect 32284 8374 32510 8426
rect 32562 8374 32564 8426
rect 32284 8372 32564 8374
rect 31388 7422 31390 7474
rect 31442 7422 31444 7474
rect 31388 7410 31444 7422
rect 31724 7586 31780 7598
rect 31724 7534 31726 7586
rect 31778 7534 31780 7586
rect 31724 7028 31780 7534
rect 32172 7588 32228 7598
rect 32284 7588 32340 8372
rect 32508 8362 32564 8372
rect 32732 8036 32788 12572
rect 32956 11956 33012 12684
rect 33292 12962 33348 12974
rect 33292 12910 33294 12962
rect 33346 12910 33348 12962
rect 33292 12628 33348 12910
rect 33740 12964 33796 12974
rect 33740 12870 33796 12908
rect 33292 12572 33684 12628
rect 33516 12404 33572 12414
rect 33292 12292 33348 12302
rect 33068 11956 33124 11966
rect 32956 11900 33068 11956
rect 32956 11172 33012 11900
rect 33068 11890 33124 11900
rect 33180 11172 33236 11182
rect 32956 11170 33236 11172
rect 32956 11118 33182 11170
rect 33234 11118 33236 11170
rect 32956 11116 33236 11118
rect 33180 11106 33236 11116
rect 32172 7586 32340 7588
rect 32172 7534 32174 7586
rect 32226 7534 32340 7586
rect 32172 7532 32340 7534
rect 32396 7980 32788 8036
rect 32956 9826 33012 9838
rect 32956 9774 32958 9826
rect 33010 9774 33012 9826
rect 32956 8484 33012 9774
rect 32172 7522 32228 7532
rect 31724 6962 31780 6972
rect 32172 6018 32228 6030
rect 32172 5966 32174 6018
rect 32226 5966 32228 6018
rect 31948 5124 32004 5134
rect 32172 5124 32228 5966
rect 32004 5068 32228 5124
rect 31948 5030 32004 5068
rect 30324 4956 30772 5012
rect 31612 5012 31668 5022
rect 30268 4946 30324 4956
rect 31612 4918 31668 4956
rect 31276 4900 31332 4910
rect 30380 4898 31332 4900
rect 30380 4846 31278 4898
rect 31330 4846 31332 4898
rect 30380 4844 31332 4846
rect 30380 4450 30436 4844
rect 31276 4834 31332 4844
rect 30380 4398 30382 4450
rect 30434 4398 30436 4450
rect 30380 4386 30436 4398
rect 29708 4286 29710 4338
rect 29762 4286 29764 4338
rect 29708 4274 29764 4286
rect 32284 4340 32340 4350
rect 30192 3948 30456 3958
rect 30248 3892 30296 3948
rect 30352 3892 30400 3948
rect 30192 3882 30456 3892
rect 31724 3444 31780 3454
rect 32172 3444 32228 3454
rect 31724 3442 32228 3444
rect 31724 3390 31726 3442
rect 31778 3390 32174 3442
rect 32226 3390 32228 3442
rect 31724 3388 32228 3390
rect 31724 3378 31780 3388
rect 29372 2594 29428 2604
rect 31836 800 31892 3388
rect 32172 3378 32228 3388
rect 32284 2884 32340 4284
rect 32396 4228 32452 7980
rect 32956 7812 33012 8428
rect 32508 7756 33012 7812
rect 33180 8596 33236 8606
rect 32508 6018 32564 7756
rect 33180 7698 33236 8540
rect 33180 7646 33182 7698
rect 33234 7646 33236 7698
rect 33180 7634 33236 7646
rect 32620 7028 32676 7038
rect 32620 6690 32676 6972
rect 32620 6638 32622 6690
rect 32674 6638 32676 6690
rect 32620 6626 32676 6638
rect 33292 6356 33348 12236
rect 33516 11788 33572 12348
rect 33628 12402 33684 12572
rect 33628 12350 33630 12402
rect 33682 12350 33684 12402
rect 33628 12338 33684 12350
rect 33852 12404 33908 12414
rect 33852 12310 33908 12348
rect 33740 12180 33796 12190
rect 34412 12180 34468 13806
rect 34524 12850 34580 14140
rect 34636 13524 34692 14478
rect 34860 13972 34916 13982
rect 34860 13878 34916 13916
rect 34636 13458 34692 13468
rect 34748 13748 34804 13758
rect 34748 13076 34804 13692
rect 34972 13748 35028 17836
rect 34972 13682 35028 13692
rect 34748 13020 35028 13076
rect 34636 12964 34692 12974
rect 34636 12870 34692 12908
rect 34972 12962 35028 13020
rect 34972 12910 34974 12962
rect 35026 12910 35028 12962
rect 34524 12798 34526 12850
rect 34578 12798 34580 12850
rect 34524 12786 34580 12798
rect 34972 12516 35028 12910
rect 34636 12460 35028 12516
rect 34524 12404 34580 12414
rect 34524 12310 34580 12348
rect 33404 11732 33572 11788
rect 33628 12178 34468 12180
rect 33628 12126 33742 12178
rect 33794 12126 34468 12178
rect 33628 12124 34468 12126
rect 33404 11666 33460 11676
rect 33628 7364 33684 12124
rect 33740 12114 33796 12124
rect 34188 11732 34244 11742
rect 34188 11506 34244 11676
rect 34188 11454 34190 11506
rect 34242 11454 34244 11506
rect 34188 11284 34244 11454
rect 34188 11218 34244 11228
rect 33964 10724 34020 10734
rect 33740 10722 34020 10724
rect 33740 10670 33966 10722
rect 34018 10670 34020 10722
rect 33740 10668 34020 10670
rect 33740 9938 33796 10668
rect 33964 10658 34020 10668
rect 34300 10612 34356 10622
rect 34300 10610 34580 10612
rect 34300 10558 34302 10610
rect 34354 10558 34580 10610
rect 34300 10556 34580 10558
rect 34300 10546 34356 10556
rect 33740 9886 33742 9938
rect 33794 9886 33796 9938
rect 33740 9874 33796 9886
rect 34524 9266 34580 10556
rect 34524 9214 34526 9266
rect 34578 9214 34580 9266
rect 34524 9202 34580 9214
rect 34076 8930 34132 8942
rect 34076 8878 34078 8930
rect 34130 8878 34132 8930
rect 34076 8596 34132 8878
rect 34132 8540 34468 8596
rect 34076 8530 34132 8540
rect 34412 8370 34468 8540
rect 34412 8318 34414 8370
rect 34466 8318 34468 8370
rect 34412 8306 34468 8318
rect 33740 7364 33796 7374
rect 33628 7308 33740 7364
rect 33740 7298 33796 7308
rect 34412 7364 34468 7374
rect 34412 7270 34468 7308
rect 33292 6290 33348 6300
rect 34188 6916 34244 6926
rect 33292 6020 33348 6030
rect 32508 5966 32510 6018
rect 32562 5966 32564 6018
rect 32508 5954 32564 5966
rect 32732 6018 33348 6020
rect 32732 5966 33294 6018
rect 33346 5966 33348 6018
rect 32732 5964 33348 5966
rect 32732 5234 32788 5964
rect 33292 5954 33348 5964
rect 33628 5908 33684 5918
rect 33628 5814 33684 5852
rect 32732 5182 32734 5234
rect 32786 5182 32788 5234
rect 32732 5170 32788 5182
rect 33292 5012 33348 5022
rect 33292 4562 33348 4956
rect 33292 4510 33294 4562
rect 33346 4510 33348 4562
rect 33292 4498 33348 4510
rect 34188 4450 34244 6860
rect 34300 5908 34356 5918
rect 34300 5814 34356 5852
rect 34636 5908 34692 12460
rect 35084 12404 35140 21756
rect 35308 21746 35364 21756
rect 35980 22036 36036 22046
rect 35980 21586 36036 21980
rect 35980 21534 35982 21586
rect 36034 21534 36036 21586
rect 35980 21522 36036 21534
rect 36092 20802 36148 23326
rect 36428 23380 36484 23390
rect 36204 22370 36260 22382
rect 36204 22318 36206 22370
rect 36258 22318 36260 22370
rect 36204 21812 36260 22318
rect 36428 22258 36484 23324
rect 36428 22206 36430 22258
rect 36482 22206 36484 22258
rect 36428 22194 36484 22206
rect 36540 23154 36596 23436
rect 36652 23268 36708 23278
rect 36652 23174 36708 23212
rect 36540 23102 36542 23154
rect 36594 23102 36596 23154
rect 36540 22036 36596 23102
rect 36540 21970 36596 21980
rect 36764 22932 36820 24558
rect 37212 24052 37268 25004
rect 37212 23986 37268 23996
rect 37100 23714 37156 23726
rect 37100 23662 37102 23714
rect 37154 23662 37156 23714
rect 37100 23604 37156 23662
rect 37100 23538 37156 23548
rect 37212 23154 37268 23166
rect 37212 23102 37214 23154
rect 37266 23102 37268 23154
rect 37212 22932 37268 23102
rect 37324 23044 37380 26852
rect 37436 26178 37492 27468
rect 37548 27186 37604 28140
rect 37548 27134 37550 27186
rect 37602 27134 37604 27186
rect 37548 26908 37604 27134
rect 37660 27076 37716 28700
rect 38556 28690 38612 28700
rect 38220 28644 38276 28654
rect 38220 28420 38276 28588
rect 38668 28644 38724 28654
rect 38668 28530 38724 28588
rect 38668 28478 38670 28530
rect 38722 28478 38724 28530
rect 38668 28466 38724 28478
rect 38780 28420 38836 28430
rect 38220 28364 38500 28420
rect 38108 28196 38164 28206
rect 37996 27858 38052 27870
rect 37996 27806 37998 27858
rect 38050 27806 38052 27858
rect 37996 27748 38052 27806
rect 37996 27682 38052 27692
rect 38108 27524 38164 28140
rect 38444 27970 38500 28364
rect 38780 28082 38836 28364
rect 38892 28196 38948 29374
rect 39004 29650 39060 29662
rect 39004 29598 39006 29650
rect 39058 29598 39060 29650
rect 39004 29540 39060 29598
rect 39004 28756 39060 29484
rect 39116 29092 39172 29820
rect 39340 29428 39396 29438
rect 39116 29036 39284 29092
rect 39004 28530 39060 28700
rect 39004 28478 39006 28530
rect 39058 28478 39060 28530
rect 39004 28466 39060 28478
rect 39116 28644 39172 28654
rect 38892 28130 38948 28140
rect 38780 28030 38782 28082
rect 38834 28030 38836 28082
rect 38780 28018 38836 28030
rect 38444 27918 38446 27970
rect 38498 27918 38500 27970
rect 38444 27906 38500 27918
rect 38668 27972 38724 27982
rect 37996 27468 38164 27524
rect 38332 27858 38388 27870
rect 38332 27806 38334 27858
rect 38386 27806 38388 27858
rect 37660 27010 37716 27020
rect 37884 27076 37940 27114
rect 37884 27010 37940 27020
rect 37548 26852 37940 26908
rect 37884 26402 37940 26852
rect 37996 26628 38052 27468
rect 38332 27412 38388 27806
rect 38332 27346 38388 27356
rect 38556 27636 38612 27646
rect 38220 27188 38276 27198
rect 38556 27188 38612 27580
rect 38220 27186 38612 27188
rect 38220 27134 38222 27186
rect 38274 27134 38612 27186
rect 38220 27132 38612 27134
rect 38220 27122 38276 27132
rect 38556 27074 38612 27132
rect 38556 27022 38558 27074
rect 38610 27022 38612 27074
rect 38556 27010 38612 27022
rect 38108 26852 38164 26862
rect 38108 26850 38500 26852
rect 38108 26798 38110 26850
rect 38162 26798 38500 26850
rect 38108 26796 38500 26798
rect 38108 26786 38164 26796
rect 37996 26572 38276 26628
rect 37884 26350 37886 26402
rect 37938 26350 37940 26402
rect 37884 26338 37940 26350
rect 37996 26290 38052 26302
rect 37996 26238 37998 26290
rect 38050 26238 38052 26290
rect 37436 26126 37438 26178
rect 37490 26126 37492 26178
rect 37436 24500 37492 26126
rect 37548 26180 37604 26190
rect 37996 26180 38052 26238
rect 37548 26178 38052 26180
rect 37548 26126 37550 26178
rect 37602 26126 38052 26178
rect 37548 26124 38052 26126
rect 37548 26114 37604 26124
rect 37548 25956 37604 25966
rect 37548 25282 37604 25900
rect 37996 25844 38052 26124
rect 37996 25778 38052 25788
rect 38108 25956 38164 25966
rect 38108 25396 38164 25900
rect 38108 25330 38164 25340
rect 37548 25230 37550 25282
rect 37602 25230 37604 25282
rect 37548 24834 37604 25230
rect 38220 25284 38276 26572
rect 38444 26292 38500 26796
rect 38668 26628 38724 27916
rect 38780 27860 38836 27870
rect 39116 27860 39172 28588
rect 39228 28084 39284 29036
rect 39340 28642 39396 29372
rect 39340 28590 39342 28642
rect 39394 28590 39396 28642
rect 39340 28578 39396 28590
rect 39564 28644 39620 37548
rect 41020 36594 41076 39200
rect 41020 36542 41022 36594
rect 41074 36542 41076 36594
rect 41020 36530 41076 36542
rect 41580 37492 41636 37502
rect 40012 36260 40068 36270
rect 40012 36258 40292 36260
rect 40012 36206 40014 36258
rect 40066 36206 40292 36258
rect 40012 36204 40292 36206
rect 40012 36194 40068 36204
rect 39852 36092 40116 36102
rect 39908 36036 39956 36092
rect 40012 36036 40060 36092
rect 39852 36026 40116 36036
rect 39900 35586 39956 35598
rect 39900 35534 39902 35586
rect 39954 35534 39956 35586
rect 39900 34692 39956 35534
rect 40012 35474 40068 35486
rect 40012 35422 40014 35474
rect 40066 35422 40068 35474
rect 40012 34916 40068 35422
rect 40236 35252 40292 36204
rect 40236 34916 40292 35196
rect 40572 35588 40628 35598
rect 40460 35140 40516 35150
rect 40348 34916 40404 34926
rect 40236 34914 40404 34916
rect 40236 34862 40350 34914
rect 40402 34862 40404 34914
rect 40236 34860 40404 34862
rect 40460 34916 40516 35084
rect 40572 35140 40628 35532
rect 40572 35138 40852 35140
rect 40572 35086 40574 35138
rect 40626 35086 40852 35138
rect 40572 35084 40852 35086
rect 40572 35074 40628 35084
rect 40572 34916 40628 34926
rect 40460 34914 40628 34916
rect 40460 34862 40574 34914
rect 40626 34862 40628 34914
rect 40460 34860 40628 34862
rect 40012 34850 40068 34860
rect 40348 34804 40404 34860
rect 40348 34738 40404 34748
rect 39900 34636 40292 34692
rect 39852 34524 40116 34534
rect 39908 34468 39956 34524
rect 40012 34468 40060 34524
rect 39852 34458 40116 34468
rect 40124 34132 40180 34142
rect 40236 34132 40292 34636
rect 40124 34130 40292 34132
rect 40124 34078 40126 34130
rect 40178 34078 40292 34130
rect 40124 34076 40292 34078
rect 39676 34020 39732 34030
rect 39676 32788 39732 33964
rect 40124 33684 40180 34076
rect 40124 33628 40516 33684
rect 39852 32956 40116 32966
rect 39908 32900 39956 32956
rect 40012 32900 40060 32956
rect 39852 32890 40116 32900
rect 39676 32732 39844 32788
rect 39676 32564 39732 32574
rect 39676 32470 39732 32508
rect 39788 31892 39844 32732
rect 39900 32676 39956 32686
rect 39900 32562 39956 32620
rect 39900 32510 39902 32562
rect 39954 32510 39956 32562
rect 39900 32498 39956 32510
rect 40236 32676 40292 32686
rect 39788 31826 39844 31836
rect 39852 31388 40116 31398
rect 39908 31332 39956 31388
rect 40012 31332 40060 31388
rect 39852 31322 40116 31332
rect 40012 31220 40068 31230
rect 40012 31126 40068 31164
rect 40236 31218 40292 32620
rect 40236 31166 40238 31218
rect 40290 31166 40292 31218
rect 40236 31154 40292 31166
rect 39788 30996 39844 31006
rect 39788 30902 39844 30940
rect 40236 29988 40292 29998
rect 39852 29820 40116 29830
rect 39908 29764 39956 29820
rect 40012 29764 40060 29820
rect 39852 29754 40116 29764
rect 40012 29652 40068 29662
rect 40012 29558 40068 29596
rect 40236 29538 40292 29932
rect 40236 29486 40238 29538
rect 40290 29486 40292 29538
rect 39788 29428 39844 29438
rect 39564 28578 39620 28588
rect 39676 29372 39788 29428
rect 39228 28018 39284 28028
rect 39564 28418 39620 28430
rect 39564 28366 39566 28418
rect 39618 28366 39620 28418
rect 39564 27972 39620 28366
rect 39676 27972 39732 29372
rect 39788 29362 39844 29372
rect 40124 29426 40180 29438
rect 40124 29374 40126 29426
rect 40178 29374 40180 29426
rect 40124 28868 40180 29374
rect 40124 28802 40180 28812
rect 39788 28756 39844 28766
rect 39788 28642 39844 28700
rect 39788 28590 39790 28642
rect 39842 28590 39844 28642
rect 39788 28578 39844 28590
rect 40236 28532 40292 29486
rect 40348 29428 40404 29438
rect 40348 28866 40404 29372
rect 40348 28814 40350 28866
rect 40402 28814 40404 28866
rect 40348 28802 40404 28814
rect 40460 28644 40516 33628
rect 40460 28578 40516 28588
rect 40236 28476 40404 28532
rect 39900 28420 39956 28458
rect 39900 28354 39956 28364
rect 40124 28420 40180 28430
rect 40124 28418 40292 28420
rect 40124 28366 40126 28418
rect 40178 28366 40292 28418
rect 40124 28364 40292 28366
rect 40124 28354 40180 28364
rect 39852 28252 40116 28262
rect 39908 28196 39956 28252
rect 40012 28196 40060 28252
rect 39852 28186 40116 28196
rect 39900 28084 39956 28094
rect 39788 27972 39844 27982
rect 39676 27970 39844 27972
rect 39676 27918 39790 27970
rect 39842 27918 39844 27970
rect 39676 27916 39844 27918
rect 39564 27906 39620 27916
rect 39788 27906 39844 27916
rect 38780 27074 38836 27804
rect 38780 27022 38782 27074
rect 38834 27022 38836 27074
rect 38780 27010 38836 27022
rect 38892 27804 39172 27860
rect 38444 26290 38612 26292
rect 38444 26238 38446 26290
rect 38498 26238 38612 26290
rect 38444 26236 38612 26238
rect 38444 26226 38500 26236
rect 38444 25844 38500 25854
rect 38444 25506 38500 25788
rect 38444 25454 38446 25506
rect 38498 25454 38500 25506
rect 38444 25442 38500 25454
rect 38556 25396 38612 26236
rect 38668 26290 38724 26572
rect 38780 26740 38836 26750
rect 38780 26514 38836 26684
rect 38780 26462 38782 26514
rect 38834 26462 38836 26514
rect 38780 26450 38836 26462
rect 38892 26404 38948 27804
rect 39340 27748 39396 27758
rect 39340 27654 39396 27692
rect 39116 27634 39172 27646
rect 39116 27582 39118 27634
rect 39170 27582 39172 27634
rect 39004 27524 39060 27534
rect 39004 27298 39060 27468
rect 39116 27412 39172 27582
rect 39676 27634 39732 27646
rect 39676 27582 39678 27634
rect 39730 27582 39732 27634
rect 39116 27346 39172 27356
rect 39340 27524 39396 27534
rect 39004 27246 39006 27298
rect 39058 27246 39060 27298
rect 39004 27234 39060 27246
rect 39340 27076 39396 27468
rect 39676 27524 39732 27582
rect 39676 27458 39732 27468
rect 39900 27300 39956 28028
rect 40236 27970 40292 28364
rect 40236 27918 40238 27970
rect 40290 27918 40292 27970
rect 40236 27906 40292 27918
rect 40124 27636 40180 27646
rect 40124 27542 40180 27580
rect 39340 27010 39396 27020
rect 39452 27244 39956 27300
rect 39340 26852 39396 26862
rect 39340 26758 39396 26796
rect 38892 26348 39060 26404
rect 38668 26238 38670 26290
rect 38722 26238 38724 26290
rect 38668 26226 38724 26238
rect 38556 25330 38612 25340
rect 38668 25956 38724 25966
rect 38276 25228 38500 25284
rect 38220 25190 38276 25228
rect 38444 25060 38500 25228
rect 38444 25004 38612 25060
rect 37548 24782 37550 24834
rect 37602 24782 37604 24834
rect 37548 24770 37604 24782
rect 38444 24836 38500 24846
rect 37436 24434 37492 24444
rect 37660 24722 37716 24734
rect 37660 24670 37662 24722
rect 37714 24670 37716 24722
rect 37660 24164 37716 24670
rect 37884 24722 37940 24734
rect 37884 24670 37886 24722
rect 37938 24670 37940 24722
rect 37884 24500 37940 24670
rect 37884 24434 37940 24444
rect 38220 24724 38276 24734
rect 37660 24108 38164 24164
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 38108 23938 38164 24108
rect 38108 23886 38110 23938
rect 38162 23886 38164 23938
rect 38108 23828 38164 23886
rect 38220 23938 38276 24668
rect 38220 23886 38222 23938
rect 38274 23886 38276 23938
rect 38220 23874 38276 23886
rect 38332 24610 38388 24622
rect 38332 24558 38334 24610
rect 38386 24558 38388 24610
rect 38108 23762 38164 23772
rect 38108 23604 38164 23614
rect 37324 22988 37940 23044
rect 37212 22876 37604 22932
rect 36204 21252 36260 21756
rect 36428 21588 36484 21598
rect 36204 21186 36260 21196
rect 36316 21476 36372 21486
rect 36092 20750 36094 20802
rect 36146 20750 36148 20802
rect 36092 20738 36148 20750
rect 35420 20692 35476 20702
rect 35420 20018 35476 20636
rect 36316 20580 36372 21420
rect 36428 20916 36484 21532
rect 36428 20692 36484 20860
rect 36428 20626 36484 20636
rect 36316 20130 36372 20524
rect 36316 20078 36318 20130
rect 36370 20078 36372 20130
rect 36316 20066 36372 20078
rect 35420 19966 35422 20018
rect 35474 19966 35476 20018
rect 35420 19954 35476 19966
rect 35532 19906 35588 19918
rect 35532 19854 35534 19906
rect 35586 19854 35588 19906
rect 35420 19796 35476 19806
rect 35308 19684 35364 19694
rect 35196 17666 35252 17678
rect 35196 17614 35198 17666
rect 35250 17614 35252 17666
rect 35196 17444 35252 17614
rect 35196 17378 35252 17388
rect 35308 16436 35364 19628
rect 35420 19234 35476 19740
rect 35420 19182 35422 19234
rect 35474 19182 35476 19234
rect 35420 19170 35476 19182
rect 35532 18562 35588 19854
rect 36764 19908 36820 22876
rect 37212 22482 37268 22494
rect 37212 22430 37214 22482
rect 37266 22430 37268 22482
rect 37100 22370 37156 22382
rect 37100 22318 37102 22370
rect 37154 22318 37156 22370
rect 36988 22260 37044 22270
rect 36988 22166 37044 22204
rect 36988 21698 37044 21710
rect 36988 21646 36990 21698
rect 37042 21646 37044 21698
rect 36764 19842 36820 19852
rect 36876 21474 36932 21486
rect 36876 21422 36878 21474
rect 36930 21422 36932 21474
rect 36428 19236 36484 19246
rect 36428 19142 36484 19180
rect 35532 18510 35534 18562
rect 35586 18510 35588 18562
rect 35420 17554 35476 17566
rect 35420 17502 35422 17554
rect 35474 17502 35476 17554
rect 35420 17108 35476 17502
rect 35532 17556 35588 18510
rect 35532 17490 35588 17500
rect 35644 19122 35700 19134
rect 35644 19070 35646 19122
rect 35698 19070 35700 19122
rect 35644 17780 35700 19070
rect 36876 18788 36932 21422
rect 36988 21476 37044 21646
rect 37100 21588 37156 22318
rect 37100 21522 37156 21532
rect 36988 21410 37044 21420
rect 36652 18732 36876 18788
rect 36428 18676 36484 18686
rect 36316 18674 36484 18676
rect 36316 18622 36430 18674
rect 36482 18622 36484 18674
rect 36316 18620 36484 18622
rect 35420 17042 35476 17052
rect 35644 16882 35700 17724
rect 35644 16830 35646 16882
rect 35698 16830 35700 16882
rect 35532 16772 35588 16782
rect 35532 16678 35588 16716
rect 35196 15876 35252 15886
rect 35196 15538 35252 15820
rect 35196 15486 35198 15538
rect 35250 15486 35252 15538
rect 35196 15474 35252 15486
rect 35196 13748 35252 13758
rect 35196 12962 35252 13692
rect 35308 13188 35364 16380
rect 35420 16658 35476 16670
rect 35420 16606 35422 16658
rect 35474 16606 35476 16658
rect 35420 16212 35476 16606
rect 35420 16146 35476 16156
rect 35644 16100 35700 16830
rect 35644 16034 35700 16044
rect 35868 18004 35924 18014
rect 35868 16098 35924 17948
rect 36092 17892 36148 17902
rect 36092 17554 36148 17836
rect 36092 17502 36094 17554
rect 36146 17502 36148 17554
rect 36092 17490 36148 17502
rect 36204 17666 36260 17678
rect 36204 17614 36206 17666
rect 36258 17614 36260 17666
rect 36204 17556 36260 17614
rect 36204 17490 36260 17500
rect 36316 16324 36372 18620
rect 36428 18610 36484 18620
rect 36540 18450 36596 18462
rect 36540 18398 36542 18450
rect 36594 18398 36596 18450
rect 36540 17892 36596 18398
rect 36540 17826 36596 17836
rect 36316 16258 36372 16268
rect 36428 17220 36484 17230
rect 35868 16046 35870 16098
rect 35922 16046 35924 16098
rect 35756 15316 35812 15326
rect 35868 15316 35924 16046
rect 36428 15988 36484 17164
rect 36092 15986 36484 15988
rect 36092 15934 36430 15986
rect 36482 15934 36484 15986
rect 36092 15932 36484 15934
rect 35980 15876 36036 15886
rect 35980 15782 36036 15820
rect 36092 15428 36148 15932
rect 36428 15922 36484 15932
rect 36652 15988 36708 18732
rect 36876 18722 36932 18732
rect 37212 18676 37268 22430
rect 37100 18620 37268 18676
rect 37324 20802 37380 20814
rect 37324 20750 37326 20802
rect 37378 20750 37380 20802
rect 37324 19012 37380 20750
rect 37548 20356 37604 22876
rect 37548 20018 37604 20300
rect 37548 19966 37550 20018
rect 37602 19966 37604 20018
rect 37548 19954 37604 19966
rect 37772 20018 37828 20030
rect 37772 19966 37774 20018
rect 37826 19966 37828 20018
rect 37772 19012 37828 19966
rect 37324 19010 37828 19012
rect 37324 18958 37326 19010
rect 37378 18958 37828 19010
rect 37324 18956 37828 18958
rect 37100 18228 37156 18620
rect 37324 18564 37380 18956
rect 37324 18498 37380 18508
rect 37436 18788 37492 18798
rect 37436 18562 37492 18732
rect 37436 18510 37438 18562
rect 37490 18510 37492 18562
rect 37436 18498 37492 18510
rect 37660 18788 37716 18798
rect 37100 18172 37268 18228
rect 36988 18004 37044 18014
rect 36988 17666 37044 17948
rect 36988 17614 36990 17666
rect 37042 17614 37044 17666
rect 36988 17602 37044 17614
rect 37212 17668 37268 18172
rect 37548 17780 37604 17790
rect 37660 17780 37716 18732
rect 37548 17778 37716 17780
rect 37548 17726 37550 17778
rect 37602 17726 37716 17778
rect 37548 17724 37716 17726
rect 37548 17714 37604 17724
rect 35756 15314 35924 15316
rect 35756 15262 35758 15314
rect 35810 15262 35924 15314
rect 35756 15260 35924 15262
rect 35980 15372 36148 15428
rect 35756 15250 35812 15260
rect 35532 15202 35588 15214
rect 35532 15150 35534 15202
rect 35586 15150 35588 15202
rect 35532 15148 35588 15150
rect 35980 15148 36036 15372
rect 36652 15314 36708 15932
rect 36764 16884 36820 16894
rect 36764 15426 36820 16828
rect 37212 16882 37268 17612
rect 37212 16830 37214 16882
rect 37266 16830 37268 16882
rect 37212 16818 37268 16830
rect 37548 17332 37604 17342
rect 36988 16772 37044 16782
rect 37436 16772 37492 16782
rect 36988 16098 37044 16716
rect 36988 16046 36990 16098
rect 37042 16046 37044 16098
rect 36988 16034 37044 16046
rect 37324 16716 37436 16772
rect 37324 15988 37380 16716
rect 37436 16706 37492 16716
rect 36764 15374 36766 15426
rect 36818 15374 36820 15426
rect 36764 15362 36820 15374
rect 37212 15932 37380 15988
rect 36652 15262 36654 15314
rect 36706 15262 36708 15314
rect 36652 15250 36708 15262
rect 35532 15092 36036 15148
rect 36764 15204 36820 15242
rect 36764 15138 36820 15148
rect 36092 15090 36148 15102
rect 36092 15038 36094 15090
rect 36146 15038 36148 15090
rect 35644 14532 35700 14542
rect 36092 14532 36148 15038
rect 36204 14532 36260 14542
rect 36092 14476 36204 14532
rect 35644 14438 35700 14476
rect 36204 14438 36260 14476
rect 37100 14084 37156 14094
rect 35308 13122 35364 13132
rect 35420 13860 35476 13870
rect 35196 12910 35198 12962
rect 35250 12910 35252 12962
rect 35196 12898 35252 12910
rect 35308 12964 35364 12974
rect 35308 12870 35364 12908
rect 35420 12964 35476 13804
rect 35644 13860 35700 13870
rect 35644 13766 35700 13804
rect 36092 13636 36148 13646
rect 35980 13634 36148 13636
rect 35980 13582 36094 13634
rect 36146 13582 36148 13634
rect 35980 13580 36148 13582
rect 35420 12962 35924 12964
rect 35420 12910 35422 12962
rect 35474 12910 35924 12962
rect 35420 12908 35924 12910
rect 35420 12898 35476 12908
rect 35532 12740 35588 12750
rect 35644 12740 35700 12750
rect 35532 12738 35644 12740
rect 35532 12686 35534 12738
rect 35586 12686 35644 12738
rect 35532 12684 35644 12686
rect 35532 12674 35588 12684
rect 34972 12348 35140 12404
rect 34860 9828 34916 9838
rect 34860 9042 34916 9772
rect 34972 9268 35028 12348
rect 34972 9202 35028 9212
rect 35084 12180 35140 12190
rect 34860 8990 34862 9042
rect 34914 8990 34916 9042
rect 34860 8978 34916 8990
rect 35084 8820 35140 12124
rect 35420 12068 35476 12078
rect 35420 12066 35588 12068
rect 35420 12014 35422 12066
rect 35474 12014 35588 12066
rect 35420 12012 35588 12014
rect 35420 12002 35476 12012
rect 34860 8764 35140 8820
rect 35420 9154 35476 9166
rect 35420 9102 35422 9154
rect 35474 9102 35476 9154
rect 34748 8034 34804 8046
rect 34748 7982 34750 8034
rect 34802 7982 34804 8034
rect 34748 6916 34804 7982
rect 34860 7252 34916 8764
rect 34972 8596 35028 8606
rect 35420 8596 35476 9102
rect 35028 8540 35476 8596
rect 34972 8258 35028 8540
rect 34972 8206 34974 8258
rect 35026 8206 35028 8258
rect 34972 8194 35028 8206
rect 34860 7186 34916 7196
rect 34748 6850 34804 6860
rect 35196 6916 35252 6926
rect 35084 6468 35140 6478
rect 34636 5906 34916 5908
rect 34636 5854 34638 5906
rect 34690 5854 34916 5906
rect 34636 5852 34916 5854
rect 34636 5842 34692 5852
rect 34860 5234 34916 5852
rect 34860 5182 34862 5234
rect 34914 5182 34916 5234
rect 34860 5170 34916 5182
rect 35084 4564 35140 6412
rect 35196 6018 35252 6860
rect 35420 6468 35476 6478
rect 35196 5966 35198 6018
rect 35250 5966 35252 6018
rect 35196 5954 35252 5966
rect 35308 6466 35476 6468
rect 35308 6414 35422 6466
rect 35474 6414 35476 6466
rect 35308 6412 35476 6414
rect 34188 4398 34190 4450
rect 34242 4398 34244 4450
rect 34188 4386 34244 4398
rect 34412 4562 35140 4564
rect 34412 4510 35086 4562
rect 35138 4510 35140 4562
rect 34412 4508 35140 4510
rect 32508 4340 32564 4350
rect 32508 4228 32564 4284
rect 33628 4340 33684 4350
rect 33628 4246 33684 4284
rect 34412 4338 34468 4508
rect 35084 4498 35140 4508
rect 35308 5906 35364 6412
rect 35420 6402 35476 6412
rect 35308 5854 35310 5906
rect 35362 5854 35364 5906
rect 34412 4286 34414 4338
rect 34466 4286 34468 4338
rect 34412 4274 34468 4286
rect 32396 4226 32564 4228
rect 32396 4174 32510 4226
rect 32562 4174 32564 4226
rect 32396 4172 32564 4174
rect 32508 4162 32564 4172
rect 35308 4228 35364 5854
rect 35420 5124 35476 5134
rect 35420 5030 35476 5068
rect 35532 4900 35588 12012
rect 35644 11396 35700 12684
rect 35644 11340 35812 11396
rect 35644 9044 35700 9054
rect 35644 8950 35700 8988
rect 35644 8258 35700 8270
rect 35644 8206 35646 8258
rect 35698 8206 35700 8258
rect 35644 8148 35700 8206
rect 35644 8082 35700 8092
rect 35756 7812 35812 11340
rect 35868 9938 35924 12908
rect 35980 12740 36036 13580
rect 36092 13570 36148 13580
rect 36652 13634 36708 13646
rect 36652 13582 36654 13634
rect 36706 13582 36708 13634
rect 36316 13188 36372 13198
rect 36652 13188 36708 13582
rect 37100 13634 37156 14028
rect 37100 13582 37102 13634
rect 37154 13582 37156 13634
rect 37100 13524 37156 13582
rect 37100 13458 37156 13468
rect 37212 13300 37268 15932
rect 37548 15876 37604 17276
rect 36372 13132 36708 13188
rect 37100 13244 37268 13300
rect 37324 15820 37604 15876
rect 35980 12674 36036 12684
rect 36092 12740 36148 12750
rect 36316 12740 36372 13132
rect 37100 12852 37156 13244
rect 37212 13076 37268 13086
rect 37212 12982 37268 13020
rect 37100 12796 37268 12852
rect 36092 12738 36372 12740
rect 36092 12686 36094 12738
rect 36146 12686 36372 12738
rect 36092 12684 36372 12686
rect 36428 12738 36484 12750
rect 36428 12686 36430 12738
rect 36482 12686 36484 12738
rect 36092 12404 36148 12684
rect 36428 12516 36484 12686
rect 36428 12450 36484 12460
rect 36092 12338 36148 12348
rect 36204 12178 36260 12190
rect 36204 12126 36206 12178
rect 36258 12126 36260 12178
rect 36204 11844 36260 12126
rect 36988 12068 37044 12078
rect 36988 12066 37156 12068
rect 36988 12014 36990 12066
rect 37042 12014 37156 12066
rect 36988 12012 37156 12014
rect 36988 12002 37044 12012
rect 35980 11788 36204 11844
rect 35980 11506 36036 11788
rect 36204 11778 36260 11788
rect 35980 11454 35982 11506
rect 36034 11454 36036 11506
rect 35980 11442 36036 11454
rect 36428 11172 36484 11182
rect 36428 11078 36484 11116
rect 36988 11170 37044 11182
rect 36988 11118 36990 11170
rect 37042 11118 37044 11170
rect 36988 11060 37044 11118
rect 36988 10994 37044 11004
rect 35868 9886 35870 9938
rect 35922 9886 35924 9938
rect 35868 9828 35924 9886
rect 35868 9762 35924 9772
rect 36204 9044 36260 9054
rect 36204 8950 36260 8988
rect 36988 8372 37044 8382
rect 37100 8372 37156 12012
rect 37212 11396 37268 12796
rect 37324 11732 37380 15820
rect 37436 15652 37492 15662
rect 37436 15314 37492 15596
rect 37436 15262 37438 15314
rect 37490 15262 37492 15314
rect 37436 14530 37492 15262
rect 37660 14642 37716 17724
rect 37660 14590 37662 14642
rect 37714 14590 37716 14642
rect 37660 14578 37716 14590
rect 37772 15204 37828 15214
rect 37436 14478 37438 14530
rect 37490 14478 37492 14530
rect 37436 14466 37492 14478
rect 37548 13972 37604 13982
rect 37548 12964 37604 13916
rect 37772 13860 37828 15148
rect 37884 14084 37940 22988
rect 38108 19236 38164 23548
rect 38220 23042 38276 23054
rect 38220 22990 38222 23042
rect 38274 22990 38276 23042
rect 38220 20690 38276 22990
rect 38332 21924 38388 24558
rect 38444 23938 38500 24780
rect 38556 24164 38612 25004
rect 38668 24948 38724 25900
rect 39004 25956 39060 26348
rect 39004 25890 39060 25900
rect 38780 25844 38836 25854
rect 38780 25508 38836 25788
rect 39004 25620 39060 25630
rect 39004 25618 39396 25620
rect 39004 25566 39006 25618
rect 39058 25566 39396 25618
rect 39004 25564 39396 25566
rect 39004 25554 39060 25564
rect 38780 25442 38836 25452
rect 38892 25396 38948 25406
rect 38892 25302 38948 25340
rect 39116 25396 39172 25434
rect 39116 25330 39172 25340
rect 38780 24948 38836 24958
rect 38668 24946 38948 24948
rect 38668 24894 38782 24946
rect 38834 24894 38948 24946
rect 38668 24892 38948 24894
rect 38780 24882 38836 24892
rect 38556 24098 38612 24108
rect 38444 23886 38446 23938
rect 38498 23886 38500 23938
rect 38444 23874 38500 23886
rect 38780 23940 38836 23950
rect 38780 23846 38836 23884
rect 38780 23268 38836 23278
rect 38780 22596 38836 23212
rect 38892 23044 38948 24892
rect 39228 24722 39284 24734
rect 39228 24670 39230 24722
rect 39282 24670 39284 24722
rect 39116 23940 39172 23950
rect 38892 22978 38948 22988
rect 39004 23042 39060 23054
rect 39004 22990 39006 23042
rect 39058 22990 39060 23042
rect 39004 22932 39060 22990
rect 39004 22866 39060 22876
rect 38780 22540 39060 22596
rect 38332 21868 38612 21924
rect 38444 21700 38500 21710
rect 38444 21606 38500 21644
rect 38556 21588 38612 21868
rect 38780 21812 38836 21822
rect 38780 21718 38836 21756
rect 38668 21588 38724 21598
rect 38556 21586 38836 21588
rect 38556 21534 38670 21586
rect 38722 21534 38836 21586
rect 38556 21532 38836 21534
rect 38668 21494 38724 21532
rect 38220 20638 38222 20690
rect 38274 20638 38276 20690
rect 38220 19460 38276 20638
rect 38668 20580 38724 20590
rect 38220 19394 38276 19404
rect 38556 20578 38724 20580
rect 38556 20526 38670 20578
rect 38722 20526 38724 20578
rect 38556 20524 38724 20526
rect 38108 19180 38500 19236
rect 38108 19012 38164 19022
rect 38108 18918 38164 18956
rect 37996 18452 38052 18462
rect 37996 18358 38052 18396
rect 38220 16100 38276 16110
rect 38220 16006 38276 16044
rect 38332 15652 38388 15662
rect 38220 15202 38276 15214
rect 38220 15150 38222 15202
rect 38274 15150 38276 15202
rect 38108 14756 38164 14766
rect 37996 14644 38052 14654
rect 37996 14550 38052 14588
rect 37884 14028 38052 14084
rect 37884 13860 37940 13870
rect 37772 13858 37940 13860
rect 37772 13806 37886 13858
rect 37938 13806 37940 13858
rect 37772 13804 37940 13806
rect 37884 13794 37940 13804
rect 37772 13188 37828 13198
rect 37660 12964 37716 12974
rect 37548 12962 37716 12964
rect 37548 12910 37662 12962
rect 37714 12910 37716 12962
rect 37548 12908 37716 12910
rect 37660 12898 37716 12908
rect 37436 12740 37492 12750
rect 37436 12738 37716 12740
rect 37436 12686 37438 12738
rect 37490 12686 37716 12738
rect 37436 12684 37716 12686
rect 37436 12674 37492 12684
rect 37324 11666 37380 11676
rect 37212 11340 37604 11396
rect 37324 11172 37380 11182
rect 37044 8316 37156 8372
rect 37212 9938 37268 9950
rect 37212 9886 37214 9938
rect 37266 9886 37268 9938
rect 37212 9044 37268 9886
rect 37324 9828 37380 11116
rect 37324 9762 37380 9772
rect 37548 9826 37604 11340
rect 37660 10612 37716 12684
rect 37772 12180 37828 13132
rect 37772 12114 37828 12124
rect 37996 11620 38052 14028
rect 38108 13746 38164 14700
rect 38108 13694 38110 13746
rect 38162 13694 38164 13746
rect 38108 13682 38164 13694
rect 38220 13188 38276 15150
rect 38332 14530 38388 15596
rect 38332 14478 38334 14530
rect 38386 14478 38388 14530
rect 38332 14466 38388 14478
rect 38444 13860 38500 19180
rect 38556 17444 38612 20524
rect 38668 20514 38724 20524
rect 38780 20468 38836 21532
rect 38892 21586 38948 21598
rect 38892 21534 38894 21586
rect 38946 21534 38948 21586
rect 38892 21476 38948 21534
rect 38892 21410 38948 21420
rect 39004 20914 39060 22540
rect 39004 20862 39006 20914
rect 39058 20862 39060 20914
rect 39004 20850 39060 20862
rect 39116 20692 39172 23884
rect 39228 23828 39284 24670
rect 39340 24724 39396 25564
rect 39340 24658 39396 24668
rect 39452 23938 39508 27244
rect 40236 27074 40292 27086
rect 40236 27022 40238 27074
rect 40290 27022 40292 27074
rect 39676 26962 39732 26974
rect 39676 26910 39678 26962
rect 39730 26910 39732 26962
rect 39676 26740 39732 26910
rect 39900 26964 39956 27002
rect 39900 26898 39956 26908
rect 39788 26852 39844 26890
rect 39788 26786 39844 26796
rect 39676 26674 39732 26684
rect 39852 26684 40116 26694
rect 39564 26628 39620 26638
rect 39908 26628 39956 26684
rect 40012 26628 40060 26684
rect 39852 26618 40116 26628
rect 39564 26516 39620 26572
rect 40124 26516 40180 26526
rect 39564 26460 39844 26516
rect 39676 26292 39732 26302
rect 39676 26178 39732 26236
rect 39676 26126 39678 26178
rect 39730 26126 39732 26178
rect 39676 26114 39732 26126
rect 39452 23886 39454 23938
rect 39506 23886 39508 23938
rect 39452 23874 39508 23886
rect 39564 25844 39620 25854
rect 39228 21698 39284 23772
rect 39340 23492 39396 23502
rect 39340 23268 39396 23436
rect 39340 23202 39396 23212
rect 39228 21646 39230 21698
rect 39282 21646 39284 21698
rect 39228 21634 39284 21646
rect 39340 22370 39396 22382
rect 39340 22318 39342 22370
rect 39394 22318 39396 22370
rect 38780 20402 38836 20412
rect 39004 20636 39172 20692
rect 39228 21476 39284 21486
rect 38780 19794 38836 19806
rect 38780 19742 38782 19794
rect 38834 19742 38836 19794
rect 38556 16882 38612 17388
rect 38668 17556 38724 17566
rect 38780 17556 38836 19742
rect 38668 17554 38836 17556
rect 38668 17502 38670 17554
rect 38722 17502 38836 17554
rect 38668 17500 38836 17502
rect 38892 19346 38948 19358
rect 38892 19294 38894 19346
rect 38946 19294 38948 19346
rect 38892 18452 38948 19294
rect 38668 17220 38724 17500
rect 38668 17154 38724 17164
rect 38556 16830 38558 16882
rect 38610 16830 38612 16882
rect 38556 16818 38612 16830
rect 38892 16884 38948 18396
rect 38668 16548 38724 16558
rect 38556 14756 38612 14766
rect 38556 14662 38612 14700
rect 38668 14196 38724 16492
rect 38892 16098 38948 16828
rect 38892 16046 38894 16098
rect 38946 16046 38948 16098
rect 38892 16034 38948 16046
rect 39004 15148 39060 20636
rect 39116 19234 39172 19246
rect 39116 19182 39118 19234
rect 39170 19182 39172 19234
rect 39116 19124 39172 19182
rect 39116 17108 39172 19068
rect 39228 18450 39284 21420
rect 39340 21028 39396 22318
rect 39340 20962 39396 20972
rect 39452 22260 39508 22270
rect 39452 19236 39508 22204
rect 39452 19170 39508 19180
rect 39228 18398 39230 18450
rect 39282 18398 39284 18450
rect 39228 18386 39284 18398
rect 39340 17556 39396 17566
rect 39340 17462 39396 17500
rect 39340 17108 39396 17118
rect 39116 17106 39396 17108
rect 39116 17054 39342 17106
rect 39394 17054 39396 17106
rect 39116 17052 39396 17054
rect 39340 17042 39396 17052
rect 39228 16658 39284 16670
rect 39228 16606 39230 16658
rect 39282 16606 39284 16658
rect 39116 16100 39172 16110
rect 39116 16006 39172 16044
rect 39228 15538 39284 16606
rect 39228 15486 39230 15538
rect 39282 15486 39284 15538
rect 39228 15474 39284 15486
rect 39564 15148 39620 25788
rect 39788 25508 39844 26460
rect 40124 26290 40180 26460
rect 40124 26238 40126 26290
rect 40178 26238 40180 26290
rect 40124 26226 40180 26238
rect 40012 26068 40068 26078
rect 40236 26068 40292 27022
rect 40012 25508 40068 26012
rect 40124 26012 40292 26068
rect 40348 26068 40404 28476
rect 40572 28308 40628 34860
rect 40796 34130 40852 35084
rect 41244 34916 41300 34926
rect 40796 34078 40798 34130
rect 40850 34078 40852 34130
rect 40796 33346 40852 34078
rect 41132 34804 41188 34814
rect 41132 34690 41188 34748
rect 41132 34638 41134 34690
rect 41186 34638 41188 34690
rect 41132 33908 41188 34638
rect 41244 34356 41300 34860
rect 41244 34262 41300 34300
rect 41468 34130 41524 34142
rect 41468 34078 41470 34130
rect 41522 34078 41524 34130
rect 41132 33842 41188 33852
rect 41356 34018 41412 34030
rect 41356 33966 41358 34018
rect 41410 33966 41412 34018
rect 40796 33294 40798 33346
rect 40850 33294 40852 33346
rect 40796 33282 40852 33294
rect 41356 32564 41412 33966
rect 41468 34020 41524 34078
rect 41468 33954 41524 33964
rect 41356 32498 41412 32508
rect 41244 31778 41300 31790
rect 41244 31726 41246 31778
rect 41298 31726 41300 31778
rect 41020 31668 41076 31678
rect 40796 31666 41076 31668
rect 40796 31614 41022 31666
rect 41074 31614 41076 31666
rect 40796 31612 41076 31614
rect 40796 31332 40852 31612
rect 41020 31602 41076 31612
rect 40684 28868 40740 28878
rect 40684 28774 40740 28812
rect 40124 25844 40180 26012
rect 40348 26002 40404 26012
rect 40460 28252 40628 28308
rect 40124 25788 40292 25844
rect 40236 25618 40292 25788
rect 40236 25566 40238 25618
rect 40290 25566 40292 25618
rect 40236 25554 40292 25566
rect 40124 25508 40180 25518
rect 40012 25506 40180 25508
rect 40012 25454 40126 25506
rect 40178 25454 40180 25506
rect 40012 25452 40180 25454
rect 39788 25442 39844 25452
rect 40124 25442 40180 25452
rect 40348 25506 40404 25518
rect 40348 25454 40350 25506
rect 40402 25454 40404 25506
rect 39676 25394 39732 25406
rect 39676 25342 39678 25394
rect 39730 25342 39732 25394
rect 39676 24948 39732 25342
rect 40348 25396 40404 25454
rect 40348 25330 40404 25340
rect 39900 25284 39956 25294
rect 39900 25282 40292 25284
rect 39900 25230 39902 25282
rect 39954 25230 40292 25282
rect 39900 25228 40292 25230
rect 39900 25218 39956 25228
rect 39852 25116 40116 25126
rect 39908 25060 39956 25116
rect 40012 25060 40060 25116
rect 39852 25050 40116 25060
rect 39676 24892 39956 24948
rect 39676 24724 39732 24734
rect 39676 24630 39732 24668
rect 39788 24610 39844 24622
rect 39788 24558 39790 24610
rect 39842 24558 39844 24610
rect 39788 24050 39844 24558
rect 39900 24164 39956 24892
rect 40012 24836 40068 24846
rect 40236 24836 40292 25228
rect 40068 24780 40292 24836
rect 40012 24742 40068 24780
rect 40460 24388 40516 28252
rect 40796 28084 40852 31276
rect 41244 31220 41300 31726
rect 41244 31154 41300 31164
rect 41020 30996 41076 31006
rect 41020 30902 41076 30940
rect 41468 30210 41524 30222
rect 41468 30158 41470 30210
rect 41522 30158 41524 30210
rect 41468 29652 41524 30158
rect 41580 30212 41636 37436
rect 42476 37380 42532 37390
rect 42140 35586 42196 35598
rect 42140 35534 42142 35586
rect 42194 35534 42196 35586
rect 42140 35364 42196 35534
rect 42140 35298 42196 35308
rect 41916 34356 41972 34366
rect 41916 34262 41972 34300
rect 41692 34130 41748 34142
rect 41692 34078 41694 34130
rect 41746 34078 41748 34130
rect 41692 32676 41748 34078
rect 42028 34130 42084 34142
rect 42028 34078 42030 34130
rect 42082 34078 42084 34130
rect 42028 34020 42084 34078
rect 42028 33954 42084 33964
rect 41692 32610 41748 32620
rect 42028 32450 42084 32462
rect 42028 32398 42030 32450
rect 42082 32398 42084 32450
rect 42028 31668 42084 32398
rect 42364 32452 42420 32462
rect 42364 31892 42420 32396
rect 42252 31668 42308 31678
rect 42028 31666 42308 31668
rect 42028 31614 42254 31666
rect 42306 31614 42308 31666
rect 42028 31612 42308 31614
rect 42140 30994 42196 31006
rect 42140 30942 42142 30994
rect 42194 30942 42196 30994
rect 41804 30884 41860 30894
rect 42140 30884 42196 30942
rect 41804 30882 42196 30884
rect 41804 30830 41806 30882
rect 41858 30830 42196 30882
rect 41804 30828 42196 30830
rect 42252 30884 42308 31612
rect 42364 31666 42420 31836
rect 42364 31614 42366 31666
rect 42418 31614 42420 31666
rect 42364 31602 42420 31614
rect 42476 30996 42532 37324
rect 43484 36708 43540 39200
rect 45948 39060 46004 39200
rect 46172 39060 46228 39228
rect 45948 39004 46228 39060
rect 44380 37268 44436 37278
rect 44436 37212 44548 37268
rect 44380 37202 44436 37212
rect 43932 36708 43988 36718
rect 43484 36706 43988 36708
rect 43484 36654 43934 36706
rect 43986 36654 43988 36706
rect 43484 36652 43988 36654
rect 43932 36642 43988 36652
rect 43036 36484 43092 36494
rect 43036 36390 43092 36428
rect 43260 35588 43316 35598
rect 43036 35028 43092 35038
rect 43036 34934 43092 34972
rect 42588 34804 42644 34814
rect 42588 33796 42644 34748
rect 42588 33730 42644 33740
rect 43036 33460 43092 33470
rect 43036 33234 43092 33404
rect 43036 33182 43038 33234
rect 43090 33182 43092 33234
rect 43036 33170 43092 33182
rect 42700 33122 42756 33134
rect 42700 33070 42702 33122
rect 42754 33070 42756 33122
rect 42700 32788 42756 33070
rect 42700 32722 42756 32732
rect 43036 32788 43092 32798
rect 43036 32694 43092 32732
rect 42700 32452 42756 32462
rect 42700 32358 42756 32396
rect 42588 31836 43204 31892
rect 42588 31778 42644 31836
rect 42588 31726 42590 31778
rect 42642 31726 42644 31778
rect 42588 31714 42644 31726
rect 43148 31778 43204 31836
rect 43148 31726 43150 31778
rect 43202 31726 43204 31778
rect 43148 31714 43204 31726
rect 42476 30884 42532 30940
rect 42924 31666 42980 31678
rect 42924 31614 42926 31666
rect 42978 31614 42980 31666
rect 42588 30884 42644 30894
rect 42476 30882 42644 30884
rect 42476 30830 42590 30882
rect 42642 30830 42644 30882
rect 42476 30828 42644 30830
rect 41804 30324 41860 30828
rect 41804 30258 41860 30268
rect 41916 30322 41972 30334
rect 41916 30270 41918 30322
rect 41970 30270 41972 30322
rect 41580 30146 41636 30156
rect 41468 29586 41524 29596
rect 41916 29764 41972 30270
rect 41244 29316 41300 29326
rect 41692 29316 41748 29326
rect 41244 29314 41748 29316
rect 41244 29262 41246 29314
rect 41298 29262 41694 29314
rect 41746 29262 41748 29314
rect 41244 29260 41748 29262
rect 41244 29250 41300 29260
rect 41692 28868 41748 29260
rect 40908 28812 41524 28868
rect 40908 28754 40964 28812
rect 40908 28702 40910 28754
rect 40962 28702 40964 28754
rect 40908 28690 40964 28702
rect 40348 24332 40516 24388
rect 40572 28028 40852 28084
rect 41020 28644 41076 28654
rect 40348 24276 40404 24332
rect 39900 24098 39956 24108
rect 40236 24220 40404 24276
rect 39788 23998 39790 24050
rect 39842 23998 39844 24050
rect 39788 23986 39844 23998
rect 39852 23548 40116 23558
rect 39908 23492 39956 23548
rect 40012 23492 40060 23548
rect 39852 23482 40116 23492
rect 40236 23378 40292 24220
rect 40236 23326 40238 23378
rect 40290 23326 40292 23378
rect 40236 23314 40292 23326
rect 40460 23940 40516 23950
rect 39676 23268 39732 23278
rect 39676 23174 39732 23212
rect 39788 23154 39844 23166
rect 39788 23102 39790 23154
rect 39842 23102 39844 23154
rect 39788 22932 39844 23102
rect 40124 23156 40180 23166
rect 40124 23062 40180 23100
rect 39788 22866 39844 22876
rect 39900 23044 39956 23054
rect 39676 22596 39732 22606
rect 39676 21474 39732 22540
rect 39788 22482 39844 22494
rect 39788 22430 39790 22482
rect 39842 22430 39844 22482
rect 39788 22260 39844 22430
rect 39900 22372 39956 22988
rect 40460 22594 40516 23884
rect 40460 22542 40462 22594
rect 40514 22542 40516 22594
rect 40460 22530 40516 22542
rect 39900 22278 39956 22316
rect 39788 22194 39844 22204
rect 40348 22258 40404 22270
rect 40348 22206 40350 22258
rect 40402 22206 40404 22258
rect 39852 21980 40116 21990
rect 39908 21924 39956 21980
rect 40012 21924 40060 21980
rect 39852 21914 40116 21924
rect 40348 21812 40404 22206
rect 40348 21746 40404 21756
rect 40460 21924 40516 21934
rect 39676 21422 39678 21474
rect 39730 21422 39732 21474
rect 39676 21410 39732 21422
rect 40124 21588 40180 21598
rect 40460 21588 40516 21868
rect 40124 21586 40516 21588
rect 40124 21534 40126 21586
rect 40178 21534 40516 21586
rect 40124 21532 40516 21534
rect 40124 21476 40180 21532
rect 40124 21410 40180 21420
rect 40236 20916 40292 20926
rect 40124 20692 40180 20702
rect 40124 20598 40180 20636
rect 40236 20690 40292 20860
rect 40236 20638 40238 20690
rect 40290 20638 40292 20690
rect 40236 20626 40292 20638
rect 40460 20578 40516 20590
rect 40460 20526 40462 20578
rect 40514 20526 40516 20578
rect 39852 20412 40116 20422
rect 39908 20356 39956 20412
rect 40012 20356 40060 20412
rect 39852 20346 40116 20356
rect 40460 20132 40516 20526
rect 40460 20066 40516 20076
rect 40236 20020 40292 20030
rect 40236 20018 40404 20020
rect 40236 19966 40238 20018
rect 40290 19966 40404 20018
rect 40236 19964 40404 19966
rect 40236 19954 40292 19964
rect 39852 18844 40116 18854
rect 39908 18788 39956 18844
rect 40012 18788 40060 18844
rect 39852 18778 40116 18788
rect 40012 18452 40068 18462
rect 40012 18358 40068 18396
rect 40348 18340 40404 19964
rect 40572 19684 40628 28028
rect 40684 27748 40740 27758
rect 40684 26516 40740 27692
rect 40796 27412 40852 27422
rect 40796 26850 40852 27356
rect 41020 26908 41076 28588
rect 41132 28082 41188 28812
rect 41468 28532 41524 28812
rect 41580 28756 41636 28794
rect 41580 28690 41636 28700
rect 41692 28642 41748 28812
rect 41692 28590 41694 28642
rect 41746 28590 41748 28642
rect 41692 28578 41748 28590
rect 41804 29092 41860 29102
rect 41580 28532 41636 28542
rect 41468 28530 41636 28532
rect 41468 28478 41582 28530
rect 41634 28478 41636 28530
rect 41468 28476 41636 28478
rect 41580 28466 41636 28476
rect 41132 28030 41134 28082
rect 41186 28030 41188 28082
rect 41132 28018 41188 28030
rect 41356 27970 41412 27982
rect 41356 27918 41358 27970
rect 41410 27918 41412 27970
rect 41356 27300 41412 27918
rect 41468 27860 41524 27870
rect 41468 27766 41524 27804
rect 41356 27234 41412 27244
rect 41356 27076 41412 27086
rect 41356 26962 41412 27020
rect 41356 26910 41358 26962
rect 41410 26910 41412 26962
rect 41020 26852 41188 26908
rect 40796 26798 40798 26850
rect 40850 26798 40852 26850
rect 40796 26786 40852 26798
rect 40684 26450 40740 26460
rect 40684 26292 40740 26302
rect 40684 23828 40740 26236
rect 40908 25396 40964 25406
rect 40908 25282 40964 25340
rect 40908 25230 40910 25282
rect 40962 25230 40964 25282
rect 40908 25172 40964 25230
rect 40908 25106 40964 25116
rect 40908 24836 40964 24846
rect 40908 24500 40964 24780
rect 40908 24434 40964 24444
rect 40684 23762 40740 23772
rect 40908 24164 40964 24174
rect 40796 23380 40852 23390
rect 40796 22596 40852 23324
rect 40796 22530 40852 22540
rect 40908 23154 40964 24108
rect 40908 23102 40910 23154
rect 40962 23102 40964 23154
rect 40684 22372 40740 22382
rect 40684 21812 40740 22316
rect 40908 21812 40964 23102
rect 41020 23156 41076 23166
rect 41020 22370 41076 23100
rect 41020 22318 41022 22370
rect 41074 22318 41076 22370
rect 41020 22306 41076 22318
rect 41132 22146 41188 26852
rect 41356 25620 41412 26910
rect 41692 26964 41748 27002
rect 41804 26964 41860 29036
rect 41748 26908 41860 26964
rect 41692 26898 41748 26908
rect 41916 25844 41972 29708
rect 42028 29650 42084 30828
rect 42252 30818 42308 30828
rect 42588 30818 42644 30828
rect 42028 29598 42030 29650
rect 42082 29598 42084 29650
rect 42028 29586 42084 29598
rect 42252 30660 42308 30670
rect 42252 27300 42308 30604
rect 42476 30324 42532 30334
rect 42476 29650 42532 30268
rect 42588 30212 42644 30222
rect 42588 30118 42644 30156
rect 42476 29598 42478 29650
rect 42530 29598 42532 29650
rect 42476 29586 42532 29598
rect 42924 29652 42980 31614
rect 43148 31556 43204 31566
rect 43260 31556 43316 35532
rect 44268 35588 44324 35598
rect 44268 35494 44324 35532
rect 44156 35364 44212 35374
rect 43708 34916 43764 34926
rect 43484 34804 43540 34814
rect 43484 34710 43540 34748
rect 43484 34244 43540 34254
rect 43708 34244 43764 34860
rect 44044 34804 44100 34814
rect 44044 34710 44100 34748
rect 44156 34356 44212 35308
rect 44380 35252 44436 35262
rect 44380 35138 44436 35196
rect 44380 35086 44382 35138
rect 44434 35086 44436 35138
rect 44380 35074 44436 35086
rect 44268 35028 44324 35038
rect 44268 34802 44324 34972
rect 44268 34750 44270 34802
rect 44322 34750 44324 34802
rect 44268 34738 44324 34750
rect 44156 34262 44212 34300
rect 43540 34188 43764 34244
rect 43484 34150 43540 34188
rect 44380 34132 44436 34142
rect 44268 34130 44436 34132
rect 44268 34078 44382 34130
rect 44434 34078 44436 34130
rect 44268 34076 44436 34078
rect 43484 33460 43540 33470
rect 43540 33404 43764 33460
rect 43484 33366 43540 33404
rect 43372 32562 43428 32574
rect 43372 32510 43374 32562
rect 43426 32510 43428 32562
rect 43372 32004 43428 32510
rect 43708 32562 43764 33404
rect 43932 33122 43988 33134
rect 43932 33070 43934 33122
rect 43986 33070 43988 33122
rect 43932 32788 43988 33070
rect 43932 32722 43988 32732
rect 44268 32786 44324 34076
rect 44380 34066 44436 34076
rect 44268 32734 44270 32786
rect 44322 32734 44324 32786
rect 44268 32722 44324 32734
rect 43708 32510 43710 32562
rect 43762 32510 43764 32562
rect 43708 32498 43764 32510
rect 43932 32340 43988 32350
rect 43820 32338 43988 32340
rect 43820 32286 43934 32338
rect 43986 32286 43988 32338
rect 43820 32284 43988 32286
rect 43372 31948 43764 32004
rect 43484 31668 43540 31678
rect 43484 31574 43540 31612
rect 43148 31554 43316 31556
rect 43148 31502 43150 31554
rect 43202 31502 43316 31554
rect 43148 31500 43316 31502
rect 43708 31556 43764 31948
rect 43148 31490 43204 31500
rect 43708 31490 43764 31500
rect 43708 31220 43764 31230
rect 43820 31220 43876 32284
rect 43932 32274 43988 32284
rect 43932 31556 43988 31566
rect 43932 31462 43988 31500
rect 43708 31218 43876 31220
rect 43708 31166 43710 31218
rect 43762 31166 43876 31218
rect 43708 31164 43876 31166
rect 43708 31154 43764 31164
rect 43596 30994 43652 31006
rect 43596 30942 43598 30994
rect 43650 30942 43652 30994
rect 43148 30884 43204 30894
rect 43596 30884 43652 30942
rect 43820 30996 43876 31006
rect 43820 30902 43876 30940
rect 44268 30996 44324 31006
rect 44268 30902 44324 30940
rect 43148 30882 43652 30884
rect 43148 30830 43150 30882
rect 43202 30830 43652 30882
rect 43148 30828 43652 30830
rect 43148 30772 43204 30828
rect 43148 30706 43204 30716
rect 43148 30100 43204 30110
rect 43148 29986 43204 30044
rect 43148 29934 43150 29986
rect 43202 29934 43204 29986
rect 43036 29652 43092 29662
rect 42924 29650 43092 29652
rect 42924 29598 43038 29650
rect 43090 29598 43092 29650
rect 42924 29596 43092 29598
rect 43148 29652 43204 29934
rect 43260 29876 43316 30828
rect 44380 30770 44436 30782
rect 44380 30718 44382 30770
rect 44434 30718 44436 30770
rect 43708 30324 43764 30334
rect 44380 30324 44436 30718
rect 43708 30322 44436 30324
rect 43708 30270 43710 30322
rect 43762 30270 44436 30322
rect 43708 30268 44436 30270
rect 43708 30258 43764 30268
rect 43596 30100 43652 30110
rect 43596 30006 43652 30044
rect 43820 30100 43876 30110
rect 43820 30006 43876 30044
rect 44044 29988 44100 29998
rect 44044 29894 44100 29932
rect 43260 29810 43316 29820
rect 43820 29876 43876 29886
rect 43148 29596 43652 29652
rect 43036 29586 43092 29596
rect 42364 29428 42420 29438
rect 42588 29428 42644 29438
rect 42364 29426 42588 29428
rect 42364 29374 42366 29426
rect 42418 29374 42588 29426
rect 42364 29372 42588 29374
rect 42364 29362 42420 29372
rect 42364 28868 42420 28878
rect 42364 28754 42420 28812
rect 42364 28702 42366 28754
rect 42418 28702 42420 28754
rect 42364 28690 42420 28702
rect 42588 28756 42644 29372
rect 42700 29428 42756 29438
rect 43372 29428 43428 29438
rect 42700 29426 43428 29428
rect 42700 29374 42702 29426
rect 42754 29374 43374 29426
rect 43426 29374 43428 29426
rect 42700 29372 43428 29374
rect 42700 29362 42756 29372
rect 43372 29362 43428 29372
rect 42812 28756 42868 28766
rect 42588 28754 42868 28756
rect 42588 28702 42814 28754
rect 42866 28702 42868 28754
rect 42588 28700 42868 28702
rect 42812 28690 42868 28700
rect 43484 28420 43540 28430
rect 43372 28364 43484 28420
rect 43260 28196 43316 28206
rect 43260 28084 43316 28140
rect 42812 28082 43316 28084
rect 42812 28030 43262 28082
rect 43314 28030 43316 28082
rect 42812 28028 43316 28030
rect 42700 27970 42756 27982
rect 42700 27918 42702 27970
rect 42754 27918 42756 27970
rect 42476 27860 42532 27870
rect 42476 27766 42532 27804
rect 42700 27412 42756 27918
rect 42812 27970 42868 28028
rect 43260 28018 43316 28028
rect 42812 27918 42814 27970
rect 42866 27918 42868 27970
rect 42812 27906 42868 27918
rect 42700 27356 42868 27412
rect 42364 27300 42420 27310
rect 42252 27298 42420 27300
rect 42252 27246 42366 27298
rect 42418 27246 42420 27298
rect 42252 27244 42420 27246
rect 42364 27234 42420 27244
rect 42700 27076 42756 27086
rect 41916 25778 41972 25788
rect 42252 27074 42756 27076
rect 42252 27022 42702 27074
rect 42754 27022 42756 27074
rect 42252 27020 42756 27022
rect 41356 25554 41412 25564
rect 41804 25284 41860 25294
rect 41692 25282 41860 25284
rect 41692 25230 41806 25282
rect 41858 25230 41860 25282
rect 41692 25228 41860 25230
rect 41692 25172 41748 25228
rect 41804 25218 41860 25228
rect 41356 24836 41412 24846
rect 41244 24834 41412 24836
rect 41244 24782 41358 24834
rect 41410 24782 41412 24834
rect 41244 24780 41412 24782
rect 41244 23828 41300 24780
rect 41356 24770 41412 24780
rect 41468 24724 41524 24734
rect 41692 24724 41748 25116
rect 41468 24722 41748 24724
rect 41468 24670 41470 24722
rect 41522 24670 41748 24722
rect 41468 24668 41748 24670
rect 41356 24500 41412 24510
rect 41356 24406 41412 24444
rect 41468 24276 41524 24668
rect 41804 24610 41860 24622
rect 41804 24558 41806 24610
rect 41858 24558 41860 24610
rect 41804 24388 41860 24558
rect 41804 24322 41860 24332
rect 41468 24210 41524 24220
rect 41692 23940 41748 23950
rect 41692 23846 41748 23884
rect 41244 23762 41300 23772
rect 41468 23828 41524 23838
rect 41468 23826 41636 23828
rect 41468 23774 41470 23826
rect 41522 23774 41636 23826
rect 41468 23772 41636 23774
rect 41468 23762 41524 23772
rect 41468 23380 41524 23390
rect 41468 23286 41524 23324
rect 41244 23154 41300 23166
rect 41244 23102 41246 23154
rect 41298 23102 41300 23154
rect 41244 23044 41300 23102
rect 41244 22978 41300 22988
rect 41356 23042 41412 23054
rect 41356 22990 41358 23042
rect 41410 22990 41412 23042
rect 41132 22094 41134 22146
rect 41186 22094 41188 22146
rect 41132 22082 41188 22094
rect 41020 21812 41076 21822
rect 40908 21810 41076 21812
rect 40908 21758 41022 21810
rect 41074 21758 41076 21810
rect 40908 21756 41076 21758
rect 40684 21746 40740 21756
rect 41020 21746 41076 21756
rect 41356 21700 41412 22990
rect 41580 22484 41636 23772
rect 41468 22428 41636 22484
rect 41916 23044 41972 23054
rect 41468 21700 41524 22428
rect 41692 22258 41748 22270
rect 41692 22206 41694 22258
rect 41746 22206 41748 22258
rect 41468 21644 41636 21700
rect 41356 21634 41412 21644
rect 41468 21474 41524 21486
rect 41468 21422 41470 21474
rect 41522 21422 41524 21474
rect 41468 21362 41524 21422
rect 41468 21310 41470 21362
rect 41522 21310 41524 21362
rect 41468 21140 41524 21310
rect 41244 21084 41524 21140
rect 40460 19628 40628 19684
rect 41020 20914 41076 20926
rect 41020 20862 41022 20914
rect 41074 20862 41076 20914
rect 40460 19348 40516 19628
rect 40460 19282 40516 19292
rect 40572 19460 40628 19470
rect 40572 19346 40628 19404
rect 40572 19294 40574 19346
rect 40626 19294 40628 19346
rect 40348 18246 40404 18284
rect 40348 18116 40404 18126
rect 40236 17892 40292 17902
rect 40236 17666 40292 17836
rect 40236 17614 40238 17666
rect 40290 17614 40292 17666
rect 40236 17602 40292 17614
rect 39852 17276 40116 17286
rect 39908 17220 39956 17276
rect 40012 17220 40060 17276
rect 39852 17210 40116 17220
rect 40236 17108 40292 17118
rect 40348 17108 40404 18060
rect 40572 17778 40628 19294
rect 40684 19234 40740 19246
rect 40684 19182 40686 19234
rect 40738 19182 40740 19234
rect 40684 19012 40740 19182
rect 40684 18116 40740 18956
rect 41020 18900 41076 20862
rect 41132 19572 41188 19582
rect 41244 19572 41300 21084
rect 41580 20692 41636 21644
rect 41692 21362 41748 22206
rect 41916 21924 41972 22988
rect 42140 22372 42196 22382
rect 42140 22278 42196 22316
rect 41692 21310 41694 21362
rect 41746 21310 41748 21362
rect 41692 21298 41748 21310
rect 41804 21812 41860 21822
rect 41804 20802 41860 21756
rect 41916 21810 41972 21868
rect 41916 21758 41918 21810
rect 41970 21758 41972 21810
rect 41916 21746 41972 21758
rect 41804 20750 41806 20802
rect 41858 20750 41860 20802
rect 41804 20738 41860 20750
rect 42140 21028 42196 21038
rect 41580 20636 41748 20692
rect 41468 20580 41524 20590
rect 41468 20578 41636 20580
rect 41468 20526 41470 20578
rect 41522 20526 41636 20578
rect 41468 20524 41636 20526
rect 41468 20514 41524 20524
rect 41356 20132 41412 20142
rect 41412 20076 41524 20132
rect 41356 20066 41412 20076
rect 41188 19516 41300 19572
rect 41356 19906 41412 19918
rect 41356 19854 41358 19906
rect 41410 19854 41412 19906
rect 41132 19506 41188 19516
rect 41020 18844 41300 18900
rect 40684 18050 40740 18060
rect 40796 18340 40852 18350
rect 41020 18340 41076 18350
rect 40684 17892 40740 17902
rect 40684 17798 40740 17836
rect 40572 17726 40574 17778
rect 40626 17726 40628 17778
rect 40572 17332 40628 17726
rect 40572 17266 40628 17276
rect 39788 17106 40516 17108
rect 39788 17054 40238 17106
rect 40290 17054 40516 17106
rect 39788 17052 40516 17054
rect 39676 16996 39732 17006
rect 39788 16996 39844 17052
rect 40236 17042 40292 17052
rect 39676 16994 39844 16996
rect 39676 16942 39678 16994
rect 39730 16942 39844 16994
rect 39676 16940 39844 16942
rect 39676 16658 39732 16940
rect 39676 16606 39678 16658
rect 39730 16606 39732 16658
rect 39676 16594 39732 16606
rect 40236 16322 40292 16334
rect 40236 16270 40238 16322
rect 40290 16270 40292 16322
rect 38668 14130 38724 14140
rect 38780 15092 39060 15148
rect 39116 15092 39620 15148
rect 39676 16212 39732 16222
rect 39676 15148 39732 16156
rect 39852 15708 40116 15718
rect 39908 15652 39956 15708
rect 40012 15652 40060 15708
rect 39852 15642 40116 15652
rect 40012 15540 40068 15550
rect 40012 15314 40068 15484
rect 40012 15262 40014 15314
rect 40066 15262 40068 15314
rect 40012 15250 40068 15262
rect 40236 15314 40292 16270
rect 40236 15262 40238 15314
rect 40290 15262 40292 15314
rect 39676 15092 39844 15148
rect 38668 13972 38724 13982
rect 38444 13804 38612 13860
rect 38444 13636 38500 13646
rect 38444 13542 38500 13580
rect 38220 13122 38276 13132
rect 37660 10546 37716 10556
rect 37772 11564 38052 11620
rect 38108 12628 38164 12638
rect 38108 12178 38164 12572
rect 38108 12126 38110 12178
rect 38162 12126 38164 12178
rect 37548 9774 37550 9826
rect 37602 9774 37604 9826
rect 37212 8372 37268 8988
rect 37548 8708 37604 9774
rect 37548 8642 37604 8652
rect 36988 8306 37044 8316
rect 37212 8306 37268 8316
rect 37324 8484 37380 8494
rect 37100 8148 37156 8158
rect 37100 8054 37156 8092
rect 35868 8036 35924 8046
rect 35868 8034 36596 8036
rect 35868 7982 35870 8034
rect 35922 7982 36596 8034
rect 35868 7980 36596 7982
rect 35868 7970 35924 7980
rect 35756 7756 35924 7812
rect 35756 6578 35812 6590
rect 35756 6526 35758 6578
rect 35810 6526 35812 6578
rect 35644 6356 35700 6366
rect 35644 5236 35700 6300
rect 35756 6020 35812 6526
rect 35868 6244 35924 7756
rect 36540 7586 36596 7980
rect 36540 7534 36542 7586
rect 36594 7534 36596 7586
rect 36540 7522 36596 7534
rect 37324 7474 37380 8428
rect 37324 7422 37326 7474
rect 37378 7422 37380 7474
rect 37324 7410 37380 7422
rect 37436 8258 37492 8270
rect 37436 8206 37438 8258
rect 37490 8206 37492 8258
rect 37436 7364 37492 8206
rect 37436 7298 37492 7308
rect 36092 6804 36148 6814
rect 36092 6578 36148 6748
rect 36092 6526 36094 6578
rect 36146 6526 36148 6578
rect 36092 6514 36148 6526
rect 36204 6580 36260 6590
rect 35868 6178 35924 6188
rect 36204 6132 36260 6524
rect 36204 6038 36260 6076
rect 37100 6132 37156 6142
rect 37100 6038 37156 6076
rect 37436 6132 37492 6142
rect 35812 5964 36036 6020
rect 35756 5954 35812 5964
rect 35644 5124 35700 5180
rect 35644 5068 35812 5124
rect 35308 4162 35364 4172
rect 35420 4844 35588 4900
rect 35644 4900 35700 4910
rect 32508 3444 32564 3482
rect 32508 3378 32564 3388
rect 32284 2818 32340 2828
rect 35420 2436 35476 4844
rect 35644 4806 35700 4844
rect 35756 4676 35812 5068
rect 35980 5010 36036 5964
rect 37436 6018 37492 6076
rect 37436 5966 37438 6018
rect 37490 5966 37492 6018
rect 37436 5954 37492 5966
rect 36652 5794 36708 5806
rect 36652 5742 36654 5794
rect 36706 5742 36708 5794
rect 36204 5348 36260 5358
rect 36204 5122 36260 5292
rect 36652 5348 36708 5742
rect 36708 5292 36932 5348
rect 36652 5282 36708 5292
rect 36204 5070 36206 5122
rect 36258 5070 36260 5122
rect 36204 5058 36260 5070
rect 35980 4958 35982 5010
rect 36034 4958 36036 5010
rect 35980 4946 36036 4958
rect 35532 4620 35812 4676
rect 35532 4226 35588 4620
rect 35532 4174 35534 4226
rect 35586 4174 35588 4226
rect 35532 4162 35588 4174
rect 36428 4116 36484 4126
rect 35532 3444 35588 3454
rect 36092 3444 36148 3454
rect 35532 3442 36148 3444
rect 35532 3390 35534 3442
rect 35586 3390 36094 3442
rect 36146 3390 36148 3442
rect 35532 3388 36148 3390
rect 35532 3378 35588 3388
rect 35420 2370 35476 2380
rect 35868 800 35924 3388
rect 36092 3378 36148 3388
rect 36428 3442 36484 4060
rect 36876 3666 36932 5292
rect 37436 5236 37492 5246
rect 37436 5142 37492 5180
rect 37100 5124 37156 5134
rect 37100 5030 37156 5068
rect 37772 5012 37828 11564
rect 37996 11396 38052 11406
rect 37884 11284 37940 11294
rect 37884 10834 37940 11228
rect 37996 11282 38052 11340
rect 37996 11230 37998 11282
rect 38050 11230 38052 11282
rect 37996 11218 38052 11230
rect 37884 10782 37886 10834
rect 37938 10782 37940 10834
rect 37884 10052 37940 10782
rect 38108 10836 38164 12126
rect 38220 11394 38276 11406
rect 38220 11342 38222 11394
rect 38274 11342 38276 11394
rect 38220 11284 38276 11342
rect 38220 11218 38276 11228
rect 38220 10836 38276 10846
rect 38108 10834 38276 10836
rect 38108 10782 38222 10834
rect 38274 10782 38276 10834
rect 38108 10780 38276 10782
rect 38220 10770 38276 10780
rect 38556 10388 38612 13804
rect 38668 12402 38724 13916
rect 38668 12350 38670 12402
rect 38722 12350 38724 12402
rect 38668 11956 38724 12350
rect 38668 11890 38724 11900
rect 38668 11732 38724 11742
rect 38668 10500 38724 11676
rect 38668 10406 38724 10444
rect 38556 10322 38612 10332
rect 37884 9986 37940 9996
rect 38332 9826 38388 9838
rect 38332 9774 38334 9826
rect 38386 9774 38388 9826
rect 38332 9156 38388 9774
rect 38444 9156 38500 9166
rect 38332 9154 38500 9156
rect 38332 9102 38446 9154
rect 38498 9102 38500 9154
rect 38332 9100 38500 9102
rect 37996 8930 38052 8942
rect 37996 8878 37998 8930
rect 38050 8878 38052 8930
rect 37996 8708 38052 8878
rect 37996 8642 38052 8652
rect 38332 8484 38388 9100
rect 38444 9090 38500 9100
rect 38668 9042 38724 9054
rect 38668 8990 38670 9042
rect 38722 8990 38724 9042
rect 38668 8428 38724 8990
rect 38332 8418 38388 8428
rect 38444 8372 38724 8428
rect 38220 8258 38276 8270
rect 38220 8206 38222 8258
rect 38274 8206 38276 8258
rect 38108 8146 38164 8158
rect 38108 8094 38110 8146
rect 38162 8094 38164 8146
rect 38108 6916 38164 8094
rect 38220 7924 38276 8206
rect 38220 7858 38276 7868
rect 37996 6132 38052 6142
rect 37996 6038 38052 6076
rect 37772 4946 37828 4956
rect 38108 5010 38164 6860
rect 38444 6804 38500 8372
rect 38780 8260 38836 15092
rect 38892 14308 38948 14318
rect 38892 14214 38948 14252
rect 39116 13300 39172 15092
rect 39676 14530 39732 14542
rect 39676 14478 39678 14530
rect 39730 14478 39732 14530
rect 39228 13972 39284 13982
rect 39228 13878 39284 13916
rect 39676 13972 39732 14478
rect 39788 14306 39844 15092
rect 39900 14532 39956 14542
rect 39900 14438 39956 14476
rect 39788 14254 39790 14306
rect 39842 14254 39844 14306
rect 39788 14242 39844 14254
rect 39852 14140 40116 14150
rect 39908 14084 39956 14140
rect 40012 14084 40060 14140
rect 39852 14074 40116 14084
rect 40236 13972 40292 15262
rect 40348 15204 40404 15242
rect 40348 15138 40404 15148
rect 39676 13916 40292 13972
rect 38220 5124 38276 5134
rect 38220 5030 38276 5068
rect 38108 4958 38110 5010
rect 38162 4958 38164 5010
rect 38108 4946 38164 4958
rect 37660 4900 37716 4910
rect 37660 4450 37716 4844
rect 37660 4398 37662 4450
rect 37714 4398 37716 4450
rect 37660 4386 37716 4398
rect 38444 4338 38500 6748
rect 38668 8204 38836 8260
rect 38892 13244 39172 13300
rect 38668 6020 38724 8204
rect 38780 8034 38836 8046
rect 38780 7982 38782 8034
rect 38834 7982 38836 8034
rect 38780 7924 38836 7982
rect 38780 7140 38836 7868
rect 38780 7074 38836 7084
rect 38892 6692 38948 13244
rect 39116 13076 39172 13086
rect 39116 12982 39172 13020
rect 39340 13076 39396 13086
rect 39340 12628 39396 13020
rect 39340 12562 39396 12572
rect 39452 12964 39508 12974
rect 39452 12402 39508 12908
rect 39676 12962 39732 13916
rect 39676 12910 39678 12962
rect 39730 12910 39732 12962
rect 39676 12898 39732 12910
rect 40012 13634 40068 13646
rect 40012 13582 40014 13634
rect 40066 13582 40068 13634
rect 40012 12740 40068 13582
rect 40124 13524 40180 13534
rect 40124 13522 40404 13524
rect 40124 13470 40126 13522
rect 40178 13470 40404 13522
rect 40124 13468 40404 13470
rect 40124 13458 40180 13468
rect 40348 12962 40404 13468
rect 40348 12910 40350 12962
rect 40402 12910 40404 12962
rect 40348 12898 40404 12910
rect 40012 12674 40068 12684
rect 39852 12572 40116 12582
rect 39908 12516 39956 12572
rect 40012 12516 40060 12572
rect 39852 12506 40116 12516
rect 39452 12350 39454 12402
rect 39506 12350 39508 12402
rect 39452 12338 39508 12350
rect 39900 12404 39956 12414
rect 39004 12290 39060 12302
rect 39004 12238 39006 12290
rect 39058 12238 39060 12290
rect 39004 12068 39060 12238
rect 39900 12178 39956 12348
rect 39900 12126 39902 12178
rect 39954 12126 39956 12178
rect 39004 12002 39060 12012
rect 39340 12066 39396 12078
rect 39340 12014 39342 12066
rect 39394 12014 39396 12066
rect 39004 11508 39060 11518
rect 39004 11414 39060 11452
rect 39340 11284 39396 12014
rect 39900 11508 39956 12126
rect 40124 12290 40180 12302
rect 40124 12238 40126 12290
rect 40178 12238 40180 12290
rect 40012 11508 40068 11518
rect 39900 11506 40068 11508
rect 39900 11454 40014 11506
rect 40066 11454 40068 11506
rect 39900 11452 40068 11454
rect 40012 11442 40068 11452
rect 40124 11508 40180 12238
rect 40124 11442 40180 11452
rect 40348 12292 40404 12302
rect 40348 11506 40404 12236
rect 40348 11454 40350 11506
rect 40402 11454 40404 11506
rect 40348 11442 40404 11454
rect 39340 10724 39396 11228
rect 39452 11170 39508 11182
rect 39452 11118 39454 11170
rect 39506 11118 39508 11170
rect 39452 11060 39508 11118
rect 39452 10994 39508 11004
rect 39852 11004 40116 11014
rect 39908 10948 39956 11004
rect 40012 10948 40060 11004
rect 39852 10938 40116 10948
rect 39340 10658 39396 10668
rect 39676 10722 39732 10734
rect 39676 10670 39678 10722
rect 39730 10670 39732 10722
rect 39676 10500 39732 10670
rect 40012 10724 40068 10734
rect 40012 10630 40068 10668
rect 39676 10434 39732 10444
rect 39116 10388 39172 10398
rect 39116 10386 39396 10388
rect 39116 10334 39118 10386
rect 39170 10334 39396 10386
rect 39116 10332 39396 10334
rect 39116 10322 39172 10332
rect 39116 9714 39172 9726
rect 39116 9662 39118 9714
rect 39170 9662 39172 9714
rect 39116 9266 39172 9662
rect 39116 9214 39118 9266
rect 39170 9214 39172 9266
rect 39116 9202 39172 9214
rect 39340 9042 39396 10332
rect 39340 8990 39342 9042
rect 39394 8990 39396 9042
rect 39340 8978 39396 8990
rect 39452 10386 39508 10398
rect 39452 10334 39454 10386
rect 39506 10334 39508 10386
rect 39452 7476 39508 10334
rect 39852 9436 40116 9446
rect 39908 9380 39956 9436
rect 40012 9380 40060 9436
rect 39852 9370 40116 9380
rect 39452 7382 39508 7420
rect 39564 8146 39620 8158
rect 39564 8094 39566 8146
rect 39618 8094 39620 8146
rect 39116 7252 39172 7262
rect 39564 7252 39620 8094
rect 40460 8148 40516 17052
rect 40796 16996 40852 18284
rect 40796 16930 40852 16940
rect 40908 18338 41076 18340
rect 40908 18286 41022 18338
rect 41074 18286 41076 18338
rect 40908 18284 41076 18286
rect 40908 16772 40964 18284
rect 41020 18274 41076 18284
rect 41020 18116 41076 18126
rect 41020 17666 41076 18060
rect 41244 18004 41300 18844
rect 41244 17938 41300 17948
rect 41020 17614 41022 17666
rect 41074 17614 41076 17666
rect 41020 17556 41076 17614
rect 41020 17500 41300 17556
rect 41020 17332 41076 17342
rect 41076 17276 41188 17332
rect 41020 17266 41076 17276
rect 41020 16996 41076 17006
rect 41020 16902 41076 16940
rect 40460 8082 40516 8092
rect 40572 16716 40964 16772
rect 40572 8370 40628 16716
rect 40684 16324 40740 16334
rect 40684 15148 40740 16268
rect 41132 16210 41188 17276
rect 41132 16158 41134 16210
rect 41186 16158 41188 16210
rect 41132 16146 41188 16158
rect 41244 16098 41300 17500
rect 41244 16046 41246 16098
rect 41298 16046 41300 16098
rect 41244 16034 41300 16046
rect 41020 15876 41076 15886
rect 40908 15314 40964 15326
rect 40908 15262 40910 15314
rect 40962 15262 40964 15314
rect 40908 15148 40964 15262
rect 41020 15316 41076 15820
rect 41356 15428 41412 19854
rect 41468 19122 41524 20076
rect 41468 19070 41470 19122
rect 41522 19070 41524 19122
rect 41468 19058 41524 19070
rect 41580 19012 41636 20524
rect 41580 18918 41636 18956
rect 41692 19348 41748 20636
rect 41916 20018 41972 20030
rect 41916 19966 41918 20018
rect 41970 19966 41972 20018
rect 41916 19796 41972 19966
rect 42028 19796 42084 19806
rect 41916 19740 42028 19796
rect 41468 18452 41524 18462
rect 41468 17106 41524 18396
rect 41468 17054 41470 17106
rect 41522 17054 41524 17106
rect 41468 17042 41524 17054
rect 41244 15372 41412 15428
rect 41132 15316 41188 15326
rect 41020 15314 41188 15316
rect 41020 15262 41134 15314
rect 41186 15262 41188 15314
rect 41020 15260 41188 15262
rect 41132 15250 41188 15260
rect 41244 15148 41300 15372
rect 40684 15092 40964 15148
rect 40908 14642 40964 15092
rect 40908 14590 40910 14642
rect 40962 14590 40964 14642
rect 40908 14578 40964 14590
rect 41132 15092 41300 15148
rect 41020 14532 41076 14542
rect 41020 14438 41076 14476
rect 40572 8318 40574 8370
rect 40626 8318 40628 8370
rect 39900 8036 39956 8046
rect 39116 7250 39620 7252
rect 39116 7198 39118 7250
rect 39170 7198 39620 7250
rect 39116 7196 39620 7198
rect 39676 8034 39956 8036
rect 39676 7982 39902 8034
rect 39954 7982 39956 8034
rect 39676 7980 39956 7982
rect 39116 7186 39172 7196
rect 39676 6802 39732 7980
rect 39900 7970 39956 7980
rect 39852 7868 40116 7878
rect 39908 7812 39956 7868
rect 40012 7812 40060 7868
rect 39852 7802 40116 7812
rect 40124 7588 40180 7598
rect 40124 7494 40180 7532
rect 40236 7476 40292 7486
rect 40572 7476 40628 8318
rect 40236 7474 40628 7476
rect 40236 7422 40238 7474
rect 40290 7422 40628 7474
rect 40236 7420 40628 7422
rect 40684 14420 40740 14430
rect 40236 7028 40292 7420
rect 40236 6962 40292 6972
rect 39676 6750 39678 6802
rect 39730 6750 39732 6802
rect 39676 6738 39732 6750
rect 38892 6626 38948 6636
rect 39004 6690 39060 6702
rect 39004 6638 39006 6690
rect 39058 6638 39060 6690
rect 38444 4286 38446 4338
rect 38498 4286 38500 4338
rect 38444 4274 38500 4286
rect 38556 5964 38724 6020
rect 38556 3780 38612 5964
rect 39004 5908 39060 6638
rect 39852 6300 40116 6310
rect 39908 6244 39956 6300
rect 40012 6244 40060 6300
rect 39852 6234 40116 6244
rect 38668 5794 38724 5806
rect 38668 5742 38670 5794
rect 38722 5742 38724 5794
rect 38668 5124 38724 5742
rect 38668 4452 38724 5068
rect 39004 5122 39060 5852
rect 40684 5124 40740 14364
rect 40908 13860 40964 13870
rect 40908 13766 40964 13804
rect 41132 12964 41188 15092
rect 41580 14418 41636 14430
rect 41580 14366 41582 14418
rect 41634 14366 41636 14418
rect 41580 14308 41636 14366
rect 41692 14420 41748 19292
rect 42028 18452 42084 19740
rect 42028 18358 42084 18396
rect 42140 19234 42196 20972
rect 42252 19572 42308 27020
rect 42700 27010 42756 27020
rect 42700 26516 42756 26554
rect 42700 26450 42756 26460
rect 42476 26292 42532 26302
rect 42700 26292 42756 26302
rect 42812 26292 42868 27356
rect 43372 26964 43428 28364
rect 43484 28354 43540 28364
rect 43484 27076 43540 27086
rect 43484 26982 43540 27020
rect 43372 26898 43428 26908
rect 42476 26290 42644 26292
rect 42476 26238 42478 26290
rect 42530 26238 42644 26290
rect 42476 26236 42644 26238
rect 42476 26226 42532 26236
rect 42476 24724 42532 24734
rect 42476 24630 42532 24668
rect 42588 24164 42644 26236
rect 42700 26290 42868 26292
rect 42700 26238 42702 26290
rect 42754 26238 42868 26290
rect 42700 26236 42868 26238
rect 42700 26226 42756 26236
rect 42700 24610 42756 24622
rect 42700 24558 42702 24610
rect 42754 24558 42756 24610
rect 42700 24276 42756 24558
rect 42700 24210 42756 24220
rect 42588 23940 42644 24108
rect 42700 23940 42756 23950
rect 42588 23938 42756 23940
rect 42588 23886 42702 23938
rect 42754 23886 42756 23938
rect 42588 23884 42756 23886
rect 42588 23548 42644 23884
rect 42700 23874 42756 23884
rect 42812 23940 42868 26236
rect 43036 26290 43092 26302
rect 43036 26238 43038 26290
rect 43090 26238 43092 26290
rect 43036 26180 43092 26238
rect 43484 26180 43540 26190
rect 43036 26178 43540 26180
rect 43036 26126 43486 26178
rect 43538 26126 43540 26178
rect 43036 26124 43540 26126
rect 43372 25956 43428 25966
rect 43372 25396 43428 25900
rect 43484 25620 43540 26124
rect 43484 25554 43540 25564
rect 43596 25396 43652 29596
rect 43820 28196 43876 29820
rect 43932 29538 43988 29550
rect 43932 29486 43934 29538
rect 43986 29486 43988 29538
rect 43932 29428 43988 29486
rect 43988 29372 44100 29428
rect 43932 29362 43988 29372
rect 43372 25340 43652 25396
rect 43708 28140 43876 28196
rect 43708 25396 43764 28140
rect 43932 28084 43988 28094
rect 43820 28028 43932 28084
rect 43820 25956 43876 28028
rect 43932 27990 43988 28028
rect 43932 26962 43988 26974
rect 43932 26910 43934 26962
rect 43986 26910 43988 26962
rect 43932 26908 43988 26910
rect 44044 26908 44100 29372
rect 44156 29426 44212 29438
rect 44156 29374 44158 29426
rect 44210 29374 44212 29426
rect 44156 28082 44212 29374
rect 44156 28030 44158 28082
rect 44210 28030 44212 28082
rect 44156 28018 44212 28030
rect 44268 29316 44324 29326
rect 44268 27860 44324 29260
rect 44380 28084 44436 28094
rect 44492 28084 44548 37212
rect 46956 36932 47012 39228
rect 48384 39200 48496 40000
rect 50848 39200 50960 40000
rect 53312 39200 53424 40000
rect 55776 39200 55888 40000
rect 58240 39200 58352 40000
rect 60704 39200 60816 40000
rect 63168 39200 63280 40000
rect 65632 39200 65744 40000
rect 68096 39200 68208 40000
rect 70560 39200 70672 40000
rect 73024 39200 73136 40000
rect 75488 39200 75600 40000
rect 77952 39200 78064 40000
rect 46956 36876 47684 36932
rect 47628 36706 47684 36876
rect 47628 36654 47630 36706
rect 47682 36654 47684 36706
rect 47628 36642 47684 36654
rect 45836 36484 45892 36494
rect 45052 35698 45108 35710
rect 45052 35646 45054 35698
rect 45106 35646 45108 35698
rect 44940 35028 44996 35038
rect 44940 34934 44996 34972
rect 45052 34692 45108 35646
rect 45612 35586 45668 35598
rect 45612 35534 45614 35586
rect 45666 35534 45668 35586
rect 45164 35476 45220 35486
rect 45220 35420 45332 35476
rect 45164 35410 45220 35420
rect 45164 34692 45220 34702
rect 45052 34636 45164 34692
rect 44716 34244 44772 34254
rect 44716 34150 44772 34188
rect 45164 34130 45220 34636
rect 45164 34078 45166 34130
rect 45218 34078 45220 34130
rect 45164 34066 45220 34078
rect 44828 33460 44884 33470
rect 44828 33366 44884 33404
rect 45052 33348 45108 33358
rect 44940 33346 45108 33348
rect 44940 33294 45054 33346
rect 45106 33294 45108 33346
rect 44940 33292 45108 33294
rect 44940 32900 44996 33292
rect 45052 33282 45108 33292
rect 44716 32844 44996 32900
rect 44604 31108 44660 31118
rect 44604 31014 44660 31052
rect 44716 30770 44772 32844
rect 45276 32788 45332 35420
rect 45500 35474 45556 35486
rect 45500 35422 45502 35474
rect 45554 35422 45556 35474
rect 45388 35028 45444 35038
rect 45388 34934 45444 34972
rect 45388 33460 45444 33470
rect 45388 33366 45444 33404
rect 44828 32676 44884 32686
rect 45164 32676 45220 32686
rect 45276 32676 45332 32732
rect 44828 32674 45108 32676
rect 44828 32622 44830 32674
rect 44882 32622 45108 32674
rect 44828 32620 45108 32622
rect 44828 32610 44884 32620
rect 44828 32452 44884 32462
rect 44828 32002 44884 32396
rect 44828 31950 44830 32002
rect 44882 31950 44884 32002
rect 44828 31938 44884 31950
rect 44940 31666 44996 31678
rect 44940 31614 44942 31666
rect 44994 31614 44996 31666
rect 44940 31556 44996 31614
rect 45052 31668 45108 32620
rect 45164 32674 45332 32676
rect 45164 32622 45166 32674
rect 45218 32622 45332 32674
rect 45164 32620 45332 32622
rect 45164 32452 45220 32620
rect 45164 32386 45220 32396
rect 45500 32004 45556 35422
rect 45612 35252 45668 35534
rect 45612 35186 45668 35196
rect 45724 35028 45780 35038
rect 45612 34972 45724 35028
rect 45612 34914 45668 34972
rect 45724 34962 45780 34972
rect 45612 34862 45614 34914
rect 45666 34862 45668 34914
rect 45612 34804 45668 34862
rect 45612 34738 45668 34748
rect 45724 34802 45780 34814
rect 45724 34750 45726 34802
rect 45778 34750 45780 34802
rect 45724 34580 45780 34750
rect 45836 34804 45892 36428
rect 46284 36482 46340 36494
rect 46284 36430 46286 36482
rect 46338 36430 46340 36482
rect 46284 36260 46340 36430
rect 46284 36194 46340 36204
rect 46844 36258 46900 36270
rect 46844 36206 46846 36258
rect 46898 36206 46900 36258
rect 46284 35924 46340 35934
rect 46284 35700 46340 35868
rect 46844 35924 46900 36206
rect 46844 35858 46900 35868
rect 48188 35812 48244 35822
rect 48188 35718 48244 35756
rect 46060 35698 46340 35700
rect 46060 35646 46286 35698
rect 46338 35646 46340 35698
rect 46060 35644 46340 35646
rect 45948 34916 46004 34926
rect 45948 34822 46004 34860
rect 45836 34738 45892 34748
rect 46060 34580 46116 35644
rect 46284 35634 46340 35644
rect 47628 35700 47684 35710
rect 46956 35588 47012 35598
rect 46844 35586 47012 35588
rect 46844 35534 46958 35586
rect 47010 35534 47012 35586
rect 46844 35532 47012 35534
rect 45724 34524 46116 34580
rect 46172 35364 46228 35374
rect 45724 34356 45780 34524
rect 45724 34290 45780 34300
rect 45836 34244 45892 34254
rect 45836 34150 45892 34188
rect 45836 33348 45892 33358
rect 45836 33254 45892 33292
rect 45612 32788 45668 32798
rect 45612 32694 45668 32732
rect 46172 32564 46228 35308
rect 46396 35028 46452 35038
rect 46396 34934 46452 34972
rect 46732 34916 46788 34926
rect 46844 34916 46900 35532
rect 46956 35522 47012 35532
rect 46788 34860 46900 34916
rect 47628 35028 47684 35644
rect 47964 35698 48020 35710
rect 47964 35646 47966 35698
rect 48018 35646 48020 35698
rect 47628 34914 47684 34972
rect 47628 34862 47630 34914
rect 47682 34862 47684 34914
rect 46732 34850 46788 34860
rect 47628 34850 47684 34862
rect 47740 35586 47796 35598
rect 47740 35534 47742 35586
rect 47794 35534 47796 35586
rect 46956 34804 47012 34814
rect 46844 34802 47012 34804
rect 46844 34750 46958 34802
rect 47010 34750 47012 34802
rect 46844 34748 47012 34750
rect 46284 33122 46340 33134
rect 46284 33070 46286 33122
rect 46338 33070 46340 33122
rect 46284 32788 46340 33070
rect 46284 32694 46340 32732
rect 46620 32674 46676 32686
rect 46620 32622 46622 32674
rect 46674 32622 46676 32674
rect 46172 32508 46340 32564
rect 45052 31602 45108 31612
rect 45164 31948 45556 32004
rect 44940 31490 44996 31500
rect 44716 30718 44718 30770
rect 44770 30718 44772 30770
rect 44716 30706 44772 30718
rect 44940 29986 44996 29998
rect 44940 29934 44942 29986
rect 44994 29934 44996 29986
rect 44940 29876 44996 29934
rect 44716 29428 44772 29438
rect 44716 29334 44772 29372
rect 44940 29204 44996 29820
rect 44940 29138 44996 29148
rect 44940 28756 44996 28766
rect 44436 28028 44660 28084
rect 44380 27990 44436 28028
rect 43932 26852 44100 26908
rect 44156 27804 44324 27860
rect 44492 27858 44548 27870
rect 44492 27806 44494 27858
rect 44546 27806 44548 27858
rect 44156 26908 44212 27804
rect 44492 27748 44548 27806
rect 44492 27682 44548 27692
rect 44492 27412 44548 27422
rect 44268 27356 44492 27412
rect 44268 27074 44324 27356
rect 44492 27346 44548 27356
rect 44268 27022 44270 27074
rect 44322 27022 44324 27074
rect 44268 27010 44324 27022
rect 44156 26852 44436 26908
rect 43932 26180 43988 26852
rect 43988 26124 44324 26180
rect 43932 26114 43988 26124
rect 43820 25618 43876 25900
rect 43820 25566 43822 25618
rect 43874 25566 43876 25618
rect 43820 25554 43876 25566
rect 44268 25618 44324 26124
rect 44268 25566 44270 25618
rect 44322 25566 44324 25618
rect 44268 25508 44324 25566
rect 44268 25442 44324 25452
rect 43708 25340 43988 25396
rect 43036 24724 43092 24734
rect 42924 23940 42980 23950
rect 42812 23938 42980 23940
rect 42812 23886 42926 23938
rect 42978 23886 42980 23938
rect 42812 23884 42980 23886
rect 42812 23604 42868 23884
rect 42924 23874 42980 23884
rect 43036 23940 43092 24668
rect 43260 24610 43316 24622
rect 43260 24558 43262 24610
rect 43314 24558 43316 24610
rect 43260 24276 43316 24558
rect 43260 24210 43316 24220
rect 43036 23714 43092 23884
rect 43036 23662 43038 23714
rect 43090 23662 43092 23714
rect 43036 23650 43092 23662
rect 43260 23826 43316 23838
rect 43260 23774 43262 23826
rect 43314 23774 43316 23826
rect 42364 23492 42644 23548
rect 42700 23548 42868 23604
rect 43260 23604 43316 23774
rect 43372 23604 43428 23614
rect 43260 23548 43372 23604
rect 42364 23266 42420 23492
rect 42364 23214 42366 23266
rect 42418 23214 42420 23266
rect 42364 23202 42420 23214
rect 42476 23268 42532 23278
rect 42476 22370 42532 23212
rect 42476 22318 42478 22370
rect 42530 22318 42532 22370
rect 42476 22306 42532 22318
rect 42700 23154 42756 23548
rect 43372 23538 43428 23548
rect 42812 23380 42868 23390
rect 42812 23286 42868 23324
rect 42700 23102 42702 23154
rect 42754 23102 42756 23154
rect 42700 22260 42756 23102
rect 43036 23154 43092 23166
rect 43036 23102 43038 23154
rect 43090 23102 43092 23154
rect 43036 23044 43092 23102
rect 43372 23044 43428 23054
rect 43036 23042 43428 23044
rect 43036 22990 43374 23042
rect 43426 22990 43428 23042
rect 43036 22988 43428 22990
rect 43372 22596 43428 22988
rect 43372 22530 43428 22540
rect 43260 22372 43316 22382
rect 43260 22278 43316 22316
rect 42812 22260 42868 22270
rect 42700 22258 42868 22260
rect 42700 22206 42814 22258
rect 42866 22206 42868 22258
rect 42700 22204 42868 22206
rect 42812 22194 42868 22204
rect 42364 21812 42420 21822
rect 42364 21718 42420 21756
rect 42812 21588 42868 21598
rect 42812 21494 42868 21532
rect 43372 21588 43428 21598
rect 43484 21588 43540 25340
rect 43708 23940 43764 23950
rect 43708 23846 43764 23884
rect 43596 23828 43652 23838
rect 43596 23734 43652 23772
rect 43820 23044 43876 23054
rect 43708 22988 43820 23044
rect 43708 22148 43764 22988
rect 43820 22950 43876 22988
rect 43708 22054 43764 22092
rect 43596 21588 43652 21598
rect 43484 21586 43652 21588
rect 43484 21534 43598 21586
rect 43650 21534 43652 21586
rect 43484 21532 43652 21534
rect 43372 21494 43428 21532
rect 42700 21028 42756 21038
rect 42700 20914 42756 20972
rect 42700 20862 42702 20914
rect 42754 20862 42756 20914
rect 42700 20850 42756 20862
rect 43596 20914 43652 21532
rect 43932 21588 43988 25340
rect 44156 25172 44212 25182
rect 44044 24612 44100 24622
rect 44044 24052 44100 24556
rect 44044 23986 44100 23996
rect 44156 24050 44212 25116
rect 44156 23998 44158 24050
rect 44210 23998 44212 24050
rect 44156 23604 44212 23998
rect 44156 23538 44212 23548
rect 44380 23380 44436 26852
rect 44604 26514 44660 28028
rect 44940 27186 44996 28700
rect 44940 27134 44942 27186
rect 44994 27134 44996 27186
rect 44940 27122 44996 27134
rect 45052 27746 45108 27758
rect 45052 27694 45054 27746
rect 45106 27694 45108 27746
rect 44828 26964 44884 27002
rect 44828 26740 44884 26908
rect 44828 26674 44884 26684
rect 45052 26850 45108 27694
rect 45052 26798 45054 26850
rect 45106 26798 45108 26850
rect 45052 26516 45108 26798
rect 44604 26462 44606 26514
rect 44658 26462 44660 26514
rect 44604 26450 44660 26462
rect 44828 26460 45108 26516
rect 45164 27412 45220 31948
rect 46172 31892 46228 31902
rect 46172 31798 46228 31836
rect 45388 31556 45444 31566
rect 45388 31220 45444 31500
rect 45388 31154 45444 31164
rect 45276 29986 45332 29998
rect 45276 29934 45278 29986
rect 45330 29934 45332 29986
rect 45276 29540 45332 29934
rect 45724 29986 45780 29998
rect 45724 29934 45726 29986
rect 45778 29934 45780 29986
rect 45724 29876 45780 29934
rect 45724 29810 45780 29820
rect 46060 29988 46116 29998
rect 45276 29474 45332 29484
rect 45948 29316 46004 29326
rect 45948 29222 46004 29260
rect 46060 28754 46116 29932
rect 46172 29540 46228 29550
rect 46172 29446 46228 29484
rect 46060 28702 46062 28754
rect 46114 28702 46116 28754
rect 46060 28690 46116 28702
rect 46060 28418 46116 28430
rect 46060 28366 46062 28418
rect 46114 28366 46116 28418
rect 45388 27748 45444 27758
rect 45388 27412 45444 27692
rect 45388 27356 45668 27412
rect 44828 26292 44884 26460
rect 45164 26402 45220 27356
rect 45500 26964 45556 27002
rect 45612 26964 45668 27356
rect 45836 26964 45892 27002
rect 45612 26908 45836 26964
rect 45500 26898 45556 26908
rect 45836 26898 45892 26908
rect 46060 26628 46116 28366
rect 46172 28418 46228 28430
rect 46172 28366 46174 28418
rect 46226 28366 46228 28418
rect 46172 27972 46228 28366
rect 46172 27906 46228 27916
rect 46284 27636 46340 32508
rect 46620 31780 46676 32622
rect 46620 31714 46676 31724
rect 46732 31556 46788 31566
rect 46732 31462 46788 31500
rect 46844 31220 46900 34748
rect 46956 34738 47012 34748
rect 47740 33572 47796 35534
rect 47964 35476 48020 35646
rect 47964 34914 48020 35420
rect 48412 35140 48468 39200
rect 49512 36876 49776 36886
rect 49568 36820 49616 36876
rect 49672 36820 49720 36876
rect 49512 36810 49776 36820
rect 49868 36482 49924 36494
rect 49868 36430 49870 36482
rect 49922 36430 49924 36482
rect 48972 35812 49028 35822
rect 48972 35718 49028 35756
rect 48860 35698 48916 35710
rect 48860 35646 48862 35698
rect 48914 35646 48916 35698
rect 48860 35476 48916 35646
rect 49084 35700 49140 35710
rect 49084 35606 49140 35644
rect 49532 35476 49588 35486
rect 48860 35410 48916 35420
rect 49308 35474 49588 35476
rect 49308 35422 49534 35474
rect 49586 35422 49588 35474
rect 49308 35420 49588 35422
rect 48412 35074 48468 35084
rect 47964 34862 47966 34914
rect 48018 34862 48020 34914
rect 47964 34850 48020 34862
rect 49196 34914 49252 34926
rect 49196 34862 49198 34914
rect 49250 34862 49252 34914
rect 49196 34692 49252 34862
rect 49196 34626 49252 34636
rect 48076 34468 48132 34478
rect 48076 34354 48132 34412
rect 48076 34302 48078 34354
rect 48130 34302 48132 34354
rect 48076 34290 48132 34302
rect 47740 33506 47796 33516
rect 48748 34018 48804 34030
rect 48748 33966 48750 34018
rect 48802 33966 48804 34018
rect 48524 32004 48580 32014
rect 47964 31892 48020 31902
rect 46620 31164 46900 31220
rect 47516 31556 47572 31566
rect 46396 28644 46452 28654
rect 46620 28644 46676 31164
rect 46844 30996 46900 31006
rect 46844 30322 46900 30940
rect 47516 30994 47572 31500
rect 47516 30942 47518 30994
rect 47570 30942 47572 30994
rect 47516 30436 47572 30942
rect 47964 30884 48020 31836
rect 47964 30790 48020 30828
rect 46844 30270 46846 30322
rect 46898 30270 46900 30322
rect 46844 30258 46900 30270
rect 47068 30380 47572 30436
rect 46844 29986 46900 29998
rect 46844 29934 46846 29986
rect 46898 29934 46900 29986
rect 46396 28530 46452 28588
rect 46396 28478 46398 28530
rect 46450 28478 46452 28530
rect 46396 28466 46452 28478
rect 46508 28642 46676 28644
rect 46508 28590 46622 28642
rect 46674 28590 46676 28642
rect 46508 28588 46676 28590
rect 46284 27570 46340 27580
rect 46060 26572 46340 26628
rect 46284 26514 46340 26572
rect 46284 26462 46286 26514
rect 46338 26462 46340 26514
rect 46284 26450 46340 26462
rect 45164 26350 45166 26402
rect 45218 26350 45220 26402
rect 45164 26338 45220 26350
rect 44604 26236 44884 26292
rect 45052 26290 45108 26302
rect 45052 26238 45054 26290
rect 45106 26238 45108 26290
rect 44604 23548 44660 26236
rect 45052 25956 45108 26238
rect 45276 26292 45332 26302
rect 46060 26292 46116 26302
rect 46508 26292 46564 28588
rect 46620 28578 46676 28588
rect 46732 29428 46788 29438
rect 46732 27972 46788 29372
rect 46844 28756 46900 29934
rect 46956 29988 47012 29998
rect 46956 29316 47012 29932
rect 46956 29250 47012 29260
rect 46844 28690 46900 28700
rect 46956 28980 47012 28990
rect 46956 28084 47012 28924
rect 46956 28018 47012 28028
rect 46732 27916 46900 27972
rect 46844 27860 46900 27916
rect 46956 27860 47012 27870
rect 46844 27858 47012 27860
rect 46844 27806 46958 27858
rect 47010 27806 47012 27858
rect 46844 27804 47012 27806
rect 46956 27794 47012 27804
rect 46956 27636 47012 27646
rect 45276 26290 45444 26292
rect 45276 26238 45278 26290
rect 45330 26238 45444 26290
rect 45276 26236 45444 26238
rect 45276 26226 45332 26236
rect 45108 25900 45220 25956
rect 45052 25890 45108 25900
rect 44940 25844 44996 25854
rect 44828 25508 44884 25518
rect 44828 25414 44884 25452
rect 44940 25284 44996 25788
rect 45164 25506 45220 25900
rect 45164 25454 45166 25506
rect 45218 25454 45220 25506
rect 45164 25442 45220 25454
rect 45388 25506 45444 26236
rect 45612 26290 46116 26292
rect 45612 26238 46062 26290
rect 46114 26238 46116 26290
rect 45612 26236 46116 26238
rect 45612 25844 45668 26236
rect 46060 26226 46116 26236
rect 46172 26236 46564 26292
rect 46844 27076 46900 27086
rect 45724 26068 45780 26078
rect 45724 25974 45780 26012
rect 45612 25778 45668 25788
rect 45388 25454 45390 25506
rect 45442 25454 45444 25506
rect 45052 25284 45108 25294
rect 44940 25282 45108 25284
rect 44940 25230 45054 25282
rect 45106 25230 45108 25282
rect 44940 25228 45108 25230
rect 45052 25218 45108 25228
rect 45388 24834 45444 25454
rect 45948 25284 46004 25294
rect 45388 24782 45390 24834
rect 45442 24782 45444 24834
rect 45388 24770 45444 24782
rect 45836 24834 45892 24846
rect 45836 24782 45838 24834
rect 45890 24782 45892 24834
rect 44716 24722 44772 24734
rect 44716 24670 44718 24722
rect 44770 24670 44772 24722
rect 44716 24612 44772 24670
rect 44716 24546 44772 24556
rect 45276 24724 45332 24734
rect 44380 23314 44436 23324
rect 44492 23492 44660 23548
rect 43932 21522 43988 21532
rect 44268 22372 44324 22382
rect 44492 22372 44548 23492
rect 44268 22370 44548 22372
rect 44268 22318 44270 22370
rect 44322 22318 44548 22370
rect 44268 22316 44548 22318
rect 44604 23042 44660 23054
rect 44604 22990 44606 23042
rect 44658 22990 44660 23042
rect 44604 22708 44660 22990
rect 45052 23044 45108 23054
rect 45052 23042 45220 23044
rect 45052 22990 45054 23042
rect 45106 22990 45220 23042
rect 45052 22988 45220 22990
rect 45052 22978 45108 22988
rect 45164 22708 45220 22988
rect 44604 22652 45108 22708
rect 43596 20862 43598 20914
rect 43650 20862 43652 20914
rect 43596 20850 43652 20862
rect 44156 21362 44212 21374
rect 44156 21310 44158 21362
rect 44210 21310 44212 21362
rect 42364 20802 42420 20814
rect 42364 20750 42366 20802
rect 42418 20750 42420 20802
rect 42364 20356 42420 20750
rect 43036 20690 43092 20702
rect 43036 20638 43038 20690
rect 43090 20638 43092 20690
rect 43036 20580 43092 20638
rect 43036 20514 43092 20524
rect 43932 20580 43988 20590
rect 42364 20300 42980 20356
rect 42476 20132 42532 20142
rect 42700 20132 42756 20142
rect 42476 20038 42532 20076
rect 42588 20076 42700 20132
rect 42364 19572 42420 19582
rect 42252 19516 42364 19572
rect 42364 19506 42420 19516
rect 42140 19182 42142 19234
rect 42194 19182 42196 19234
rect 42028 16996 42084 17006
rect 42140 16996 42196 19182
rect 42252 19236 42308 19246
rect 42308 19180 42420 19236
rect 42252 19170 42308 19180
rect 42364 18116 42420 19180
rect 42588 19234 42644 20076
rect 42700 20038 42756 20076
rect 42588 19182 42590 19234
rect 42642 19182 42644 19234
rect 42476 19012 42532 19022
rect 42476 18674 42532 18956
rect 42476 18622 42478 18674
rect 42530 18622 42532 18674
rect 42476 18610 42532 18622
rect 42364 18060 42532 18116
rect 42028 16994 42196 16996
rect 42028 16942 42030 16994
rect 42082 16942 42196 16994
rect 42028 16940 42196 16942
rect 42476 17220 42532 18060
rect 42476 16994 42532 17164
rect 42476 16942 42478 16994
rect 42530 16942 42532 16994
rect 42028 16930 42084 16940
rect 42476 16930 42532 16942
rect 42588 16996 42644 19182
rect 42812 19794 42868 19806
rect 42812 19742 42814 19794
rect 42866 19742 42868 19794
rect 41804 16882 41860 16894
rect 42364 16884 42420 16894
rect 41804 16830 41806 16882
rect 41858 16830 41860 16882
rect 41804 16772 41860 16830
rect 41804 16210 41860 16716
rect 41804 16158 41806 16210
rect 41858 16158 41860 16210
rect 41804 16146 41860 16158
rect 42140 16828 42364 16884
rect 42140 15986 42196 16828
rect 42364 16790 42420 16828
rect 42476 16100 42532 16110
rect 42588 16100 42644 16940
rect 42476 16098 42644 16100
rect 42476 16046 42478 16098
rect 42530 16046 42644 16098
rect 42476 16044 42644 16046
rect 42700 18228 42756 18238
rect 42476 16034 42532 16044
rect 42140 15934 42142 15986
rect 42194 15934 42196 15986
rect 42140 15922 42196 15934
rect 42364 15988 42420 15998
rect 42700 15988 42756 18172
rect 42812 16100 42868 19742
rect 42924 19124 42980 20300
rect 43260 20132 43316 20142
rect 43260 20038 43316 20076
rect 43708 19906 43764 19918
rect 43708 19854 43710 19906
rect 43762 19854 43764 19906
rect 43708 19796 43764 19854
rect 43708 19730 43764 19740
rect 43484 19234 43540 19246
rect 43484 19182 43486 19234
rect 43538 19182 43540 19234
rect 43036 19124 43092 19134
rect 42924 19122 43092 19124
rect 42924 19070 43038 19122
rect 43090 19070 43092 19122
rect 42924 19068 43092 19070
rect 42924 18338 42980 18350
rect 42924 18286 42926 18338
rect 42978 18286 42980 18338
rect 42924 17556 42980 18286
rect 43036 18340 43092 19068
rect 43484 18564 43540 19182
rect 43932 19234 43988 20524
rect 43932 19182 43934 19234
rect 43986 19182 43988 19234
rect 43932 19124 43988 19182
rect 43932 19058 43988 19068
rect 43036 18274 43092 18284
rect 43148 18562 43540 18564
rect 43148 18510 43486 18562
rect 43538 18510 43540 18562
rect 43148 18508 43540 18510
rect 42924 17490 42980 17500
rect 42812 16034 42868 16044
rect 42924 17220 42980 17230
rect 42924 16882 42980 17164
rect 43036 16996 43092 17006
rect 43148 16996 43204 18508
rect 43484 18498 43540 18508
rect 43596 18450 43652 18462
rect 43596 18398 43598 18450
rect 43650 18398 43652 18450
rect 43484 18340 43540 18350
rect 43596 18340 43652 18398
rect 43540 18284 43652 18340
rect 44044 18452 44100 18462
rect 43260 17668 43316 17678
rect 43484 17668 43540 18284
rect 43260 17666 43540 17668
rect 43260 17614 43262 17666
rect 43314 17614 43540 17666
rect 43260 17612 43540 17614
rect 43708 17666 43764 17678
rect 43708 17614 43710 17666
rect 43762 17614 43764 17666
rect 43260 17220 43316 17612
rect 43596 17556 43652 17566
rect 43260 17154 43316 17164
rect 43372 17444 43428 17454
rect 43372 16996 43428 17388
rect 43036 16994 43148 16996
rect 43036 16942 43038 16994
rect 43090 16942 43148 16994
rect 43036 16940 43148 16942
rect 43036 16930 43092 16940
rect 43148 16902 43204 16940
rect 43260 16940 43428 16996
rect 42924 16830 42926 16882
rect 42978 16830 42980 16882
rect 42028 15540 42084 15550
rect 42028 14642 42084 15484
rect 42028 14590 42030 14642
rect 42082 14590 42084 14642
rect 42028 14578 42084 14590
rect 41692 14354 41748 14364
rect 41916 14532 41972 14542
rect 41580 14242 41636 14252
rect 40908 12908 41188 12964
rect 41244 13972 41300 13982
rect 41244 13858 41300 13916
rect 41244 13806 41246 13858
rect 41298 13806 41300 13858
rect 40796 11508 40852 11518
rect 40796 11414 40852 11452
rect 40796 10948 40852 10958
rect 40796 7700 40852 10892
rect 40908 8260 40964 12908
rect 41244 12852 41300 13806
rect 41692 13860 41748 13870
rect 41692 13766 41748 13804
rect 41468 13524 41524 13534
rect 41468 12962 41524 13468
rect 41468 12910 41470 12962
rect 41522 12910 41524 12962
rect 41468 12898 41524 12910
rect 41692 13300 41748 13310
rect 41356 12852 41412 12862
rect 41244 12796 41356 12852
rect 41132 12740 41188 12750
rect 41132 12292 41188 12684
rect 41356 12404 41412 12796
rect 41468 12404 41524 12414
rect 41356 12402 41524 12404
rect 41356 12350 41470 12402
rect 41522 12350 41524 12402
rect 41356 12348 41524 12350
rect 41468 12338 41524 12348
rect 41692 12402 41748 13244
rect 41916 13074 41972 14476
rect 42364 13860 42420 15932
rect 42588 15932 42756 15988
rect 42588 15148 42644 15932
rect 42812 15874 42868 15886
rect 42812 15822 42814 15874
rect 42866 15822 42868 15874
rect 42812 15540 42868 15822
rect 42924 15764 42980 16830
rect 43036 16098 43092 16110
rect 43036 16046 43038 16098
rect 43090 16046 43092 16098
rect 43036 15876 43092 16046
rect 43036 15810 43092 15820
rect 42924 15698 42980 15708
rect 42812 15474 42868 15484
rect 42700 15428 42756 15438
rect 42700 15334 42756 15372
rect 43260 15148 43316 16940
rect 43596 16884 43652 17500
rect 43596 16790 43652 16828
rect 43484 16100 43540 16110
rect 43372 16044 43484 16100
rect 43372 15316 43428 16044
rect 43484 16006 43540 16044
rect 43484 15764 43540 15774
rect 43484 15538 43540 15708
rect 43484 15486 43486 15538
rect 43538 15486 43540 15538
rect 43484 15474 43540 15486
rect 43596 15540 43652 15550
rect 43708 15540 43764 17614
rect 44044 17444 44100 18396
rect 43932 17442 44100 17444
rect 43932 17390 44046 17442
rect 44098 17390 44100 17442
rect 43932 17388 44100 17390
rect 43596 15538 43708 15540
rect 43596 15486 43598 15538
rect 43650 15486 43708 15538
rect 43596 15484 43708 15486
rect 43596 15474 43652 15484
rect 43708 15474 43764 15484
rect 43820 16996 43876 17006
rect 43820 16098 43876 16940
rect 43932 16884 43988 17388
rect 44044 17378 44100 17388
rect 43932 16818 43988 16828
rect 44044 17220 44100 17230
rect 43820 16046 43822 16098
rect 43874 16046 43876 16098
rect 43372 15250 43428 15260
rect 43708 15316 43764 15326
rect 43820 15316 43876 16046
rect 43932 16548 43988 16558
rect 43932 16100 43988 16492
rect 43932 16034 43988 16044
rect 44044 15986 44100 17164
rect 44156 17108 44212 21310
rect 44268 21364 44324 22316
rect 44268 21298 44324 21308
rect 44492 21476 44548 21486
rect 44492 20242 44548 21420
rect 44492 20190 44494 20242
rect 44546 20190 44548 20242
rect 44492 20178 44548 20190
rect 44492 19572 44548 19582
rect 44268 18450 44324 18462
rect 44268 18398 44270 18450
rect 44322 18398 44324 18450
rect 44268 17556 44324 18398
rect 44268 17462 44324 17500
rect 44380 17444 44436 17454
rect 44380 17350 44436 17388
rect 44156 17052 44324 17108
rect 44156 16884 44212 16894
rect 44156 16790 44212 16828
rect 44044 15934 44046 15986
rect 44098 15934 44100 15986
rect 44044 15922 44100 15934
rect 44156 15874 44212 15886
rect 44156 15822 44158 15874
rect 44210 15822 44212 15874
rect 44156 15764 44212 15822
rect 44156 15698 44212 15708
rect 43708 15314 43876 15316
rect 43708 15262 43710 15314
rect 43762 15262 43876 15314
rect 43708 15260 43876 15262
rect 43932 15652 43988 15662
rect 43708 15250 43764 15260
rect 42364 13794 42420 13804
rect 42476 15092 42644 15148
rect 43148 15092 43316 15148
rect 41916 13022 41918 13074
rect 41970 13022 41972 13074
rect 41916 13010 41972 13022
rect 42140 13634 42196 13646
rect 42140 13582 42142 13634
rect 42194 13582 42196 13634
rect 42140 13412 42196 13582
rect 41692 12350 41694 12402
rect 41746 12350 41748 12402
rect 41692 12338 41748 12350
rect 41244 12292 41300 12302
rect 41020 12290 41300 12292
rect 41020 12238 41246 12290
rect 41298 12238 41300 12290
rect 41020 12236 41300 12238
rect 41020 8820 41076 12236
rect 41244 12226 41300 12236
rect 41804 12292 41860 12302
rect 42140 12292 42196 13356
rect 42252 13188 42308 13198
rect 42252 13074 42308 13132
rect 42252 13022 42254 13074
rect 42306 13022 42308 13074
rect 42252 13010 42308 13022
rect 42364 12964 42420 12974
rect 42364 12870 42420 12908
rect 42476 12628 42532 15092
rect 42588 14306 42644 14318
rect 42588 14254 42590 14306
rect 42642 14254 42644 14306
rect 42588 13972 42644 14254
rect 43036 13972 43092 13982
rect 42644 13916 42756 13972
rect 42588 13906 42644 13916
rect 42588 13746 42644 13758
rect 42588 13694 42590 13746
rect 42642 13694 42644 13746
rect 42588 13412 42644 13694
rect 42588 13346 42644 13356
rect 41860 12236 42196 12292
rect 42252 12572 42532 12628
rect 41804 12198 41860 12236
rect 41692 12068 41748 12078
rect 41692 11394 41748 12012
rect 41804 12068 41860 12078
rect 41804 12066 41972 12068
rect 41804 12014 41806 12066
rect 41858 12014 41972 12066
rect 41804 12012 41972 12014
rect 41804 12002 41860 12012
rect 41692 11342 41694 11394
rect 41746 11342 41748 11394
rect 41132 11284 41188 11294
rect 41132 10836 41188 11228
rect 41244 11170 41300 11182
rect 41244 11118 41246 11170
rect 41298 11118 41300 11170
rect 41244 10948 41300 11118
rect 41356 11172 41412 11182
rect 41692 11172 41748 11342
rect 41916 11396 41972 12012
rect 42140 11508 42196 11518
rect 42140 11414 42196 11452
rect 41916 11340 42084 11396
rect 41804 11284 41860 11294
rect 41804 11190 41860 11228
rect 41356 11078 41412 11116
rect 41468 11116 41748 11172
rect 41916 11170 41972 11182
rect 41916 11118 41918 11170
rect 41970 11118 41972 11170
rect 41356 10948 41412 10958
rect 41244 10892 41356 10948
rect 41356 10882 41412 10892
rect 41132 10780 41300 10836
rect 41132 10498 41188 10510
rect 41132 10446 41134 10498
rect 41186 10446 41188 10498
rect 41132 10386 41188 10446
rect 41132 10334 41134 10386
rect 41186 10334 41188 10386
rect 41132 10322 41188 10334
rect 41244 9938 41300 10780
rect 41468 10386 41524 11116
rect 41916 10948 41972 11118
rect 41692 10892 41972 10948
rect 41692 10834 41748 10892
rect 42028 10836 42084 11340
rect 42252 10836 42308 12572
rect 42364 12404 42420 12414
rect 42364 12310 42420 12348
rect 42476 12178 42532 12190
rect 42476 12126 42478 12178
rect 42530 12126 42532 12178
rect 41692 10782 41694 10834
rect 41746 10782 41748 10834
rect 41692 10770 41748 10782
rect 41916 10780 42084 10836
rect 42140 10780 42308 10836
rect 42364 11732 42420 11742
rect 42364 11506 42420 11676
rect 42364 11454 42366 11506
rect 42418 11454 42420 11506
rect 41916 10722 41972 10780
rect 41916 10670 41918 10722
rect 41970 10670 41972 10722
rect 41916 10658 41972 10670
rect 41468 10334 41470 10386
rect 41522 10334 41524 10386
rect 41468 10322 41524 10334
rect 41580 10388 41636 10398
rect 41580 10294 41636 10332
rect 41244 9886 41246 9938
rect 41298 9886 41300 9938
rect 41244 9874 41300 9886
rect 41692 9602 41748 9614
rect 41692 9550 41694 9602
rect 41746 9550 41748 9602
rect 41692 8932 41748 9550
rect 41692 8876 41972 8932
rect 41020 8764 41860 8820
rect 40908 8194 40964 8204
rect 41020 7700 41076 7710
rect 40796 7698 41076 7700
rect 40796 7646 41022 7698
rect 41074 7646 41076 7698
rect 40796 7644 41076 7646
rect 40796 7588 40852 7644
rect 41020 7634 41076 7644
rect 41468 7698 41524 7710
rect 41468 7646 41470 7698
rect 41522 7646 41524 7698
rect 40796 7522 40852 7532
rect 41468 7476 41524 7646
rect 41468 7028 41524 7420
rect 41468 6962 41524 6972
rect 41804 5236 41860 8764
rect 41916 8428 41972 8876
rect 41916 8372 42084 8428
rect 41916 7588 41972 7598
rect 41916 6802 41972 7532
rect 42028 7028 42084 8372
rect 42028 6962 42084 6972
rect 41916 6750 41918 6802
rect 41970 6750 41972 6802
rect 41916 6738 41972 6750
rect 39004 5070 39006 5122
rect 39058 5070 39060 5122
rect 39004 5058 39060 5070
rect 40236 5068 40740 5124
rect 41356 5234 41860 5236
rect 41356 5182 41806 5234
rect 41858 5182 41860 5234
rect 41356 5180 41860 5182
rect 39676 5010 39732 5022
rect 39676 4958 39678 5010
rect 39730 4958 39732 5010
rect 39676 4564 39732 4958
rect 39852 4732 40116 4742
rect 39908 4676 39956 4732
rect 40012 4676 40060 4732
rect 39852 4666 40116 4676
rect 40012 4564 40068 4574
rect 39676 4562 40068 4564
rect 39676 4510 40014 4562
rect 40066 4510 40068 4562
rect 39676 4508 40068 4510
rect 40012 4498 40068 4508
rect 38668 4386 38724 4396
rect 40236 4004 40292 5068
rect 40460 4788 40516 4798
rect 40348 4340 40404 4350
rect 40348 4246 40404 4284
rect 40236 3938 40292 3948
rect 38556 3714 38612 3724
rect 36876 3614 36878 3666
rect 36930 3614 36932 3666
rect 36876 3602 36932 3614
rect 36428 3390 36430 3442
rect 36482 3390 36484 3442
rect 36428 3378 36484 3390
rect 39340 3444 39396 3454
rect 40124 3444 40180 3454
rect 39340 3442 40180 3444
rect 39340 3390 39342 3442
rect 39394 3390 40126 3442
rect 40178 3390 40180 3442
rect 39340 3388 40180 3390
rect 40460 3442 40516 4732
rect 41020 4340 41076 4350
rect 41020 4246 41076 4284
rect 41356 4338 41412 5180
rect 41804 5170 41860 5180
rect 42140 5124 42196 10780
rect 42364 10724 42420 11454
rect 42476 11172 42532 12126
rect 42476 11106 42532 11116
rect 42588 10948 42644 10958
rect 42364 10668 42532 10724
rect 42252 10610 42308 10622
rect 42252 10558 42254 10610
rect 42306 10558 42308 10610
rect 42252 10388 42308 10558
rect 42364 10388 42420 10398
rect 42252 10332 42364 10388
rect 42364 10322 42420 10332
rect 42364 8148 42420 8158
rect 42364 7028 42420 8092
rect 42476 7252 42532 10668
rect 42588 9938 42644 10892
rect 42700 10834 42756 13916
rect 43036 13878 43092 13916
rect 42812 13746 42868 13758
rect 42812 13694 42814 13746
rect 42866 13694 42868 13746
rect 42812 13524 42868 13694
rect 42924 13748 42980 13758
rect 42924 13654 42980 13692
rect 42812 13458 42868 13468
rect 43148 12404 43204 15092
rect 43260 13860 43316 13870
rect 43260 13766 43316 13804
rect 43596 13858 43652 13870
rect 43596 13806 43598 13858
rect 43650 13806 43652 13858
rect 42924 12348 43204 12404
rect 43596 12402 43652 13806
rect 43820 13748 43876 13758
rect 43820 13654 43876 13692
rect 43932 13634 43988 15596
rect 44156 15540 44212 15550
rect 44156 15446 44212 15484
rect 44044 15316 44100 15326
rect 44268 15316 44324 17052
rect 44380 16772 44436 16782
rect 44380 16678 44436 16716
rect 44380 15876 44436 15886
rect 44380 15538 44436 15820
rect 44492 15652 44548 19516
rect 44492 15586 44548 15596
rect 44380 15486 44382 15538
rect 44434 15486 44436 15538
rect 44380 15474 44436 15486
rect 44268 15260 44436 15316
rect 44044 15222 44100 15260
rect 43932 13582 43934 13634
rect 43986 13582 43988 13634
rect 43932 13570 43988 13582
rect 44044 13746 44100 13758
rect 44044 13694 44046 13746
rect 44098 13694 44100 13746
rect 44044 12516 44100 13694
rect 44268 13300 44324 13310
rect 44268 13074 44324 13244
rect 44268 13022 44270 13074
rect 44322 13022 44324 13074
rect 44268 13010 44324 13022
rect 43596 12350 43598 12402
rect 43650 12350 43652 12402
rect 42812 12178 42868 12190
rect 42812 12126 42814 12178
rect 42866 12126 42868 12178
rect 42812 12068 42868 12126
rect 42812 12002 42868 12012
rect 42812 11172 42868 11182
rect 42812 11078 42868 11116
rect 42700 10782 42702 10834
rect 42754 10782 42756 10834
rect 42700 10770 42756 10782
rect 42924 10612 42980 12348
rect 43596 12338 43652 12350
rect 43708 12460 44100 12516
rect 44156 12964 44212 12974
rect 43036 12178 43092 12190
rect 43036 12126 43038 12178
rect 43090 12126 43092 12178
rect 43036 11956 43092 12126
rect 43484 12180 43540 12190
rect 43484 12086 43540 12124
rect 43036 11890 43092 11900
rect 43148 12066 43204 12078
rect 43148 12014 43150 12066
rect 43202 12014 43204 12066
rect 43148 11508 43204 12014
rect 43148 11442 43204 11452
rect 43596 11508 43652 11518
rect 43708 11508 43764 12460
rect 43932 12068 43988 12078
rect 43932 11974 43988 12012
rect 43596 11506 43764 11508
rect 43596 11454 43598 11506
rect 43650 11454 43764 11506
rect 43596 11452 43764 11454
rect 43596 11442 43652 11452
rect 43372 11396 43428 11406
rect 43260 11394 43428 11396
rect 43260 11342 43374 11394
rect 43426 11342 43428 11394
rect 43260 11340 43428 11342
rect 42588 9886 42590 9938
rect 42642 9886 42644 9938
rect 42588 9874 42644 9886
rect 42812 10556 42980 10612
rect 43148 10612 43204 10622
rect 43260 10612 43316 11340
rect 43372 11330 43428 11340
rect 43484 11396 43540 11406
rect 43484 10724 43540 11340
rect 43820 11396 43876 11406
rect 44044 11396 44100 11406
rect 44156 11396 44212 12908
rect 43876 11340 43988 11396
rect 43820 11302 43876 11340
rect 43596 11170 43652 11182
rect 43596 11118 43598 11170
rect 43650 11118 43652 11170
rect 43596 10836 43652 11118
rect 43596 10780 43764 10836
rect 43484 10668 43652 10724
rect 43204 10556 43316 10612
rect 43372 10610 43428 10622
rect 43372 10558 43374 10610
rect 43426 10558 43428 10610
rect 42812 9156 42868 10556
rect 43036 10052 43092 10062
rect 43036 9492 43092 9996
rect 43148 9938 43204 10556
rect 43148 9886 43150 9938
rect 43202 9886 43204 9938
rect 43148 9874 43204 9886
rect 43260 10052 43316 10062
rect 43036 9426 43092 9436
rect 42812 9090 42868 9100
rect 43260 8930 43316 9996
rect 43260 8878 43262 8930
rect 43314 8878 43316 8930
rect 43260 8866 43316 8878
rect 42588 8372 42644 8382
rect 42588 7588 42644 8316
rect 42588 7494 42644 7532
rect 42476 7186 42532 7196
rect 42924 7252 42980 7262
rect 43260 7252 43316 7262
rect 42924 7250 43204 7252
rect 42924 7198 42926 7250
rect 42978 7198 43204 7250
rect 42924 7196 43204 7198
rect 42924 7186 42980 7196
rect 42924 7028 42980 7038
rect 42364 6972 42532 7028
rect 42028 5068 42196 5124
rect 42364 6018 42420 6030
rect 42364 5966 42366 6018
rect 42418 5966 42420 6018
rect 42028 4788 42084 5068
rect 42364 5012 42420 5966
rect 41356 4286 41358 4338
rect 41410 4286 41412 4338
rect 41356 4274 41412 4286
rect 41916 4732 42084 4788
rect 42140 4956 42364 5012
rect 41916 4116 41972 4732
rect 42140 4450 42196 4956
rect 42364 4946 42420 4956
rect 42140 4398 42142 4450
rect 42194 4398 42196 4450
rect 42140 4386 42196 4398
rect 42028 4340 42084 4350
rect 42028 4246 42084 4284
rect 41916 4050 41972 4060
rect 42476 3780 42532 6972
rect 42924 6692 42980 6972
rect 42700 6690 42980 6692
rect 42700 6638 42926 6690
rect 42978 6638 42980 6690
rect 42700 6636 42980 6638
rect 43148 6692 43204 7196
rect 43260 7158 43316 7196
rect 43372 6916 43428 10558
rect 43596 10610 43652 10668
rect 43596 10558 43598 10610
rect 43650 10558 43652 10610
rect 43596 10546 43652 10558
rect 43484 10498 43540 10510
rect 43484 10446 43486 10498
rect 43538 10446 43540 10498
rect 43484 10388 43540 10446
rect 43708 10388 43764 10780
rect 43820 10612 43876 10622
rect 43820 10518 43876 10556
rect 43484 10322 43540 10332
rect 43596 10332 43764 10388
rect 43596 9828 43652 10332
rect 43932 10276 43988 11340
rect 44044 11394 44212 11396
rect 44044 11342 44046 11394
rect 44098 11342 44212 11394
rect 44044 11340 44212 11342
rect 44044 11330 44100 11340
rect 44268 10500 44324 10510
rect 44268 10406 44324 10444
rect 43484 9772 43652 9828
rect 43708 10220 43988 10276
rect 43484 9044 43540 9772
rect 43708 9716 43764 10220
rect 43596 9660 43764 9716
rect 43596 9602 43652 9660
rect 43596 9550 43598 9602
rect 43650 9550 43652 9602
rect 43596 9538 43652 9550
rect 43484 8978 43540 8988
rect 44380 8596 44436 15260
rect 44604 15148 44660 22652
rect 44940 22484 44996 22494
rect 44716 22482 44996 22484
rect 44716 22430 44942 22482
rect 44994 22430 44996 22482
rect 44716 22428 44996 22430
rect 44716 21586 44772 22428
rect 44940 22418 44996 22428
rect 45052 22370 45108 22652
rect 45164 22642 45220 22652
rect 45052 22318 45054 22370
rect 45106 22318 45108 22370
rect 45052 22306 45108 22318
rect 45276 22370 45332 24668
rect 45388 24612 45444 24622
rect 45388 24050 45444 24556
rect 45836 24612 45892 24782
rect 45836 24546 45892 24556
rect 45948 24052 46004 25228
rect 46172 24724 46228 26236
rect 46284 26068 46340 26078
rect 46396 26068 46452 26078
rect 46340 26066 46452 26068
rect 46340 26014 46398 26066
rect 46450 26014 46452 26066
rect 46340 26012 46452 26014
rect 46284 24724 46340 26012
rect 46396 26002 46452 26012
rect 46396 25620 46452 25630
rect 46844 25620 46900 27020
rect 46396 25618 46900 25620
rect 46396 25566 46398 25618
rect 46450 25566 46900 25618
rect 46396 25564 46900 25566
rect 46396 25554 46452 25564
rect 46844 25506 46900 25564
rect 46844 25454 46846 25506
rect 46898 25454 46900 25506
rect 46844 25442 46900 25454
rect 46620 24948 46676 24986
rect 46620 24882 46676 24892
rect 46620 24724 46676 24734
rect 46284 24722 46676 24724
rect 46284 24670 46622 24722
rect 46674 24670 46676 24722
rect 46284 24668 46676 24670
rect 46172 24630 46228 24668
rect 46620 24658 46676 24668
rect 46956 24724 47012 27580
rect 47068 26908 47124 30380
rect 48076 30212 48132 30222
rect 48076 30118 48132 30156
rect 47404 30098 47460 30110
rect 47404 30046 47406 30098
rect 47458 30046 47460 30098
rect 47180 29986 47236 29998
rect 47180 29934 47182 29986
rect 47234 29934 47236 29986
rect 47180 29540 47236 29934
rect 47180 29474 47236 29484
rect 47292 28756 47348 28766
rect 47292 28642 47348 28700
rect 47292 28590 47294 28642
rect 47346 28590 47348 28642
rect 47292 28578 47348 28590
rect 47404 27972 47460 30046
rect 47740 29988 47796 29998
rect 47796 29932 48244 29988
rect 47740 29894 47796 29932
rect 47740 29650 47796 29662
rect 47740 29598 47742 29650
rect 47794 29598 47796 29650
rect 47740 29540 47796 29598
rect 47740 29474 47796 29484
rect 47852 29538 47908 29550
rect 47852 29486 47854 29538
rect 47906 29486 47908 29538
rect 47852 29428 47908 29486
rect 47852 29362 47908 29372
rect 47852 28644 47908 28654
rect 47852 28550 47908 28588
rect 48188 28530 48244 29932
rect 48412 29652 48468 29662
rect 48300 29540 48356 29550
rect 48300 28866 48356 29484
rect 48300 28814 48302 28866
rect 48354 28814 48356 28866
rect 48300 28802 48356 28814
rect 48188 28478 48190 28530
rect 48242 28478 48244 28530
rect 48188 28466 48244 28478
rect 48300 28532 48356 28542
rect 48412 28532 48468 29596
rect 48300 28530 48468 28532
rect 48300 28478 48302 28530
rect 48354 28478 48468 28530
rect 48300 28476 48468 28478
rect 48524 28532 48580 31948
rect 48636 31556 48692 31566
rect 48636 31462 48692 31500
rect 48748 30212 48804 33966
rect 49196 34020 49252 34030
rect 49308 34020 49364 35420
rect 49532 35410 49588 35420
rect 49512 35308 49776 35318
rect 49568 35252 49616 35308
rect 49672 35252 49720 35308
rect 49512 35242 49776 35252
rect 49420 34468 49476 34478
rect 49420 34130 49476 34412
rect 49420 34078 49422 34130
rect 49474 34078 49476 34130
rect 49420 34066 49476 34078
rect 49868 34132 49924 36430
rect 50428 36260 50484 36270
rect 50484 36204 50596 36260
rect 50428 36166 50484 36204
rect 50428 35700 50484 35710
rect 50428 35606 50484 35644
rect 49868 34066 49924 34076
rect 49980 34802 50036 34814
rect 49980 34750 49982 34802
rect 50034 34750 50036 34802
rect 49196 34018 49364 34020
rect 49196 33966 49198 34018
rect 49250 33966 49364 34018
rect 49196 33964 49364 33966
rect 48860 33572 48916 33582
rect 48860 33478 48916 33516
rect 49196 33348 49252 33964
rect 49512 33740 49776 33750
rect 49568 33684 49616 33740
rect 49672 33684 49720 33740
rect 49512 33674 49776 33684
rect 49196 33254 49252 33292
rect 48972 33122 49028 33134
rect 48972 33070 48974 33122
rect 49026 33070 49028 33122
rect 48972 31892 49028 33070
rect 49868 33124 49924 33134
rect 49868 32786 49924 33068
rect 49868 32734 49870 32786
rect 49922 32734 49924 32786
rect 49868 32722 49924 32734
rect 49512 32172 49776 32182
rect 49568 32116 49616 32172
rect 49672 32116 49720 32172
rect 49512 32106 49776 32116
rect 48972 31826 49028 31836
rect 49644 31668 49700 31678
rect 49868 31668 49924 31678
rect 49644 31574 49700 31612
rect 49756 31666 49924 31668
rect 49756 31614 49870 31666
rect 49922 31614 49924 31666
rect 49756 31612 49924 31614
rect 48972 31556 49028 31566
rect 48972 31462 49028 31500
rect 49420 31556 49476 31566
rect 49420 31218 49476 31500
rect 49420 31166 49422 31218
rect 49474 31166 49476 31218
rect 49420 31154 49476 31166
rect 49644 31220 49700 31230
rect 49756 31220 49812 31612
rect 49868 31602 49924 31612
rect 49980 31554 50036 34750
rect 50540 33236 50596 36204
rect 50652 35810 50708 35822
rect 50652 35758 50654 35810
rect 50706 35758 50708 35810
rect 50652 35252 50708 35758
rect 50652 34692 50708 35196
rect 50652 34626 50708 34636
rect 50876 34020 50932 39200
rect 52556 37156 52612 37166
rect 52444 36708 52500 36718
rect 52332 36484 52388 36494
rect 52108 36372 52164 36382
rect 52108 36370 52276 36372
rect 52108 36318 52110 36370
rect 52162 36318 52276 36370
rect 52108 36316 52276 36318
rect 52108 36306 52164 36316
rect 50988 35700 51044 35710
rect 50988 35606 51044 35644
rect 51324 35698 51380 35710
rect 51324 35646 51326 35698
rect 51378 35646 51380 35698
rect 51324 35252 51380 35646
rect 52108 35588 52164 35598
rect 51324 35186 51380 35196
rect 51884 35586 52164 35588
rect 51884 35534 52110 35586
rect 52162 35534 52164 35586
rect 51884 35532 52164 35534
rect 51548 35028 51604 35038
rect 51324 34020 51380 34030
rect 50876 34018 51380 34020
rect 50876 33966 51326 34018
rect 51378 33966 51380 34018
rect 50876 33964 51380 33966
rect 51324 33954 51380 33964
rect 50540 33170 50596 33180
rect 50652 33124 50708 33134
rect 50652 32562 50708 33068
rect 50652 32510 50654 32562
rect 50706 32510 50708 32562
rect 50428 32452 50484 32462
rect 50428 32450 50596 32452
rect 50428 32398 50430 32450
rect 50482 32398 50596 32450
rect 50428 32396 50596 32398
rect 50428 32386 50484 32396
rect 49980 31502 49982 31554
rect 50034 31502 50036 31554
rect 49980 31490 50036 31502
rect 50092 31892 50148 31902
rect 49644 31218 49812 31220
rect 49644 31166 49646 31218
rect 49698 31166 49812 31218
rect 49644 31164 49812 31166
rect 49644 31154 49700 31164
rect 48972 31108 49028 31118
rect 48748 30146 48804 30156
rect 48860 31052 48972 31108
rect 48636 29428 48692 29438
rect 48636 28644 48692 29372
rect 48860 29092 48916 31052
rect 48972 31014 49028 31052
rect 49308 31108 49364 31118
rect 49308 31014 49364 31052
rect 49512 30604 49776 30614
rect 49568 30548 49616 30604
rect 49672 30548 49720 30604
rect 49512 30538 49776 30548
rect 48972 30212 49028 30222
rect 48972 29428 49028 30156
rect 49196 29708 49700 29764
rect 49084 29652 49140 29662
rect 49084 29558 49140 29596
rect 49196 29650 49252 29708
rect 49196 29598 49198 29650
rect 49250 29598 49252 29650
rect 49196 29586 49252 29598
rect 49644 29538 49700 29708
rect 49868 29652 49924 29662
rect 49644 29486 49646 29538
rect 49698 29486 49700 29538
rect 49644 29474 49700 29486
rect 49756 29540 49812 29550
rect 49756 29446 49812 29484
rect 49308 29428 49364 29438
rect 48972 29426 49364 29428
rect 48972 29374 49310 29426
rect 49362 29374 49364 29426
rect 48972 29372 49364 29374
rect 49308 29362 49364 29372
rect 49756 29204 49812 29242
rect 49756 29138 49812 29148
rect 48860 29036 49140 29092
rect 48860 28756 48916 28766
rect 48636 28588 48804 28644
rect 47404 27906 47460 27916
rect 48076 27972 48132 27982
rect 48300 27972 48356 28476
rect 48524 28466 48580 28476
rect 48076 27970 48356 27972
rect 48076 27918 48078 27970
rect 48130 27918 48356 27970
rect 48076 27916 48356 27918
rect 48076 27906 48132 27916
rect 47740 27858 47796 27870
rect 47740 27806 47742 27858
rect 47794 27806 47796 27858
rect 47292 27634 47348 27646
rect 47292 27582 47294 27634
rect 47346 27582 47348 27634
rect 47068 26852 47236 26908
rect 46956 24658 47012 24668
rect 45388 23998 45390 24050
rect 45442 23998 45444 24050
rect 45388 23986 45444 23998
rect 45612 24050 46004 24052
rect 45612 23998 45950 24050
rect 46002 23998 46004 24050
rect 45612 23996 46004 23998
rect 45612 23492 45668 23996
rect 45948 23986 46004 23996
rect 45276 22318 45278 22370
rect 45330 22318 45332 22370
rect 45276 22306 45332 22318
rect 45388 23380 45444 23390
rect 44940 22148 44996 22158
rect 45388 22148 45444 23324
rect 45500 23044 45556 23054
rect 45500 22950 45556 22988
rect 45500 22372 45556 22382
rect 45612 22372 45668 23436
rect 46172 23380 46228 23390
rect 46172 23286 46228 23324
rect 47180 23378 47236 26852
rect 47292 26852 47348 27582
rect 47740 26908 47796 27806
rect 47740 26852 47908 26908
rect 47292 26786 47348 26796
rect 47852 26740 47908 26852
rect 47852 26674 47908 26684
rect 48412 26852 48468 26862
rect 47292 26628 47348 26638
rect 47292 25618 47348 26572
rect 48188 26180 48244 26190
rect 47292 25566 47294 25618
rect 47346 25566 47348 25618
rect 47292 25554 47348 25566
rect 47516 25732 47572 25742
rect 47516 24946 47572 25676
rect 47852 25732 47908 25742
rect 48188 25732 48244 26124
rect 48412 26068 48468 26796
rect 48412 26002 48468 26012
rect 47908 25676 48244 25732
rect 47516 24894 47518 24946
rect 47570 24894 47572 24946
rect 47516 24882 47572 24894
rect 47740 25394 47796 25406
rect 47740 25342 47742 25394
rect 47794 25342 47796 25394
rect 47740 25284 47796 25342
rect 47852 25394 47908 25676
rect 48748 25618 48804 28588
rect 48860 28082 48916 28700
rect 48860 28030 48862 28082
rect 48914 28030 48916 28082
rect 48860 28018 48916 28030
rect 48972 28532 49028 28542
rect 48972 26402 49028 28476
rect 49084 26516 49140 29036
rect 49512 29036 49776 29046
rect 49568 28980 49616 29036
rect 49672 28980 49720 29036
rect 49512 28970 49776 28980
rect 49756 28084 49812 28094
rect 49756 27990 49812 28028
rect 49196 27970 49252 27982
rect 49196 27918 49198 27970
rect 49250 27918 49252 27970
rect 49196 26852 49252 27918
rect 49512 27468 49776 27478
rect 49568 27412 49616 27468
rect 49672 27412 49720 27468
rect 49512 27402 49776 27412
rect 49868 27300 49924 29596
rect 49980 28756 50036 28766
rect 49980 28662 50036 28700
rect 49980 28084 50036 28094
rect 49980 27990 50036 28028
rect 49196 26786 49252 26796
rect 49756 27244 49924 27300
rect 49532 26740 49588 26750
rect 49084 26460 49252 26516
rect 48972 26350 48974 26402
rect 49026 26350 49028 26402
rect 48972 26338 49028 26350
rect 49084 26290 49140 26302
rect 49084 26238 49086 26290
rect 49138 26238 49140 26290
rect 49084 26180 49140 26238
rect 49084 26114 49140 26124
rect 48748 25566 48750 25618
rect 48802 25566 48804 25618
rect 48748 25554 48804 25566
rect 48076 25508 48132 25518
rect 48300 25508 48356 25518
rect 48076 25506 48356 25508
rect 48076 25454 48078 25506
rect 48130 25454 48302 25506
rect 48354 25454 48356 25506
rect 48076 25452 48356 25454
rect 48076 25442 48132 25452
rect 48300 25442 48356 25452
rect 47852 25342 47854 25394
rect 47906 25342 47908 25394
rect 47852 25330 47908 25342
rect 48636 25394 48692 25406
rect 48636 25342 48638 25394
rect 48690 25342 48692 25394
rect 47740 23940 47796 25228
rect 48636 24948 48692 25342
rect 47852 23940 47908 23950
rect 47740 23938 47908 23940
rect 47740 23886 47854 23938
rect 47906 23886 47908 23938
rect 47740 23884 47908 23886
rect 48636 23940 48692 24892
rect 48748 23940 48804 23950
rect 48636 23938 48804 23940
rect 48636 23886 48750 23938
rect 48802 23886 48804 23938
rect 48636 23884 48804 23886
rect 47516 23826 47572 23838
rect 47516 23774 47518 23826
rect 47570 23774 47572 23826
rect 47516 23604 47572 23774
rect 47516 23538 47572 23548
rect 47180 23326 47182 23378
rect 47234 23326 47236 23378
rect 47180 23268 47236 23326
rect 47516 23380 47572 23390
rect 47516 23286 47572 23324
rect 47180 23202 47236 23212
rect 45948 23154 46004 23166
rect 45948 23102 45950 23154
rect 46002 23102 46004 23154
rect 45948 23044 46004 23102
rect 45948 22978 46004 22988
rect 46732 23042 46788 23054
rect 46732 22990 46734 23042
rect 46786 22990 46788 23042
rect 45500 22370 45668 22372
rect 45500 22318 45502 22370
rect 45554 22318 45668 22370
rect 45500 22316 45668 22318
rect 46172 22708 46228 22718
rect 46172 22372 46228 22652
rect 46620 22484 46676 22494
rect 46620 22390 46676 22428
rect 46172 22370 46564 22372
rect 46172 22318 46174 22370
rect 46226 22318 46564 22370
rect 46172 22316 46564 22318
rect 45500 22306 45556 22316
rect 46172 22306 46228 22316
rect 44716 21534 44718 21586
rect 44770 21534 44772 21586
rect 44716 21522 44772 21534
rect 44828 21588 44884 21598
rect 44828 20130 44884 21532
rect 44940 21140 44996 22092
rect 45276 22092 45444 22148
rect 44940 20802 44996 21084
rect 45164 21586 45220 21598
rect 45164 21534 45166 21586
rect 45218 21534 45220 21586
rect 45164 20914 45220 21534
rect 45164 20862 45166 20914
rect 45218 20862 45220 20914
rect 45164 20850 45220 20862
rect 44940 20750 44942 20802
rect 44994 20750 44996 20802
rect 44940 20738 44996 20750
rect 45276 20802 45332 22092
rect 46508 21812 46564 22316
rect 46732 22148 46788 22990
rect 47068 22820 47124 22830
rect 47068 22372 47124 22764
rect 46732 22082 46788 22092
rect 46844 22370 47124 22372
rect 46844 22318 47070 22370
rect 47122 22318 47124 22370
rect 46844 22316 47124 22318
rect 46620 21812 46676 21822
rect 46508 21810 46676 21812
rect 46508 21758 46622 21810
rect 46674 21758 46676 21810
rect 46508 21756 46676 21758
rect 45612 21588 45668 21598
rect 45612 21494 45668 21532
rect 45500 21476 45556 21486
rect 45500 21382 45556 21420
rect 45276 20750 45278 20802
rect 45330 20750 45332 20802
rect 45276 20738 45332 20750
rect 45388 21364 45444 21374
rect 45388 20802 45444 21308
rect 45948 21364 46004 21374
rect 45948 21270 46004 21308
rect 45500 21140 45556 21150
rect 45556 21084 45892 21140
rect 45500 21074 45556 21084
rect 45388 20750 45390 20802
rect 45442 20750 45444 20802
rect 45052 20580 45108 20590
rect 45164 20580 45220 20590
rect 45052 20578 45164 20580
rect 45052 20526 45054 20578
rect 45106 20526 45164 20578
rect 45052 20524 45164 20526
rect 45052 20514 45108 20524
rect 44828 20078 44830 20130
rect 44882 20078 44884 20130
rect 44828 20066 44884 20078
rect 44940 19124 44996 19134
rect 44940 19030 44996 19068
rect 44716 18452 44772 18462
rect 44716 18358 44772 18396
rect 45052 18226 45108 18238
rect 45052 18174 45054 18226
rect 45106 18174 45108 18226
rect 45052 17668 45108 18174
rect 45052 17602 45108 17612
rect 45164 17444 45220 20524
rect 45388 20244 45444 20750
rect 45276 20188 45444 20244
rect 45276 20130 45332 20188
rect 45276 20078 45278 20130
rect 45330 20078 45332 20130
rect 45276 20066 45332 20078
rect 45836 20130 45892 21084
rect 46620 21026 46676 21756
rect 46620 20974 46622 21026
rect 46674 20974 46676 21026
rect 46620 20962 46676 20974
rect 46844 20914 46900 22316
rect 47068 22306 47124 22316
rect 47180 22148 47236 22158
rect 46844 20862 46846 20914
rect 46898 20862 46900 20914
rect 46844 20850 46900 20862
rect 47068 22146 47236 22148
rect 47068 22094 47182 22146
rect 47234 22094 47236 22146
rect 47068 22092 47236 22094
rect 45948 20580 46004 20590
rect 45948 20486 46004 20524
rect 45836 20078 45838 20130
rect 45890 20078 45892 20130
rect 45836 20066 45892 20078
rect 47068 19908 47124 22092
rect 47180 22082 47236 22092
rect 47852 21812 47908 23884
rect 48748 23874 48804 23884
rect 47964 23268 48020 23278
rect 48020 23212 48132 23268
rect 47964 23202 48020 23212
rect 47964 21812 48020 21822
rect 47852 21810 48020 21812
rect 47852 21758 47966 21810
rect 48018 21758 48020 21810
rect 47852 21756 48020 21758
rect 47964 21746 48020 21756
rect 47516 21588 47572 21598
rect 47404 21532 47516 21588
rect 47180 21476 47236 21486
rect 47180 21382 47236 21420
rect 47180 21026 47236 21038
rect 47180 20974 47182 21026
rect 47234 20974 47236 21026
rect 47180 20914 47236 20974
rect 47180 20862 47182 20914
rect 47234 20862 47236 20914
rect 47180 20850 47236 20862
rect 47068 19842 47124 19852
rect 46732 19460 46788 19470
rect 46620 19404 46732 19460
rect 45052 17388 45220 17444
rect 45388 18450 45444 18462
rect 45388 18398 45390 18450
rect 45442 18398 45444 18450
rect 44940 16882 44996 16894
rect 44940 16830 44942 16882
rect 44994 16830 44996 16882
rect 44828 16772 44884 16782
rect 44940 16772 44996 16830
rect 44884 16716 44996 16772
rect 44828 16098 44884 16716
rect 44828 16046 44830 16098
rect 44882 16046 44884 16098
rect 44828 16034 44884 16046
rect 44716 15876 44772 15886
rect 44716 15314 44772 15820
rect 44716 15262 44718 15314
rect 44770 15262 44772 15314
rect 44716 15250 44772 15262
rect 44604 15092 44772 15148
rect 44604 13412 44660 13422
rect 44492 12292 44548 12302
rect 44492 12178 44548 12236
rect 44492 12126 44494 12178
rect 44546 12126 44548 12178
rect 44492 12114 44548 12126
rect 44604 11844 44660 13356
rect 44604 11060 44660 11788
rect 44604 10994 44660 11004
rect 44380 8540 44660 8596
rect 44044 8260 44100 8270
rect 43932 7812 43988 7822
rect 43932 7586 43988 7756
rect 43932 7534 43934 7586
rect 43986 7534 43988 7586
rect 43932 7028 43988 7534
rect 44044 7588 44100 8204
rect 44604 7812 44660 8540
rect 44604 7698 44660 7756
rect 44604 7646 44606 7698
rect 44658 7646 44660 7698
rect 44604 7634 44660 7646
rect 44044 7474 44100 7532
rect 44044 7422 44046 7474
rect 44098 7422 44100 7474
rect 44044 7410 44100 7422
rect 43932 6962 43988 6972
rect 43372 6850 43428 6860
rect 43260 6692 43316 6702
rect 43148 6690 43316 6692
rect 43148 6638 43262 6690
rect 43314 6638 43316 6690
rect 43148 6636 43316 6638
rect 42700 6130 42756 6636
rect 42924 6626 42980 6636
rect 43260 6626 43316 6636
rect 43932 6692 43988 6702
rect 43596 6468 43652 6478
rect 43596 6466 43876 6468
rect 43596 6414 43598 6466
rect 43650 6414 43876 6466
rect 43596 6412 43876 6414
rect 43596 6402 43652 6412
rect 42700 6078 42702 6130
rect 42754 6078 42756 6130
rect 42700 6066 42756 6078
rect 42812 6244 42868 6254
rect 42700 5124 42756 5134
rect 42700 5030 42756 5068
rect 42812 4562 42868 6188
rect 43820 6018 43876 6412
rect 43820 5966 43822 6018
rect 43874 5966 43876 6018
rect 43820 5954 43876 5966
rect 43036 5908 43092 5918
rect 43092 5852 43316 5908
rect 43036 5814 43092 5852
rect 43260 5124 43316 5852
rect 43932 5124 43988 6636
rect 43260 5068 43540 5124
rect 43260 5010 43316 5068
rect 43260 4958 43262 5010
rect 43314 4958 43316 5010
rect 43260 4946 43316 4958
rect 42924 4900 42980 4910
rect 42924 4806 42980 4844
rect 43484 4788 43540 5068
rect 43596 5068 43988 5124
rect 43596 5010 43652 5068
rect 43596 4958 43598 5010
rect 43650 4958 43652 5010
rect 43596 4946 43652 4958
rect 43932 5010 43988 5068
rect 44268 6356 44324 6366
rect 44268 5122 44324 6300
rect 44268 5070 44270 5122
rect 44322 5070 44324 5122
rect 44268 5058 44324 5070
rect 43932 4958 43934 5010
rect 43986 4958 43988 5010
rect 43932 4946 43988 4958
rect 44380 4900 44436 4910
rect 43484 4732 43764 4788
rect 42812 4510 42814 4562
rect 42866 4510 42868 4562
rect 42812 4340 42868 4510
rect 42812 4274 42868 4284
rect 43708 4338 43764 4732
rect 44380 4450 44436 4844
rect 44380 4398 44382 4450
rect 44434 4398 44436 4450
rect 44380 4386 44436 4398
rect 43708 4286 43710 4338
rect 43762 4286 43764 4338
rect 43708 4274 43764 4286
rect 42476 3714 42532 3724
rect 44716 3556 44772 15092
rect 44828 13300 44884 13310
rect 44828 5348 44884 13244
rect 44940 13188 44996 13198
rect 44940 13074 44996 13132
rect 44940 13022 44942 13074
rect 44994 13022 44996 13074
rect 44940 13010 44996 13022
rect 44940 11396 44996 11406
rect 44940 11302 44996 11340
rect 44940 9602 44996 9614
rect 44940 9550 44942 9602
rect 44994 9550 44996 9602
rect 44940 8258 44996 9550
rect 44940 8206 44942 8258
rect 44994 8206 44996 8258
rect 44940 8194 44996 8206
rect 44828 5282 44884 5292
rect 44940 5124 44996 5134
rect 44940 5030 44996 5068
rect 45052 4788 45108 17388
rect 45164 15202 45220 15214
rect 45164 15150 45166 15202
rect 45218 15150 45220 15202
rect 45164 15148 45220 15150
rect 45388 15148 45444 18398
rect 46060 18340 46116 18350
rect 46060 18338 46228 18340
rect 46060 18286 46062 18338
rect 46114 18286 46228 18338
rect 46060 18284 46228 18286
rect 46060 18274 46116 18284
rect 45500 17778 45556 17790
rect 45500 17726 45502 17778
rect 45554 17726 45556 17778
rect 45500 17108 45556 17726
rect 45500 17042 45556 17052
rect 46060 17220 46116 17230
rect 46060 16994 46116 17164
rect 46172 17108 46228 18284
rect 46396 17668 46452 17678
rect 46396 17574 46452 17612
rect 46620 17444 46676 19404
rect 46732 19394 46788 19404
rect 47068 19234 47124 19246
rect 47068 19182 47070 19234
rect 47122 19182 47124 19234
rect 47068 17668 47124 19182
rect 47404 17780 47460 21532
rect 47516 21494 47572 21532
rect 47740 21586 47796 21598
rect 47740 21534 47742 21586
rect 47794 21534 47796 21586
rect 47628 20580 47684 20590
rect 47740 20580 47796 21534
rect 48076 21586 48132 23212
rect 49196 22596 49252 26460
rect 49308 26180 49364 26190
rect 49308 24948 49364 26124
rect 49532 26178 49588 26684
rect 49532 26126 49534 26178
rect 49586 26126 49588 26178
rect 49532 26114 49588 26126
rect 49756 26068 49812 27244
rect 50092 27076 50148 31836
rect 50204 31668 50260 31678
rect 50540 31668 50596 32396
rect 50652 32004 50708 32510
rect 50652 31938 50708 31948
rect 50764 32674 50820 32686
rect 50764 32622 50766 32674
rect 50818 32622 50820 32674
rect 50652 31668 50708 31678
rect 50204 31666 50372 31668
rect 50204 31614 50206 31666
rect 50258 31614 50372 31666
rect 50204 31612 50372 31614
rect 50204 31602 50260 31612
rect 50316 28980 50372 31612
rect 50540 31666 50708 31668
rect 50540 31614 50654 31666
rect 50706 31614 50708 31666
rect 50540 31612 50708 31614
rect 50540 31332 50596 31612
rect 50652 31602 50708 31612
rect 50764 31668 50820 32622
rect 50988 32564 51044 32574
rect 50988 32562 51492 32564
rect 50988 32510 50990 32562
rect 51042 32510 51492 32562
rect 50988 32508 51492 32510
rect 50988 32498 51044 32508
rect 51212 32004 51268 32014
rect 51436 32004 51492 32508
rect 51548 32562 51604 34972
rect 51772 34580 51828 34590
rect 51660 33348 51716 33358
rect 51660 33254 51716 33292
rect 51772 33234 51828 34524
rect 51772 33182 51774 33234
rect 51826 33182 51828 33234
rect 51772 33170 51828 33182
rect 51548 32510 51550 32562
rect 51602 32510 51604 32562
rect 51548 32498 51604 32510
rect 51436 31948 51716 32004
rect 50764 31666 50932 31668
rect 50764 31614 50766 31666
rect 50818 31614 50932 31666
rect 50764 31612 50932 31614
rect 50764 31602 50820 31612
rect 50428 29652 50484 29662
rect 50540 29652 50596 31276
rect 50876 31556 50932 31612
rect 50876 31220 50932 31500
rect 50988 31554 51044 31566
rect 50988 31502 50990 31554
rect 51042 31502 51044 31554
rect 50988 31444 51044 31502
rect 50988 31378 51044 31388
rect 51100 31220 51156 31230
rect 50876 31218 51156 31220
rect 50876 31166 51102 31218
rect 51154 31166 51156 31218
rect 50876 31164 51156 31166
rect 51100 31154 51156 31164
rect 50988 30994 51044 31006
rect 50988 30942 50990 30994
rect 51042 30942 51044 30994
rect 50652 30884 50708 30894
rect 50988 30884 51044 30942
rect 50652 30882 51044 30884
rect 50652 30830 50654 30882
rect 50706 30830 51044 30882
rect 50652 30828 51044 30830
rect 50652 30818 50708 30828
rect 50484 29596 50596 29652
rect 50988 29652 51044 30828
rect 51212 30772 51268 31948
rect 51660 31778 51716 31948
rect 51660 31726 51662 31778
rect 51714 31726 51716 31778
rect 51660 31714 51716 31726
rect 51436 31668 51492 31678
rect 51324 30996 51380 31006
rect 51436 30996 51492 31612
rect 51884 31554 51940 35532
rect 52108 35522 52164 35532
rect 52220 35140 52276 36316
rect 52220 35074 52276 35084
rect 52332 35812 52388 36428
rect 52108 35026 52164 35038
rect 52108 34974 52110 35026
rect 52162 34974 52164 35026
rect 52108 34916 52164 34974
rect 52332 34916 52388 35756
rect 52108 34860 52388 34916
rect 51996 34020 52052 34030
rect 51996 33346 52052 33964
rect 51996 33294 51998 33346
rect 52050 33294 52052 33346
rect 51996 33282 52052 33294
rect 52332 32452 52388 32462
rect 52108 32450 52388 32452
rect 52108 32398 52334 32450
rect 52386 32398 52388 32450
rect 52108 32396 52388 32398
rect 51884 31502 51886 31554
rect 51938 31502 51940 31554
rect 51884 31490 51940 31502
rect 51996 31666 52052 31678
rect 51996 31614 51998 31666
rect 52050 31614 52052 31666
rect 51548 31444 51604 31454
rect 51604 31388 51828 31444
rect 51548 31378 51604 31388
rect 51772 31106 51828 31388
rect 51996 31332 52052 31614
rect 51772 31054 51774 31106
rect 51826 31054 51828 31106
rect 51772 31042 51828 31054
rect 51884 31276 52052 31332
rect 51548 30996 51604 31006
rect 51436 30994 51604 30996
rect 51436 30942 51550 30994
rect 51602 30942 51604 30994
rect 51436 30940 51604 30942
rect 51324 30902 51380 30940
rect 51548 30930 51604 30940
rect 51212 30716 51604 30772
rect 50988 29596 51268 29652
rect 50428 29586 50484 29596
rect 50316 28924 50820 28980
rect 50316 28532 50372 28542
rect 50316 28082 50372 28476
rect 50316 28030 50318 28082
rect 50370 28030 50372 28082
rect 50316 28018 50372 28030
rect 49980 27020 50148 27076
rect 50652 27970 50708 27982
rect 50652 27918 50654 27970
rect 50706 27918 50708 27970
rect 49980 26852 50036 27020
rect 50652 26964 50708 27918
rect 50652 26898 50708 26908
rect 49980 26796 50148 26852
rect 49756 26012 50036 26068
rect 49512 25900 49776 25910
rect 49568 25844 49616 25900
rect 49672 25844 49720 25900
rect 49512 25834 49776 25844
rect 49756 25620 49812 25630
rect 49420 25618 49812 25620
rect 49420 25566 49758 25618
rect 49810 25566 49812 25618
rect 49420 25564 49812 25566
rect 49420 25506 49476 25564
rect 49756 25554 49812 25564
rect 49420 25454 49422 25506
rect 49474 25454 49476 25506
rect 49420 25442 49476 25454
rect 49868 25282 49924 25294
rect 49868 25230 49870 25282
rect 49922 25230 49924 25282
rect 49532 24948 49588 24958
rect 49868 24948 49924 25230
rect 49308 24946 49924 24948
rect 49308 24894 49534 24946
rect 49586 24894 49924 24946
rect 49308 24892 49924 24894
rect 49532 24882 49588 24892
rect 49512 24332 49776 24342
rect 49568 24276 49616 24332
rect 49672 24276 49720 24332
rect 49512 24266 49776 24276
rect 49420 24052 49476 24062
rect 49420 23958 49476 23996
rect 49420 23044 49476 23054
rect 48748 22540 49252 22596
rect 49308 22988 49420 23044
rect 48188 22372 48244 22382
rect 48188 22370 48356 22372
rect 48188 22318 48190 22370
rect 48242 22318 48356 22370
rect 48188 22316 48356 22318
rect 48188 22306 48244 22316
rect 48076 21534 48078 21586
rect 48130 21534 48132 21586
rect 48076 21522 48132 21534
rect 47852 21474 47908 21486
rect 47852 21422 47854 21474
rect 47906 21422 47908 21474
rect 47852 20804 47908 21422
rect 47852 20738 47908 20748
rect 47628 20578 47796 20580
rect 47628 20526 47630 20578
rect 47682 20526 47796 20578
rect 47628 20524 47796 20526
rect 47516 19122 47572 19134
rect 47516 19070 47518 19122
rect 47570 19070 47572 19122
rect 47516 19012 47572 19070
rect 47516 18946 47572 18956
rect 47628 18228 47684 20524
rect 48188 20468 48244 20478
rect 48188 18564 48244 20412
rect 48300 20244 48356 22316
rect 48636 21476 48692 21486
rect 48636 20692 48692 21420
rect 48748 21364 48804 22540
rect 48972 22370 49028 22382
rect 48972 22318 48974 22370
rect 49026 22318 49028 22370
rect 48860 21588 48916 21598
rect 48860 21494 48916 21532
rect 48748 21308 48916 21364
rect 48748 20804 48804 20814
rect 48748 20710 48804 20748
rect 48636 20580 48692 20636
rect 48636 20524 48804 20580
rect 48300 20188 48692 20244
rect 48636 19796 48692 20188
rect 48748 20130 48804 20524
rect 48748 20078 48750 20130
rect 48802 20078 48804 20130
rect 48748 20066 48804 20078
rect 48860 20244 48916 21308
rect 48860 20130 48916 20188
rect 48860 20078 48862 20130
rect 48914 20078 48916 20130
rect 48860 20066 48916 20078
rect 48636 19740 48804 19796
rect 48188 18508 48356 18564
rect 47628 18162 47684 18172
rect 48188 18338 48244 18350
rect 48188 18286 48190 18338
rect 48242 18286 48244 18338
rect 47404 17714 47460 17724
rect 47964 17668 48020 17678
rect 48188 17668 48244 18286
rect 47068 17602 47124 17612
rect 47852 17666 48244 17668
rect 47852 17614 47966 17666
rect 48018 17614 48244 17666
rect 47852 17612 48244 17614
rect 47180 17556 47236 17566
rect 47628 17556 47684 17566
rect 47180 17554 47684 17556
rect 47180 17502 47182 17554
rect 47234 17502 47630 17554
rect 47682 17502 47684 17554
rect 47180 17500 47684 17502
rect 47180 17490 47236 17500
rect 47628 17490 47684 17500
rect 46620 17388 46788 17444
rect 46172 17042 46228 17052
rect 46620 17220 46676 17230
rect 46060 16942 46062 16994
rect 46114 16942 46116 16994
rect 46060 16930 46116 16942
rect 46508 16770 46564 16782
rect 46508 16718 46510 16770
rect 46562 16718 46564 16770
rect 45836 16212 45892 16222
rect 45724 16210 45892 16212
rect 45724 16158 45838 16210
rect 45890 16158 45892 16210
rect 45724 16156 45892 16158
rect 45612 15202 45668 15214
rect 45612 15150 45614 15202
rect 45666 15150 45668 15202
rect 45164 15092 45332 15148
rect 45388 15092 45556 15148
rect 45164 13858 45220 13870
rect 45164 13806 45166 13858
rect 45218 13806 45220 13858
rect 45164 12290 45220 13806
rect 45276 13412 45332 15092
rect 45276 13346 45332 13356
rect 45388 13746 45444 13758
rect 45388 13694 45390 13746
rect 45442 13694 45444 13746
rect 45388 13186 45444 13694
rect 45388 13134 45390 13186
rect 45442 13134 45444 13186
rect 45388 13122 45444 13134
rect 45164 12238 45166 12290
rect 45218 12238 45220 12290
rect 45164 12226 45220 12238
rect 45276 12964 45332 12974
rect 45276 10052 45332 12908
rect 45500 12292 45556 15092
rect 45612 14420 45668 15150
rect 45612 14354 45668 14364
rect 45612 14196 45668 14206
rect 45612 12740 45668 14140
rect 45724 13860 45780 16156
rect 45836 16146 45892 16156
rect 46396 15876 46452 15886
rect 46396 15782 46452 15820
rect 46060 15540 46116 15550
rect 46060 15446 46116 15484
rect 46508 15148 46564 16718
rect 46284 15092 46564 15148
rect 46060 14420 46116 14430
rect 45724 13804 45892 13860
rect 45724 13524 45780 13534
rect 45724 13186 45780 13468
rect 45724 13134 45726 13186
rect 45778 13134 45780 13186
rect 45724 13122 45780 13134
rect 45612 12674 45668 12684
rect 45500 12226 45556 12236
rect 45276 9958 45332 9996
rect 45500 11172 45556 11182
rect 45500 10500 45556 11116
rect 45388 8930 45444 8942
rect 45388 8878 45390 8930
rect 45442 8878 45444 8930
rect 45388 8428 45444 8878
rect 45164 8372 45444 8428
rect 45164 8146 45220 8372
rect 45164 8094 45166 8146
rect 45218 8094 45220 8146
rect 45164 8082 45220 8094
rect 45276 5348 45332 5358
rect 45276 5254 45332 5292
rect 45052 4722 45108 4732
rect 44716 3490 44772 3500
rect 40460 3390 40462 3442
rect 40514 3390 40516 3442
rect 39340 3378 39396 3388
rect 40124 3332 40292 3388
rect 40460 3378 40516 3390
rect 43932 3444 43988 3482
rect 44156 3444 44212 3454
rect 43932 3442 44212 3444
rect 43932 3390 43934 3442
rect 43986 3390 44158 3442
rect 44210 3390 44212 3442
rect 43932 3388 44212 3390
rect 39852 3164 40116 3174
rect 39908 3108 39956 3164
rect 40012 3108 40060 3164
rect 39852 3098 40116 3108
rect 40236 2324 40292 3332
rect 39900 2268 40292 2324
rect 39900 800 39956 2268
rect 43932 800 43988 3388
rect 44156 3378 44212 3388
rect 44492 3444 44548 3482
rect 45500 3388 45556 10444
rect 45612 7140 45668 7150
rect 45668 7084 45780 7140
rect 45612 7074 45668 7084
rect 45724 6580 45780 7084
rect 45724 5236 45780 6524
rect 45724 5122 45780 5180
rect 45724 5070 45726 5122
rect 45778 5070 45780 5122
rect 45724 5058 45780 5070
rect 45836 5796 45892 13804
rect 45948 13636 46004 13646
rect 45948 13542 46004 13580
rect 46060 13412 46116 14364
rect 45948 13356 46116 13412
rect 45948 11172 46004 13356
rect 46284 13188 46340 15092
rect 46620 14644 46676 17164
rect 46732 16212 46788 17388
rect 46844 17442 46900 17454
rect 46844 17390 46846 17442
rect 46898 17390 46900 17442
rect 46844 17108 46900 17390
rect 46844 17042 46900 17052
rect 46956 17444 47012 17454
rect 46956 16884 47012 17388
rect 46956 16790 47012 16828
rect 47404 16882 47460 16894
rect 47404 16830 47406 16882
rect 47458 16830 47460 16882
rect 46844 16212 46900 16222
rect 46732 16210 46900 16212
rect 46732 16158 46846 16210
rect 46898 16158 46900 16210
rect 46732 16156 46900 16158
rect 46508 14588 46676 14644
rect 46396 13972 46452 13982
rect 46396 13878 46452 13916
rect 46396 13188 46452 13198
rect 46284 13132 46396 13188
rect 46396 13122 46452 13132
rect 46396 12962 46452 12974
rect 46396 12910 46398 12962
rect 46450 12910 46452 12962
rect 46284 12852 46340 12862
rect 45948 11106 46004 11116
rect 46060 12850 46340 12852
rect 46060 12798 46286 12850
rect 46338 12798 46340 12850
rect 46060 12796 46340 12798
rect 46060 10948 46116 12796
rect 46284 12786 46340 12796
rect 46396 12852 46452 12910
rect 46396 12786 46452 12796
rect 45948 10892 46116 10948
rect 45948 9714 46004 10892
rect 46396 10836 46452 10846
rect 46508 10836 46564 14588
rect 46732 13858 46788 13870
rect 46732 13806 46734 13858
rect 46786 13806 46788 13858
rect 46732 13524 46788 13806
rect 46732 13458 46788 13468
rect 46844 13412 46900 16156
rect 47404 15540 47460 16830
rect 47628 16884 47684 16894
rect 47628 16098 47684 16828
rect 47628 16046 47630 16098
rect 47682 16046 47684 16098
rect 47628 16034 47684 16046
rect 47852 15876 47908 17612
rect 47964 17602 48020 17612
rect 48300 17444 48356 18508
rect 48748 18450 48804 19740
rect 48972 18564 49028 22318
rect 49308 21588 49364 22988
rect 49420 22950 49476 22988
rect 49512 22764 49776 22774
rect 49568 22708 49616 22764
rect 49672 22708 49720 22764
rect 49512 22698 49776 22708
rect 49756 22146 49812 22158
rect 49756 22094 49758 22146
rect 49810 22094 49812 22146
rect 49756 21812 49812 22094
rect 49756 21588 49812 21756
rect 49196 21586 49812 21588
rect 49196 21534 49310 21586
rect 49362 21534 49812 21586
rect 49196 21532 49812 21534
rect 49868 21588 49924 21598
rect 49084 20916 49140 20926
rect 49196 20916 49252 21532
rect 49308 21522 49364 21532
rect 49512 21196 49776 21206
rect 49568 21140 49616 21196
rect 49672 21140 49720 21196
rect 49512 21130 49776 21140
rect 49868 21028 49924 21532
rect 49140 20860 49252 20916
rect 49756 20972 49924 21028
rect 49084 20850 49140 20860
rect 49084 20690 49140 20702
rect 49084 20638 49086 20690
rect 49138 20638 49140 20690
rect 49084 20242 49140 20638
rect 49084 20190 49086 20242
rect 49138 20190 49140 20242
rect 49084 20178 49140 20190
rect 49308 20578 49364 20590
rect 49308 20526 49310 20578
rect 49362 20526 49364 20578
rect 48972 18470 49028 18508
rect 49196 19012 49252 19022
rect 48748 18398 48750 18450
rect 48802 18398 48804 18450
rect 48636 18340 48692 18350
rect 48636 17554 48692 18284
rect 48748 18004 48804 18398
rect 48748 17948 49140 18004
rect 48748 17780 48804 17790
rect 48748 17666 48804 17724
rect 48748 17614 48750 17666
rect 48802 17614 48804 17666
rect 48748 17602 48804 17614
rect 49084 17668 49140 17948
rect 49196 17780 49252 18956
rect 49308 18228 49364 20526
rect 49420 20244 49476 20254
rect 49756 20244 49812 20972
rect 49868 20804 49924 20814
rect 49980 20804 50036 26012
rect 50092 25732 50148 26796
rect 50428 26850 50484 26862
rect 50428 26798 50430 26850
rect 50482 26798 50484 26850
rect 50204 26292 50260 26302
rect 50204 26198 50260 26236
rect 50428 26292 50484 26798
rect 50540 26852 50596 26862
rect 50540 26514 50596 26796
rect 50540 26462 50542 26514
rect 50594 26462 50596 26514
rect 50540 26450 50596 26462
rect 50764 26514 50820 28924
rect 50876 27972 50932 27982
rect 50876 27858 50932 27916
rect 50876 27806 50878 27858
rect 50930 27806 50932 27858
rect 50876 27794 50932 27806
rect 50764 26462 50766 26514
rect 50818 26462 50820 26514
rect 50764 26450 50820 26462
rect 50988 27748 51044 27758
rect 50428 26226 50484 26236
rect 50652 26292 50708 26302
rect 50652 26290 50820 26292
rect 50652 26238 50654 26290
rect 50706 26238 50820 26290
rect 50652 26236 50820 26238
rect 50652 26226 50708 26236
rect 50652 25844 50708 25854
rect 50540 25788 50652 25844
rect 50092 25730 50484 25732
rect 50092 25678 50094 25730
rect 50146 25678 50484 25730
rect 50092 25676 50484 25678
rect 50092 25666 50148 25676
rect 50428 25506 50484 25676
rect 50428 25454 50430 25506
rect 50482 25454 50484 25506
rect 50428 25442 50484 25454
rect 50316 24276 50372 24286
rect 50092 23380 50148 23390
rect 50092 23286 50148 23324
rect 50316 23156 50372 24220
rect 49868 20802 49980 20804
rect 49868 20750 49870 20802
rect 49922 20750 49980 20802
rect 49868 20748 49980 20750
rect 49868 20738 49924 20748
rect 49980 20710 50036 20748
rect 50092 23100 50372 23156
rect 50092 22372 50148 23100
rect 49868 20244 49924 20254
rect 49756 20242 49924 20244
rect 49756 20190 49870 20242
rect 49922 20190 49924 20242
rect 49756 20188 49924 20190
rect 49420 20130 49476 20188
rect 49420 20078 49422 20130
rect 49474 20078 49476 20130
rect 49420 20066 49476 20078
rect 49868 20020 49924 20188
rect 49868 19954 49924 19964
rect 50092 19796 50148 22316
rect 50204 22482 50260 22494
rect 50204 22430 50206 22482
rect 50258 22430 50260 22482
rect 50204 22260 50260 22430
rect 50204 22194 50260 22204
rect 50316 21812 50372 21822
rect 50316 21718 50372 21756
rect 50316 20804 50372 20814
rect 50540 20804 50596 25788
rect 50652 25778 50708 25788
rect 50764 25396 50820 26236
rect 50764 25302 50820 25340
rect 50876 26290 50932 26302
rect 50876 26238 50878 26290
rect 50930 26238 50932 26290
rect 50764 25060 50820 25070
rect 50764 24610 50820 25004
rect 50764 24558 50766 24610
rect 50818 24558 50820 24610
rect 50764 24500 50820 24558
rect 50764 24434 50820 24444
rect 50876 24052 50932 26238
rect 50988 24276 51044 27692
rect 51100 26964 51156 26974
rect 51100 26402 51156 26908
rect 51100 26350 51102 26402
rect 51154 26350 51156 26402
rect 51100 26338 51156 26350
rect 51212 25844 51268 29596
rect 51436 29204 51492 29214
rect 51436 28642 51492 29148
rect 51436 28590 51438 28642
rect 51490 28590 51492 28642
rect 51436 28578 51492 28590
rect 51436 28420 51492 28430
rect 51436 28082 51492 28364
rect 51436 28030 51438 28082
rect 51490 28030 51492 28082
rect 51436 28018 51492 28030
rect 51212 25778 51268 25788
rect 51100 24722 51156 24734
rect 51100 24670 51102 24722
rect 51154 24670 51156 24722
rect 51100 24500 51156 24670
rect 51100 24434 51156 24444
rect 50988 24220 51268 24276
rect 50876 23986 50932 23996
rect 50764 23714 50820 23726
rect 50764 23662 50766 23714
rect 50818 23662 50820 23714
rect 50652 23492 50708 23502
rect 50652 23154 50708 23436
rect 50652 23102 50654 23154
rect 50706 23102 50708 23154
rect 50652 22372 50708 23102
rect 50764 23156 50820 23662
rect 51100 23380 51156 23390
rect 50988 23156 51044 23166
rect 50764 23154 51044 23156
rect 50764 23102 50990 23154
rect 51042 23102 51044 23154
rect 50764 23100 51044 23102
rect 50988 23044 51044 23100
rect 50988 22978 51044 22988
rect 51100 22482 51156 23324
rect 51100 22430 51102 22482
rect 51154 22430 51156 22482
rect 51100 22418 51156 22430
rect 50652 22306 50708 22316
rect 50876 22148 50932 22158
rect 50876 22146 51044 22148
rect 50876 22094 50878 22146
rect 50930 22094 51044 22146
rect 50876 22092 51044 22094
rect 50876 22082 50932 22092
rect 50876 21812 50932 21822
rect 50876 21718 50932 21756
rect 50988 21588 51044 22092
rect 51212 21810 51268 24220
rect 51324 23716 51380 23726
rect 51324 23380 51380 23660
rect 51324 23378 51492 23380
rect 51324 23326 51326 23378
rect 51378 23326 51492 23378
rect 51324 23324 51492 23326
rect 51324 23314 51380 23324
rect 51324 23156 51380 23166
rect 51324 22594 51380 23100
rect 51324 22542 51326 22594
rect 51378 22542 51380 22594
rect 51324 22530 51380 22542
rect 51212 21758 51214 21810
rect 51266 21758 51268 21810
rect 51212 21746 51268 21758
rect 51324 22036 51380 22046
rect 51324 21700 51380 21980
rect 51436 21812 51492 23324
rect 51436 21746 51492 21756
rect 50988 21586 51268 21588
rect 50988 21534 50990 21586
rect 51042 21534 51268 21586
rect 50988 21532 51268 21534
rect 50988 21522 51044 21532
rect 50876 21476 50932 21486
rect 50204 20692 50260 20702
rect 50204 20598 50260 20636
rect 50316 20690 50372 20748
rect 50316 20638 50318 20690
rect 50370 20638 50372 20690
rect 50316 20626 50372 20638
rect 50428 20748 50596 20804
rect 50764 21474 50932 21476
rect 50764 21422 50878 21474
rect 50930 21422 50932 21474
rect 50764 21420 50932 21422
rect 50764 20802 50820 21420
rect 50876 21410 50932 21420
rect 50764 20750 50766 20802
rect 50818 20750 50820 20802
rect 50428 20020 50484 20748
rect 50764 20738 50820 20750
rect 50876 20690 50932 20702
rect 50876 20638 50878 20690
rect 50930 20638 50932 20690
rect 50540 20580 50596 20590
rect 50876 20580 50932 20638
rect 50540 20578 50932 20580
rect 50540 20526 50542 20578
rect 50594 20526 50932 20578
rect 50540 20524 50932 20526
rect 50988 20692 51044 20702
rect 50540 20514 50596 20524
rect 50988 20130 51044 20636
rect 50988 20078 50990 20130
rect 51042 20078 51044 20130
rect 50988 20066 51044 20078
rect 51100 20578 51156 20590
rect 51100 20526 51102 20578
rect 51154 20526 51156 20578
rect 50876 20020 50932 20030
rect 50428 20018 50932 20020
rect 50428 19966 50878 20018
rect 50930 19966 50932 20018
rect 50428 19964 50932 19966
rect 49868 19740 50148 19796
rect 50316 19908 50372 19918
rect 49512 19628 49776 19638
rect 49568 19572 49616 19628
rect 49672 19572 49720 19628
rect 49512 19562 49776 19572
rect 49420 18900 49476 18910
rect 49420 18338 49476 18844
rect 49420 18286 49422 18338
rect 49474 18286 49476 18338
rect 49420 18274 49476 18286
rect 49308 18162 49364 18172
rect 49512 18060 49776 18070
rect 49568 18004 49616 18060
rect 49672 18004 49720 18060
rect 49512 17994 49776 18004
rect 49308 17780 49364 17790
rect 49196 17724 49308 17780
rect 49308 17686 49364 17724
rect 49084 17612 49252 17668
rect 48636 17502 48638 17554
rect 48690 17502 48692 17554
rect 48636 17490 48692 17502
rect 47964 17388 48356 17444
rect 47964 16996 48020 17388
rect 48636 17108 48692 17118
rect 47964 16994 48132 16996
rect 47964 16942 47966 16994
rect 48018 16942 48132 16994
rect 47964 16940 48132 16942
rect 47964 16930 48020 16940
rect 47404 15474 47460 15484
rect 47628 15820 47908 15876
rect 47292 15092 47348 15102
rect 46956 14532 47012 14542
rect 46956 14530 47236 14532
rect 46956 14478 46958 14530
rect 47010 14478 47236 14530
rect 46956 14476 47236 14478
rect 46956 14466 47012 14476
rect 46844 13356 47012 13412
rect 46844 13188 46900 13198
rect 46732 12740 46788 12750
rect 46060 10834 46564 10836
rect 46060 10782 46398 10834
rect 46450 10782 46564 10834
rect 46060 10780 46564 10782
rect 46620 12292 46676 12302
rect 46060 9826 46116 10780
rect 46396 10770 46452 10780
rect 46060 9774 46062 9826
rect 46114 9774 46116 9826
rect 46060 9762 46116 9774
rect 46620 9828 46676 12236
rect 46732 11506 46788 12684
rect 46732 11454 46734 11506
rect 46786 11454 46788 11506
rect 46732 11442 46788 11454
rect 46732 9828 46788 9838
rect 46620 9826 46788 9828
rect 46620 9774 46734 9826
rect 46786 9774 46788 9826
rect 46620 9772 46788 9774
rect 45948 9662 45950 9714
rect 46002 9662 46004 9714
rect 45948 9156 46004 9662
rect 45948 9090 46004 9100
rect 46172 9716 46228 9726
rect 46172 9044 46228 9660
rect 46172 9042 46564 9044
rect 46172 8990 46174 9042
rect 46226 8990 46564 9042
rect 46172 8988 46564 8990
rect 46172 8978 46228 8988
rect 46508 8258 46564 8988
rect 46508 8206 46510 8258
rect 46562 8206 46564 8258
rect 46508 8194 46564 8206
rect 44492 3378 44548 3388
rect 45388 3332 45556 3388
rect 45836 3388 45892 5740
rect 45948 7252 46004 7262
rect 45948 5794 46004 7196
rect 46620 6692 46676 9772
rect 46732 9762 46788 9772
rect 46844 7588 46900 13132
rect 46956 12852 47012 13356
rect 47068 12964 47124 12974
rect 47068 12870 47124 12908
rect 46956 12786 47012 12796
rect 47180 11732 47236 14476
rect 47292 13972 47348 15036
rect 47516 14420 47572 14430
rect 47516 14326 47572 14364
rect 47292 13746 47348 13916
rect 47292 13694 47294 13746
rect 47346 13694 47348 13746
rect 47292 13682 47348 13694
rect 47628 13746 47684 15820
rect 47964 15764 48020 15774
rect 47740 15316 47796 15326
rect 47964 15316 48020 15708
rect 47740 15314 48020 15316
rect 47740 15262 47742 15314
rect 47794 15262 48020 15314
rect 47740 15260 48020 15262
rect 47740 15250 47796 15260
rect 47964 14308 48020 15260
rect 47852 13970 47908 13982
rect 47852 13918 47854 13970
rect 47906 13918 47908 13970
rect 47852 13860 47908 13918
rect 47964 13970 48020 14252
rect 47964 13918 47966 13970
rect 48018 13918 48020 13970
rect 47964 13906 48020 13918
rect 47852 13794 47908 13804
rect 47628 13694 47630 13746
rect 47682 13694 47684 13746
rect 47292 13412 47348 13422
rect 47292 12066 47348 13356
rect 47628 12180 47684 13694
rect 47628 12114 47684 12124
rect 47740 13188 47796 13198
rect 47292 12014 47294 12066
rect 47346 12014 47348 12066
rect 47292 12002 47348 12014
rect 47180 11666 47236 11676
rect 47516 9828 47572 9838
rect 47068 9826 47572 9828
rect 47068 9774 47518 9826
rect 47570 9774 47572 9826
rect 47068 9772 47572 9774
rect 47068 9716 47124 9772
rect 47516 9762 47572 9772
rect 47068 9622 47124 9660
rect 47740 9492 47796 13132
rect 47852 12852 47908 12862
rect 47852 12402 47908 12796
rect 47852 12350 47854 12402
rect 47906 12350 47908 12402
rect 47852 12338 47908 12350
rect 47852 11170 47908 11182
rect 47852 11118 47854 11170
rect 47906 11118 47908 11170
rect 47852 10722 47908 11118
rect 47852 10670 47854 10722
rect 47906 10670 47908 10722
rect 47852 10658 47908 10670
rect 47740 9426 47796 9436
rect 48076 9268 48132 16940
rect 48188 16660 48244 16670
rect 48188 16212 48244 16604
rect 48188 16210 48580 16212
rect 48188 16158 48190 16210
rect 48242 16158 48580 16210
rect 48188 16156 48580 16158
rect 48188 16146 48244 16156
rect 48188 15202 48244 15214
rect 48188 15150 48190 15202
rect 48242 15150 48244 15202
rect 48188 14420 48244 15150
rect 48412 15204 48468 15214
rect 48300 14532 48356 14542
rect 48300 14438 48356 14476
rect 48188 14354 48244 14364
rect 48188 13748 48244 13758
rect 48188 11618 48244 13692
rect 48300 13636 48356 13646
rect 48412 13636 48468 15148
rect 48356 13580 48468 13636
rect 48300 12962 48356 13580
rect 48300 12910 48302 12962
rect 48354 12910 48356 12962
rect 48300 12898 48356 12910
rect 48188 11566 48190 11618
rect 48242 11566 48244 11618
rect 48188 11284 48244 11566
rect 48188 11218 48244 11228
rect 48524 11508 48580 16156
rect 48636 15764 48692 17052
rect 48972 16884 49028 16894
rect 48860 16828 48972 16884
rect 48860 16100 48916 16828
rect 48972 16790 49028 16828
rect 48860 16098 49028 16100
rect 48860 16046 48862 16098
rect 48914 16046 49028 16098
rect 48860 16044 49028 16046
rect 48860 16034 48916 16044
rect 48636 15698 48692 15708
rect 48860 15538 48916 15550
rect 48860 15486 48862 15538
rect 48914 15486 48916 15538
rect 48748 15314 48804 15326
rect 48748 15262 48750 15314
rect 48802 15262 48804 15314
rect 48636 12962 48692 12974
rect 48636 12910 48638 12962
rect 48690 12910 48692 12962
rect 48636 12740 48692 12910
rect 48636 12674 48692 12684
rect 48748 11956 48804 15262
rect 48860 14644 48916 15486
rect 48972 15092 49028 16044
rect 48972 15026 49028 15036
rect 49084 15538 49140 15550
rect 49084 15486 49086 15538
rect 49138 15486 49140 15538
rect 48860 14578 48916 14588
rect 48860 14196 48916 14206
rect 48860 13300 48916 14140
rect 49084 13746 49140 15486
rect 49196 14642 49252 17612
rect 49512 16492 49776 16502
rect 49568 16436 49616 16492
rect 49672 16436 49720 16492
rect 49512 16426 49776 16436
rect 49644 16212 49700 16222
rect 49196 14590 49198 14642
rect 49250 14590 49252 14642
rect 49196 14578 49252 14590
rect 49308 15986 49364 15998
rect 49308 15934 49310 15986
rect 49362 15934 49364 15986
rect 49308 14532 49364 15934
rect 49644 15314 49700 16156
rect 49644 15262 49646 15314
rect 49698 15262 49700 15314
rect 49644 15250 49700 15262
rect 49512 14924 49776 14934
rect 49568 14868 49616 14924
rect 49672 14868 49720 14924
rect 49512 14858 49776 14868
rect 49308 14466 49364 14476
rect 49084 13694 49086 13746
rect 49138 13694 49140 13746
rect 49084 13682 49140 13694
rect 49868 13634 49924 19740
rect 50316 19348 50372 19852
rect 50428 19908 50484 19964
rect 50876 19954 50932 19964
rect 50428 19842 50484 19852
rect 50316 19282 50372 19292
rect 50204 18676 50260 18686
rect 49868 13582 49870 13634
rect 49922 13582 49924 13634
rect 49868 13570 49924 13582
rect 49980 18340 50036 18350
rect 49512 13356 49776 13366
rect 49568 13300 49616 13356
rect 49672 13300 49720 13356
rect 49512 13290 49776 13300
rect 48860 13234 48916 13244
rect 48972 12964 49028 12974
rect 48972 12404 49028 12908
rect 48972 12338 49028 12348
rect 48748 11890 48804 11900
rect 49512 11788 49776 11798
rect 49568 11732 49616 11788
rect 49672 11732 49720 11788
rect 49512 11722 49776 11732
rect 48524 11282 48580 11452
rect 49756 11396 49812 11406
rect 49980 11396 50036 18284
rect 50092 16884 50148 16894
rect 50092 16790 50148 16828
rect 50204 16324 50260 18620
rect 51100 18340 51156 20526
rect 51100 18274 51156 18284
rect 50988 17444 51044 17454
rect 50764 17442 51044 17444
rect 50764 17390 50990 17442
rect 51042 17390 51044 17442
rect 50764 17388 51044 17390
rect 50764 16994 50820 17388
rect 50988 17378 51044 17388
rect 50764 16942 50766 16994
rect 50818 16942 50820 16994
rect 50764 16930 50820 16942
rect 50204 16258 50260 16268
rect 50988 16212 51044 16222
rect 50988 16098 51044 16156
rect 50988 16046 50990 16098
rect 51042 16046 51044 16098
rect 50988 16034 51044 16046
rect 50988 15540 51044 15550
rect 50988 15446 51044 15484
rect 50092 15426 50148 15438
rect 50092 15374 50094 15426
rect 50146 15374 50148 15426
rect 50092 13748 50148 15374
rect 50764 15428 50820 15438
rect 50764 14980 50820 15372
rect 50876 14980 50932 14990
rect 50764 14924 50876 14980
rect 50316 14532 50372 14542
rect 50316 14438 50372 14476
rect 50764 14418 50820 14430
rect 50764 14366 50766 14418
rect 50818 14366 50820 14418
rect 50764 14196 50820 14366
rect 50764 14130 50820 14140
rect 50428 13860 50484 13870
rect 50428 13766 50484 13804
rect 50092 13682 50148 13692
rect 50204 13746 50260 13758
rect 50204 13694 50206 13746
rect 50258 13694 50260 13746
rect 50204 13074 50260 13694
rect 50204 13022 50206 13074
rect 50258 13022 50260 13074
rect 50204 13010 50260 13022
rect 50876 12850 50932 14924
rect 51100 14644 51156 14654
rect 51100 14530 51156 14588
rect 51100 14478 51102 14530
rect 51154 14478 51156 14530
rect 51100 14466 51156 14478
rect 50876 12798 50878 12850
rect 50930 12798 50932 12850
rect 50876 12786 50932 12798
rect 51100 12964 51156 12974
rect 50652 12178 50708 12190
rect 50652 12126 50654 12178
rect 50706 12126 50708 12178
rect 49756 11394 49980 11396
rect 49756 11342 49758 11394
rect 49810 11342 49980 11394
rect 49756 11340 49980 11342
rect 49756 11330 49812 11340
rect 49980 11302 50036 11340
rect 50092 12068 50148 12078
rect 48524 11230 48526 11282
rect 48578 11230 48580 11282
rect 48524 11218 48580 11230
rect 48860 11282 48916 11294
rect 48860 11230 48862 11282
rect 48914 11230 48916 11282
rect 48860 11172 48916 11230
rect 49420 11172 49476 11182
rect 48860 11170 49476 11172
rect 48860 11118 49422 11170
rect 49474 11118 49476 11170
rect 48860 11116 49476 11118
rect 48748 11060 48804 11070
rect 48188 10722 48244 10734
rect 48188 10670 48190 10722
rect 48242 10670 48244 10722
rect 48188 9940 48244 10670
rect 48300 9940 48356 9950
rect 48188 9938 48356 9940
rect 48188 9886 48302 9938
rect 48354 9886 48356 9938
rect 48188 9884 48356 9886
rect 48300 9874 48356 9884
rect 48748 9828 48804 11004
rect 48748 9762 48804 9772
rect 47516 9212 48076 9268
rect 47180 9156 47236 9166
rect 47180 9062 47236 9100
rect 47516 9154 47572 9212
rect 48076 9202 48132 9212
rect 47516 9102 47518 9154
rect 47570 9102 47572 9154
rect 47516 9090 47572 9102
rect 48748 9154 48804 9166
rect 48748 9102 48750 9154
rect 48802 9102 48804 9154
rect 47740 9044 47796 9054
rect 47740 8950 47796 8988
rect 48076 9044 48132 9054
rect 48076 8950 48132 8988
rect 47292 8372 47348 8382
rect 47292 8278 47348 8316
rect 48748 8372 48804 9102
rect 48860 9156 48916 11116
rect 49420 11106 49476 11116
rect 50092 10948 50148 12012
rect 50204 11508 50260 11518
rect 50204 11414 50260 11452
rect 50092 10882 50148 10892
rect 50428 11284 50484 11294
rect 49512 10220 49776 10230
rect 49568 10164 49616 10220
rect 49672 10164 49720 10220
rect 49512 10154 49776 10164
rect 48860 9090 48916 9100
rect 49308 9940 49364 9950
rect 48972 9044 49028 9054
rect 48972 8950 49028 8988
rect 49308 8932 49364 9884
rect 50428 9938 50484 11228
rect 50428 9886 50430 9938
rect 50482 9886 50484 9938
rect 50428 9874 50484 9886
rect 50652 10612 50708 12126
rect 49644 9268 49700 9278
rect 49644 9174 49700 9212
rect 50540 8932 50596 8942
rect 48748 8306 48804 8316
rect 48860 8484 48916 8494
rect 46844 7522 46900 7532
rect 47404 7812 47460 7822
rect 46620 6626 46676 6636
rect 45948 5742 45950 5794
rect 46002 5742 46004 5794
rect 45948 5730 46004 5742
rect 46508 5348 46564 5358
rect 46060 5012 46116 5022
rect 46060 4918 46116 4956
rect 46508 4226 46564 5292
rect 47068 5348 47124 5358
rect 46620 5236 46676 5246
rect 46620 5142 46676 5180
rect 47068 5234 47124 5292
rect 47068 5182 47070 5234
rect 47122 5182 47124 5234
rect 47068 5170 47124 5182
rect 46508 4174 46510 4226
rect 46562 4174 46564 4226
rect 46508 4162 46564 4174
rect 47404 3444 47460 7756
rect 48860 7700 48916 8428
rect 49308 8372 49364 8876
rect 50428 8903 50540 8932
rect 50428 8851 50430 8903
rect 50482 8876 50540 8903
rect 50482 8851 50484 8876
rect 50540 8866 50596 8876
rect 50428 8839 50484 8851
rect 49512 8652 49776 8662
rect 49568 8596 49616 8652
rect 49672 8596 49720 8652
rect 49512 8586 49776 8596
rect 49420 8372 49476 8382
rect 49308 8370 49476 8372
rect 49308 8318 49422 8370
rect 49474 8318 49476 8370
rect 49308 8316 49476 8318
rect 49420 8306 49476 8316
rect 48860 7634 48916 7644
rect 48748 7252 48804 7262
rect 48636 6468 48692 6478
rect 47964 6466 48692 6468
rect 47964 6414 48638 6466
rect 48690 6414 48692 6466
rect 47964 6412 48692 6414
rect 47852 5908 47908 5918
rect 47852 5122 47908 5852
rect 47964 5906 48020 6412
rect 48636 6402 48692 6412
rect 48748 6132 48804 7196
rect 49512 7084 49776 7094
rect 49568 7028 49616 7084
rect 49672 7028 49720 7084
rect 49512 7018 49776 7028
rect 48972 6916 49028 6926
rect 48972 6822 49028 6860
rect 49196 6578 49252 6590
rect 49196 6526 49198 6578
rect 49250 6526 49252 6578
rect 49196 6468 49252 6526
rect 49756 6580 49812 6590
rect 50428 6580 50484 6590
rect 49756 6578 49924 6580
rect 49756 6526 49758 6578
rect 49810 6526 49924 6578
rect 49756 6524 49924 6526
rect 49756 6514 49812 6524
rect 49196 6402 49252 6412
rect 48748 6066 48804 6076
rect 48188 6020 48244 6030
rect 48188 5926 48244 5964
rect 49532 6020 49588 6030
rect 49532 5926 49588 5964
rect 47964 5854 47966 5906
rect 48018 5854 48020 5906
rect 47964 5842 48020 5854
rect 48860 5908 48916 5918
rect 48860 5814 48916 5852
rect 49512 5516 49776 5526
rect 49568 5460 49616 5516
rect 49672 5460 49720 5516
rect 49512 5450 49776 5460
rect 47852 5070 47854 5122
rect 47906 5070 47908 5122
rect 47852 5058 47908 5070
rect 48524 5012 48580 5022
rect 48188 5010 48580 5012
rect 48188 4958 48526 5010
rect 48578 4958 48580 5010
rect 48188 4956 48580 4958
rect 48188 4562 48244 4956
rect 48524 4946 48580 4956
rect 49868 5012 49924 6524
rect 50428 6486 50484 6524
rect 48188 4510 48190 4562
rect 48242 4510 48244 4562
rect 48188 4498 48244 4510
rect 49196 4900 49252 4910
rect 47964 4340 48020 4350
rect 47964 4246 48020 4284
rect 48860 4340 48916 4350
rect 48860 4246 48916 4284
rect 49196 4338 49252 4844
rect 49420 4788 49476 4798
rect 49420 4452 49476 4732
rect 49420 4358 49476 4396
rect 49868 4450 49924 4956
rect 50652 5234 50708 10556
rect 50876 10610 50932 10622
rect 50876 10558 50878 10610
rect 50930 10558 50932 10610
rect 50876 6468 50932 10558
rect 50988 9828 51044 9838
rect 50988 9492 51044 9772
rect 50988 9426 51044 9436
rect 51100 9714 51156 12908
rect 51100 9662 51102 9714
rect 51154 9662 51156 9714
rect 51100 8932 51156 9662
rect 51100 8866 51156 8876
rect 50876 6402 50932 6412
rect 50652 5182 50654 5234
rect 50706 5182 50708 5234
rect 50652 4900 50708 5182
rect 50652 4834 50708 4844
rect 50652 4676 50708 4686
rect 50652 4562 50708 4620
rect 50652 4510 50654 4562
rect 50706 4510 50708 4562
rect 50652 4498 50708 4510
rect 49868 4398 49870 4450
rect 49922 4398 49924 4450
rect 49868 4386 49924 4398
rect 49196 4286 49198 4338
rect 49250 4286 49252 4338
rect 49196 4274 49252 4286
rect 49512 3948 49776 3958
rect 49568 3892 49616 3948
rect 49672 3892 49720 3948
rect 49512 3882 49776 3892
rect 45836 3332 46004 3388
rect 47404 3378 47460 3388
rect 47964 3444 48020 3482
rect 48188 3444 48244 3454
rect 47964 3442 48244 3444
rect 47964 3390 47966 3442
rect 48018 3390 48190 3442
rect 48242 3390 48244 3442
rect 47964 3388 48244 3390
rect 45388 2996 45444 3332
rect 45388 2930 45444 2940
rect 45948 2772 46004 3332
rect 45948 2706 46004 2716
rect 47964 800 48020 3388
rect 48188 3378 48244 3388
rect 48524 3444 48580 3482
rect 48524 3378 48580 3388
rect 51212 3444 51268 21532
rect 51324 21586 51380 21644
rect 51324 21534 51326 21586
rect 51378 21534 51380 21586
rect 51324 21522 51380 21534
rect 51548 21588 51604 30716
rect 51772 29652 51828 29662
rect 51660 29426 51716 29438
rect 51660 29374 51662 29426
rect 51714 29374 51716 29426
rect 51660 26852 51716 29374
rect 51772 28980 51828 29596
rect 51884 29650 51940 31276
rect 51996 31108 52052 31118
rect 52108 31108 52164 32396
rect 52332 32386 52388 32396
rect 51996 31106 52164 31108
rect 51996 31054 51998 31106
rect 52050 31054 52164 31106
rect 51996 31052 52164 31054
rect 51996 31042 52052 31052
rect 52220 30994 52276 31006
rect 52220 30942 52222 30994
rect 52274 30942 52276 30994
rect 52220 29988 52276 30942
rect 52220 29922 52276 29932
rect 51884 29598 51886 29650
rect 51938 29598 51940 29650
rect 51884 29586 51940 29598
rect 51772 26908 51828 28924
rect 51996 29426 52052 29438
rect 51996 29374 51998 29426
rect 52050 29374 52052 29426
rect 51996 28418 52052 29374
rect 52220 29426 52276 29438
rect 52220 29374 52222 29426
rect 52274 29374 52276 29426
rect 51996 28366 51998 28418
rect 52050 28366 52052 28418
rect 51996 28354 52052 28366
rect 52108 28420 52164 28430
rect 52108 27858 52164 28364
rect 52220 28308 52276 29374
rect 52220 28242 52276 28252
rect 52108 27806 52110 27858
rect 52162 27806 52164 27858
rect 52108 27794 52164 27806
rect 51884 27748 51940 27758
rect 51884 27654 51940 27692
rect 51772 26852 51940 26908
rect 51660 26786 51716 26796
rect 51772 25284 51828 25294
rect 51660 24836 51716 24846
rect 51660 24722 51716 24780
rect 51660 24670 51662 24722
rect 51714 24670 51716 24722
rect 51660 23828 51716 24670
rect 51660 23762 51716 23772
rect 51660 23380 51716 23390
rect 51660 23286 51716 23324
rect 51660 23156 51716 23166
rect 51772 23156 51828 25228
rect 51716 23100 51828 23156
rect 51660 23090 51716 23100
rect 51660 22146 51716 22158
rect 51660 22094 51662 22146
rect 51714 22094 51716 22146
rect 51660 21924 51716 22094
rect 51660 21858 51716 21868
rect 51884 21812 51940 26852
rect 52108 26292 52164 26302
rect 51996 23828 52052 23838
rect 51996 23378 52052 23772
rect 51996 23326 51998 23378
rect 52050 23326 52052 23378
rect 51996 22036 52052 23326
rect 51996 21970 52052 21980
rect 51996 21812 52052 21822
rect 51884 21810 52052 21812
rect 51884 21758 51998 21810
rect 52050 21758 52052 21810
rect 51884 21756 52052 21758
rect 51996 21746 52052 21756
rect 51772 21700 51828 21738
rect 51772 21634 51828 21644
rect 51548 21522 51604 21532
rect 51884 21588 51940 21598
rect 51772 20692 51828 20702
rect 51772 20598 51828 20636
rect 51884 20690 51940 21532
rect 52108 20804 52164 26236
rect 52444 24948 52500 36652
rect 52556 27412 52612 37100
rect 53340 36708 53396 39200
rect 53340 36642 53396 36652
rect 53676 36482 53732 36494
rect 55020 36484 55076 36494
rect 53676 36430 53678 36482
rect 53730 36430 53732 36482
rect 53116 35140 53172 35150
rect 53116 34916 53172 35084
rect 53116 34850 53172 34860
rect 53564 34804 53620 34814
rect 53452 34748 53564 34804
rect 53228 33908 53284 33918
rect 52892 29988 52948 29998
rect 52948 29932 53060 29988
rect 52892 29922 52948 29932
rect 52780 29876 52836 29886
rect 52780 29316 52836 29820
rect 52892 29316 52948 29326
rect 52780 29314 52948 29316
rect 52780 29262 52894 29314
rect 52946 29262 52948 29314
rect 52780 29260 52948 29262
rect 52556 27346 52612 27356
rect 52668 28642 52724 28654
rect 52668 28590 52670 28642
rect 52722 28590 52724 28642
rect 52668 28308 52724 28590
rect 52556 26964 52612 26974
rect 52668 26908 52724 28252
rect 52780 28644 52836 29260
rect 52892 29250 52948 29260
rect 53004 28754 53060 29932
rect 53116 29652 53172 29662
rect 53116 29426 53172 29596
rect 53116 29374 53118 29426
rect 53170 29374 53172 29426
rect 53116 29362 53172 29374
rect 53228 29204 53284 33852
rect 53452 31890 53508 34748
rect 53564 34738 53620 34748
rect 53676 34468 53732 36430
rect 54236 36482 55076 36484
rect 54236 36430 55022 36482
rect 55074 36430 55076 36482
rect 54236 36428 55076 36430
rect 54236 35588 54292 36428
rect 55020 36418 55076 36428
rect 53900 35586 54292 35588
rect 53900 35534 54238 35586
rect 54290 35534 54292 35586
rect 53900 35532 54292 35534
rect 53900 35026 53956 35532
rect 54236 35522 54292 35532
rect 54572 35810 54628 35822
rect 54572 35758 54574 35810
rect 54626 35758 54628 35810
rect 53900 34974 53902 35026
rect 53954 34974 53956 35026
rect 53900 34962 53956 34974
rect 54348 35028 54404 35038
rect 54572 35028 54628 35758
rect 54908 35700 54964 35710
rect 54908 35588 54964 35644
rect 55356 35588 55412 35598
rect 54908 35586 55412 35588
rect 54908 35534 55358 35586
rect 55410 35534 55412 35586
rect 54908 35532 55412 35534
rect 54404 34972 54628 35028
rect 54348 34914 54404 34972
rect 54348 34862 54350 34914
rect 54402 34862 54404 34914
rect 54348 34850 54404 34862
rect 55132 34804 55188 34814
rect 55132 34710 55188 34748
rect 54012 34692 54068 34702
rect 54012 34690 54516 34692
rect 54012 34638 54014 34690
rect 54066 34638 54516 34690
rect 54012 34636 54516 34638
rect 54012 34626 54068 34636
rect 53676 34402 53732 34412
rect 54460 34356 54516 34636
rect 53676 34130 53732 34142
rect 53676 34078 53678 34130
rect 53730 34078 53732 34130
rect 53676 33348 53732 34078
rect 54124 34130 54180 34142
rect 54124 34078 54126 34130
rect 54178 34078 54180 34130
rect 54012 34020 54068 34030
rect 53676 33282 53732 33292
rect 53788 34018 54068 34020
rect 53788 33966 54014 34018
rect 54066 33966 54068 34018
rect 53788 33964 54068 33966
rect 53452 31838 53454 31890
rect 53506 31838 53508 31890
rect 53452 31826 53508 31838
rect 53564 31778 53620 31790
rect 53564 31726 53566 31778
rect 53618 31726 53620 31778
rect 53116 29148 53284 29204
rect 53340 31666 53396 31678
rect 53340 31614 53342 31666
rect 53394 31614 53396 31666
rect 53340 29204 53396 31614
rect 53564 30996 53620 31726
rect 53564 30930 53620 30940
rect 53788 30436 53844 33964
rect 54012 33954 54068 33964
rect 54124 34020 54180 34078
rect 54460 34130 54516 34300
rect 54460 34078 54462 34130
rect 54514 34078 54516 34130
rect 54460 34066 54516 34078
rect 54124 33954 54180 33964
rect 54348 33348 54404 33358
rect 54348 32452 54404 33292
rect 54908 33348 54964 33358
rect 54908 33254 54964 33292
rect 54460 33236 54516 33246
rect 54460 33234 54852 33236
rect 54460 33182 54462 33234
rect 54514 33182 54852 33234
rect 54460 33180 54852 33182
rect 54460 33170 54516 33180
rect 54460 32452 54516 32462
rect 54348 32450 54516 32452
rect 54348 32398 54462 32450
rect 54514 32398 54516 32450
rect 54348 32396 54516 32398
rect 54460 32386 54516 32396
rect 53900 31780 53956 31790
rect 53900 31686 53956 31724
rect 53788 30342 53844 30380
rect 53564 30210 53620 30222
rect 53564 30158 53566 30210
rect 53618 30158 53620 30210
rect 53452 29876 53508 29886
rect 53564 29876 53620 30158
rect 54124 29988 54180 29998
rect 54124 29986 54292 29988
rect 54124 29934 54126 29986
rect 54178 29934 54292 29986
rect 54124 29932 54292 29934
rect 54124 29922 54180 29932
rect 53508 29820 53620 29876
rect 53452 29810 53508 29820
rect 53452 29652 53508 29662
rect 53452 29650 53732 29652
rect 53452 29598 53454 29650
rect 53506 29598 53732 29650
rect 53452 29596 53732 29598
rect 53452 29586 53508 29596
rect 53676 29540 53732 29596
rect 53676 29484 54068 29540
rect 53676 29426 53732 29484
rect 53676 29374 53678 29426
rect 53730 29374 53732 29426
rect 53676 29362 53732 29374
rect 53900 29314 53956 29326
rect 53900 29262 53902 29314
rect 53954 29262 53956 29314
rect 53340 29148 53732 29204
rect 53116 28868 53172 29148
rect 53116 28812 53508 28868
rect 53004 28702 53006 28754
rect 53058 28702 53060 28754
rect 53004 28690 53060 28702
rect 52780 28196 52836 28588
rect 53228 28642 53284 28654
rect 53228 28590 53230 28642
rect 53282 28590 53284 28642
rect 52892 28420 52948 28430
rect 52892 28326 52948 28364
rect 53116 28418 53172 28430
rect 53116 28366 53118 28418
rect 53170 28366 53172 28418
rect 53004 28308 53060 28318
rect 52892 28196 52948 28206
rect 52780 28140 52892 28196
rect 52892 28130 52948 28140
rect 53004 26908 53060 28252
rect 53116 27748 53172 28366
rect 53116 27682 53172 27692
rect 52556 26852 52724 26908
rect 52780 26852 53060 26908
rect 53116 26852 53172 26862
rect 53228 26852 53284 28590
rect 53340 28196 53396 28206
rect 53340 27076 53396 28140
rect 53452 27298 53508 28812
rect 53564 28420 53620 28430
rect 53564 27634 53620 28364
rect 53676 28308 53732 29148
rect 53788 28532 53844 28542
rect 53788 28438 53844 28476
rect 53676 28242 53732 28252
rect 53676 27860 53732 27870
rect 53900 27860 53956 29262
rect 54012 28642 54068 29484
rect 54124 29426 54180 29438
rect 54124 29374 54126 29426
rect 54178 29374 54180 29426
rect 54124 29204 54180 29374
rect 54236 29428 54292 29932
rect 54684 29652 54740 29662
rect 54684 29558 54740 29596
rect 54796 29428 54852 33180
rect 54236 29426 54628 29428
rect 54236 29374 54238 29426
rect 54290 29374 54628 29426
rect 54236 29372 54628 29374
rect 54236 29362 54292 29372
rect 54180 29148 54404 29204
rect 54124 29138 54180 29148
rect 54012 28590 54014 28642
rect 54066 28590 54068 28642
rect 54012 28578 54068 28590
rect 54348 28642 54404 29148
rect 54348 28590 54350 28642
rect 54402 28590 54404 28642
rect 54348 28578 54404 28590
rect 54460 29092 54516 29102
rect 53676 27858 53956 27860
rect 53676 27806 53678 27858
rect 53730 27806 53956 27858
rect 53676 27804 53956 27806
rect 53676 27794 53732 27804
rect 53564 27582 53566 27634
rect 53618 27582 53620 27634
rect 53564 27570 53620 27582
rect 53564 27412 53620 27422
rect 53620 27356 53732 27412
rect 53564 27346 53620 27356
rect 53452 27246 53454 27298
rect 53506 27246 53508 27298
rect 53452 27234 53508 27246
rect 53564 27186 53620 27198
rect 53564 27134 53566 27186
rect 53618 27134 53620 27186
rect 53452 27076 53508 27086
rect 53340 27074 53508 27076
rect 53340 27022 53454 27074
rect 53506 27022 53508 27074
rect 53340 27020 53508 27022
rect 53452 27010 53508 27020
rect 52556 26290 52612 26852
rect 52780 26514 52836 26852
rect 52780 26462 52782 26514
rect 52834 26462 52836 26514
rect 52780 26450 52836 26462
rect 53172 26796 53284 26852
rect 53564 26852 53620 27134
rect 52556 26238 52558 26290
rect 52610 26238 52612 26290
rect 52556 26226 52612 26238
rect 52668 26292 52724 26302
rect 52668 26198 52724 26236
rect 52892 26290 52948 26302
rect 52892 26238 52894 26290
rect 52946 26238 52948 26290
rect 52892 25844 52948 26238
rect 53116 26290 53172 26796
rect 53564 26786 53620 26796
rect 53676 26908 53732 27356
rect 54348 27074 54404 27086
rect 54348 27022 54350 27074
rect 54402 27022 54404 27074
rect 53676 26852 54180 26908
rect 53116 26238 53118 26290
rect 53170 26238 53172 26290
rect 53116 26226 53172 26238
rect 52892 25284 52948 25788
rect 53228 25508 53284 25518
rect 53228 25414 53284 25452
rect 53676 25508 53732 26852
rect 54124 26514 54180 26852
rect 54124 26462 54126 26514
rect 54178 26462 54180 26514
rect 54124 26450 54180 26462
rect 53676 25414 53732 25452
rect 53788 25956 53844 25966
rect 52892 25218 52948 25228
rect 52668 24948 52724 24958
rect 53004 24948 53060 24958
rect 52220 24946 53060 24948
rect 52220 24894 52670 24946
rect 52722 24894 53006 24946
rect 53058 24894 53060 24946
rect 52220 24892 53060 24894
rect 52220 24050 52276 24892
rect 52668 24882 52724 24892
rect 52220 23998 52222 24050
rect 52274 23998 52276 24050
rect 52220 23986 52276 23998
rect 52780 24724 52836 24734
rect 52780 23380 52836 24668
rect 52892 24050 52948 24892
rect 53004 24882 53060 24892
rect 53788 24836 53844 25900
rect 54124 25394 54180 25406
rect 54124 25342 54126 25394
rect 54178 25342 54180 25394
rect 54124 25284 54180 25342
rect 54124 25218 54180 25228
rect 53788 24770 53844 24780
rect 53900 25060 53956 25070
rect 53900 24724 53956 25004
rect 53900 24630 53956 24668
rect 53564 24612 53620 24622
rect 53564 24610 53732 24612
rect 53564 24558 53566 24610
rect 53618 24558 53732 24610
rect 53564 24556 53732 24558
rect 53564 24546 53620 24556
rect 52892 23998 52894 24050
rect 52946 23998 52948 24050
rect 52892 23986 52948 23998
rect 53228 23940 53284 23950
rect 53228 23846 53284 23884
rect 53564 23714 53620 23726
rect 53564 23662 53566 23714
rect 53618 23662 53620 23714
rect 53116 23380 53172 23390
rect 53564 23380 53620 23662
rect 53676 23492 53732 24556
rect 54348 24276 54404 27022
rect 54012 24220 54404 24276
rect 54460 24276 54516 29036
rect 54572 28866 54628 29372
rect 54572 28814 54574 28866
rect 54626 28814 54628 28866
rect 54572 28802 54628 28814
rect 54796 28754 54852 29372
rect 54908 30436 54964 30446
rect 54908 29426 54964 30380
rect 54908 29374 54910 29426
rect 54962 29374 54964 29426
rect 54908 29362 54964 29374
rect 54796 28702 54798 28754
rect 54850 28702 54852 28754
rect 54796 28690 54852 28702
rect 54572 28532 54628 28542
rect 54572 28084 54628 28476
rect 54908 28532 54964 28542
rect 54908 28438 54964 28476
rect 55020 28530 55076 28542
rect 55020 28478 55022 28530
rect 55074 28478 55076 28530
rect 55020 28084 55076 28478
rect 54572 28082 55076 28084
rect 54572 28030 54574 28082
rect 54626 28030 55076 28082
rect 54572 28028 55076 28030
rect 54572 28018 54628 28028
rect 54908 27858 54964 28028
rect 55244 27972 55300 35532
rect 55356 35522 55412 35532
rect 55804 35252 55860 39200
rect 56028 36708 56084 36718
rect 56028 36614 56084 36652
rect 55804 35186 55860 35196
rect 57148 35700 57204 35710
rect 57148 35140 57204 35644
rect 58044 35586 58100 35598
rect 58044 35534 58046 35586
rect 58098 35534 58100 35586
rect 58044 35476 58100 35534
rect 58044 35410 58100 35420
rect 57148 35074 57204 35084
rect 58268 35140 58324 39200
rect 58268 35074 58324 35084
rect 58940 36482 58996 36494
rect 58940 36430 58942 36482
rect 58994 36430 58996 36482
rect 57260 35026 57316 35038
rect 57260 34974 57262 35026
rect 57314 34974 57316 35026
rect 57260 34916 57316 34974
rect 55580 34356 55636 34366
rect 55580 34262 55636 34300
rect 57260 34130 57316 34860
rect 57260 34078 57262 34130
rect 57314 34078 57316 34130
rect 57260 34066 57316 34078
rect 57596 34802 57652 34814
rect 57596 34750 57598 34802
rect 57650 34750 57652 34802
rect 55356 34020 55412 34030
rect 55356 33926 55412 33964
rect 55468 34018 55524 34030
rect 55468 33966 55470 34018
rect 55522 33966 55524 34018
rect 55468 33572 55524 33966
rect 57148 34018 57204 34030
rect 57148 33966 57150 34018
rect 57202 33966 57204 34018
rect 56924 33906 56980 33918
rect 56924 33854 56926 33906
rect 56978 33854 56980 33906
rect 56028 33572 56084 33582
rect 55468 33570 56084 33572
rect 55468 33518 56030 33570
rect 56082 33518 56084 33570
rect 55468 33516 56084 33518
rect 55356 33460 55412 33470
rect 55468 33460 55524 33516
rect 56028 33506 56084 33516
rect 55356 33458 55524 33460
rect 55356 33406 55358 33458
rect 55410 33406 55524 33458
rect 55356 33404 55524 33406
rect 55356 33394 55412 33404
rect 55804 33348 55860 33358
rect 55804 33254 55860 33292
rect 56364 33348 56420 33358
rect 56364 33254 56420 33292
rect 56700 30884 56756 30894
rect 55468 30660 55524 30670
rect 55132 27916 55300 27972
rect 55356 29538 55412 29550
rect 55356 29486 55358 29538
rect 55410 29486 55412 29538
rect 54908 27806 54910 27858
rect 54962 27806 54964 27858
rect 54908 27794 54964 27806
rect 55020 27860 55076 27870
rect 55020 27746 55076 27804
rect 55020 27694 55022 27746
rect 55074 27694 55076 27746
rect 55020 27682 55076 27694
rect 55132 26908 55188 27916
rect 55244 27748 55300 27758
rect 55356 27748 55412 29486
rect 55300 27692 55412 27748
rect 55244 27654 55300 27692
rect 55132 26852 55300 26908
rect 54572 25508 54628 25546
rect 54572 25442 54628 25452
rect 54796 25394 54852 25406
rect 54796 25342 54798 25394
rect 54850 25342 54852 25394
rect 54796 24724 54852 25342
rect 55132 25284 55188 25294
rect 54796 24658 54852 24668
rect 55020 25228 55132 25284
rect 53676 23436 53844 23492
rect 52780 23378 53060 23380
rect 52780 23326 52782 23378
rect 52834 23326 53060 23378
rect 52780 23324 53060 23326
rect 52780 23314 52836 23324
rect 53004 23266 53060 23324
rect 53116 23378 53620 23380
rect 53116 23326 53118 23378
rect 53170 23326 53620 23378
rect 53116 23324 53620 23326
rect 53116 23314 53172 23324
rect 53004 23214 53006 23266
rect 53058 23214 53060 23266
rect 53004 23202 53060 23214
rect 53564 23156 53620 23324
rect 53564 23090 53620 23100
rect 53788 23044 53844 23436
rect 53900 23044 53956 23054
rect 53788 22988 53900 23044
rect 53900 22978 53956 22988
rect 53564 22932 53620 22942
rect 52220 22146 52276 22158
rect 52220 22094 52222 22146
rect 52274 22094 52276 22146
rect 52220 21586 52276 22094
rect 52892 21924 52948 21934
rect 52332 21812 52388 21822
rect 52332 21718 52388 21756
rect 52220 21534 52222 21586
rect 52274 21534 52276 21586
rect 52220 20916 52276 21534
rect 52332 21476 52388 21486
rect 52332 21474 52724 21476
rect 52332 21422 52334 21474
rect 52386 21422 52724 21474
rect 52332 21420 52724 21422
rect 52332 21410 52388 21420
rect 52220 20860 52388 20916
rect 52108 20748 52276 20804
rect 51884 20638 51886 20690
rect 51938 20638 51940 20690
rect 51884 20468 51940 20638
rect 52108 20580 52164 20590
rect 52108 20486 52164 20524
rect 51436 20412 51940 20468
rect 51436 19346 51492 20412
rect 51436 19294 51438 19346
rect 51490 19294 51492 19346
rect 51436 19282 51492 19294
rect 51884 20242 51940 20254
rect 51884 20190 51886 20242
rect 51938 20190 51940 20242
rect 51324 17556 51380 17566
rect 51324 17462 51380 17500
rect 51548 16212 51604 16222
rect 51548 16118 51604 16156
rect 51436 15988 51492 15998
rect 51436 15540 51492 15932
rect 51436 15314 51492 15484
rect 51436 15262 51438 15314
rect 51490 15262 51492 15314
rect 51436 15250 51492 15262
rect 51772 15202 51828 15214
rect 51772 15150 51774 15202
rect 51826 15150 51828 15202
rect 51660 15092 51716 15102
rect 51660 14642 51716 15036
rect 51660 14590 51662 14642
rect 51714 14590 51716 14642
rect 51660 14578 51716 14590
rect 51660 13748 51716 13758
rect 51660 13076 51716 13692
rect 51660 13010 51716 13020
rect 51772 13636 51828 15150
rect 51548 12964 51604 12974
rect 51436 12962 51604 12964
rect 51436 12910 51550 12962
rect 51602 12910 51604 12962
rect 51436 12908 51604 12910
rect 51324 10052 51380 10062
rect 51324 9714 51380 9996
rect 51436 9940 51492 12908
rect 51548 12898 51604 12908
rect 51772 12178 51828 13580
rect 51884 13188 51940 20190
rect 51996 18228 52052 18238
rect 51996 13524 52052 18172
rect 52220 16548 52276 20748
rect 52220 16482 52276 16492
rect 52220 15988 52276 15998
rect 52220 15894 52276 15932
rect 52332 15148 52388 20860
rect 52668 20802 52724 21420
rect 52668 20750 52670 20802
rect 52722 20750 52724 20802
rect 52668 20738 52724 20750
rect 52780 20580 52836 20590
rect 52780 20486 52836 20524
rect 52668 20356 52724 20366
rect 52668 17332 52724 20300
rect 52892 20018 52948 21868
rect 52892 19966 52894 20018
rect 52946 19966 52948 20018
rect 52892 19954 52948 19966
rect 53004 20578 53060 20590
rect 53452 20580 53508 20590
rect 53004 20526 53006 20578
rect 53058 20526 53060 20578
rect 52780 19908 52836 19918
rect 52780 19234 52836 19852
rect 52780 19182 52782 19234
rect 52834 19182 52836 19234
rect 52780 19170 52836 19182
rect 53004 19124 53060 20526
rect 53340 20578 53508 20580
rect 53340 20526 53454 20578
rect 53506 20526 53508 20578
rect 53340 20524 53508 20526
rect 53228 19908 53284 19918
rect 53060 19068 53172 19124
rect 53004 19058 53060 19068
rect 53116 17890 53172 19068
rect 53116 17838 53118 17890
rect 53170 17838 53172 17890
rect 53116 17826 53172 17838
rect 53228 17780 53284 19852
rect 53340 19348 53396 20524
rect 53452 20514 53508 20524
rect 53452 19348 53508 19358
rect 53340 19346 53508 19348
rect 53340 19294 53454 19346
rect 53506 19294 53508 19346
rect 53340 19292 53508 19294
rect 53452 19282 53508 19292
rect 53452 18338 53508 18350
rect 53452 18286 53454 18338
rect 53506 18286 53508 18338
rect 53452 18228 53508 18286
rect 53452 18162 53508 18172
rect 53228 17724 53396 17780
rect 52780 17556 52836 17566
rect 52780 17462 52836 17500
rect 52668 17276 53172 17332
rect 52892 16772 52948 16782
rect 52892 16678 52948 16716
rect 52780 16548 52836 16558
rect 52220 15092 52388 15148
rect 52556 16100 52612 16110
rect 52556 15538 52612 16044
rect 52556 15486 52558 15538
rect 52610 15486 52612 15538
rect 51996 13458 52052 13468
rect 52108 14532 52164 14542
rect 52108 13412 52164 14476
rect 52108 13346 52164 13356
rect 51884 13132 52164 13188
rect 51772 12126 51774 12178
rect 51826 12126 51828 12178
rect 51772 12114 51828 12126
rect 52108 11732 52164 13132
rect 52108 11666 52164 11676
rect 51548 11396 51604 11406
rect 51548 10052 51604 11340
rect 52108 11284 52164 11294
rect 52108 11190 52164 11228
rect 51772 11172 51828 11182
rect 51660 11170 51828 11172
rect 51660 11118 51774 11170
rect 51826 11118 51828 11170
rect 51660 11116 51828 11118
rect 51660 10722 51716 11116
rect 51772 11106 51828 11116
rect 51660 10670 51662 10722
rect 51714 10670 51716 10722
rect 51660 10658 51716 10670
rect 51660 10052 51716 10062
rect 51548 10050 51716 10052
rect 51548 9998 51662 10050
rect 51714 9998 51716 10050
rect 51548 9996 51716 9998
rect 51660 9986 51716 9996
rect 51436 9874 51492 9884
rect 51324 9662 51326 9714
rect 51378 9662 51380 9714
rect 51324 9650 51380 9662
rect 51996 9604 52052 9614
rect 51996 9510 52052 9548
rect 51772 8372 51828 8382
rect 51772 6916 51828 8316
rect 52220 7812 52276 15092
rect 52556 13748 52612 15486
rect 52780 14868 52836 16492
rect 53004 15202 53060 15214
rect 53004 15150 53006 15202
rect 53058 15150 53060 15202
rect 52780 14802 52836 14812
rect 52892 14980 52948 14990
rect 52892 14530 52948 14924
rect 52892 14478 52894 14530
rect 52946 14478 52948 14530
rect 52892 14466 52948 14478
rect 52780 14420 52836 14430
rect 52780 13972 52836 14364
rect 53004 14196 53060 15150
rect 53004 14130 53060 14140
rect 52892 13972 52948 13982
rect 52780 13970 52948 13972
rect 52780 13918 52894 13970
rect 52946 13918 52948 13970
rect 52780 13916 52948 13918
rect 52556 13682 52612 13692
rect 52444 13522 52500 13534
rect 52444 13470 52446 13522
rect 52498 13470 52500 13522
rect 52444 12964 52500 13470
rect 52444 12898 52500 12908
rect 52892 12404 52948 13916
rect 52892 12338 52948 12348
rect 52332 12180 52388 12190
rect 52332 12086 52388 12124
rect 53116 11620 53172 17276
rect 53340 17106 53396 17724
rect 53340 17054 53342 17106
rect 53394 17054 53396 17106
rect 53340 16996 53396 17054
rect 53340 16548 53396 16940
rect 53340 16482 53396 16492
rect 53004 11564 53172 11620
rect 53228 14644 53284 14654
rect 52780 11284 52836 11294
rect 52780 11190 52836 11228
rect 53004 10724 53060 11564
rect 53116 11396 53172 11406
rect 53116 11302 53172 11340
rect 52780 10668 53060 10724
rect 52668 9604 52724 9614
rect 52556 9602 52724 9604
rect 52556 9550 52670 9602
rect 52722 9550 52724 9602
rect 52556 9548 52724 9550
rect 52556 9154 52612 9548
rect 52668 9538 52724 9548
rect 52556 9102 52558 9154
rect 52610 9102 52612 9154
rect 52556 9090 52612 9102
rect 52220 7746 52276 7756
rect 52444 7476 52500 7486
rect 52444 7474 52724 7476
rect 52444 7422 52446 7474
rect 52498 7422 52724 7474
rect 52444 7420 52724 7422
rect 52444 7410 52500 7420
rect 51772 6130 51828 6860
rect 51772 6078 51774 6130
rect 51826 6078 51828 6130
rect 51772 6066 51828 6078
rect 52668 5908 52724 7420
rect 52668 5012 52724 5852
rect 52332 5010 52724 5012
rect 52332 4958 52670 5010
rect 52722 4958 52724 5010
rect 52332 4956 52724 4958
rect 52332 4338 52388 4956
rect 52668 4946 52724 4956
rect 52332 4286 52334 4338
rect 52386 4286 52388 4338
rect 52332 4274 52388 4286
rect 51212 3378 51268 3388
rect 51996 3444 52052 3482
rect 52220 3444 52276 3454
rect 51996 3442 52276 3444
rect 51996 3390 51998 3442
rect 52050 3390 52222 3442
rect 52274 3390 52276 3442
rect 51996 3388 52276 3390
rect 51996 800 52052 3388
rect 52220 3378 52276 3388
rect 52556 3444 52612 3454
rect 52780 3444 52836 10668
rect 52892 9826 52948 9838
rect 52892 9774 52894 9826
rect 52946 9774 52948 9826
rect 52892 9604 52948 9774
rect 53228 9828 53284 14588
rect 53340 13748 53396 13758
rect 53340 13654 53396 13692
rect 53564 13188 53620 22876
rect 53676 20802 53732 20814
rect 53676 20750 53678 20802
rect 53730 20750 53732 20802
rect 53676 18676 53732 20750
rect 53676 18620 53844 18676
rect 53788 18450 53844 18620
rect 53788 18398 53790 18450
rect 53842 18398 53844 18450
rect 53788 18386 53844 18398
rect 54012 18116 54068 24220
rect 54460 24210 54516 24220
rect 54684 24498 54740 24510
rect 54684 24446 54686 24498
rect 54738 24446 54740 24498
rect 54124 24052 54180 24062
rect 54124 23958 54180 23996
rect 54460 23940 54516 23950
rect 54348 23884 54460 23940
rect 54236 23156 54292 23166
rect 54236 23062 54292 23100
rect 54124 23042 54180 23054
rect 54124 22990 54126 23042
rect 54178 22990 54180 23042
rect 54124 19348 54180 22990
rect 54348 22370 54404 23884
rect 54460 23846 54516 23884
rect 54572 23714 54628 23726
rect 54572 23662 54574 23714
rect 54626 23662 54628 23714
rect 54460 23492 54516 23502
rect 54460 22484 54516 23436
rect 54572 22932 54628 23662
rect 54572 22866 54628 22876
rect 54460 22418 54516 22428
rect 54684 22484 54740 24446
rect 54684 22418 54740 22428
rect 54796 24388 54852 24398
rect 54348 22318 54350 22370
rect 54402 22318 54404 22370
rect 54348 22306 54404 22318
rect 54460 22148 54516 22158
rect 54460 22146 54740 22148
rect 54460 22094 54462 22146
rect 54514 22094 54740 22146
rect 54460 22092 54740 22094
rect 54460 22082 54516 22092
rect 54348 20020 54404 20030
rect 54348 19926 54404 19964
rect 54124 19292 54404 19348
rect 54124 19124 54180 19134
rect 54124 18450 54180 19068
rect 54124 18398 54126 18450
rect 54178 18398 54180 18450
rect 54124 18386 54180 18398
rect 54236 18564 54292 18574
rect 54012 18050 54068 18060
rect 53676 17780 53732 17790
rect 53676 17666 53732 17724
rect 53676 17614 53678 17666
rect 53730 17614 53732 17666
rect 53676 17602 53732 17614
rect 53900 17554 53956 17566
rect 53900 17502 53902 17554
rect 53954 17502 53956 17554
rect 53676 17332 53732 17342
rect 53676 16098 53732 17276
rect 53900 16772 53956 17502
rect 53900 16706 53956 16716
rect 53676 16046 53678 16098
rect 53730 16046 53732 16098
rect 53676 16034 53732 16046
rect 54012 16098 54068 16110
rect 54012 16046 54014 16098
rect 54066 16046 54068 16098
rect 54012 15988 54068 16046
rect 54012 15922 54068 15932
rect 54236 14644 54292 18508
rect 54348 17108 54404 19292
rect 54684 18676 54740 22092
rect 54796 20244 54852 24332
rect 55020 23828 55076 25228
rect 55132 25218 55188 25228
rect 55132 25060 55188 25070
rect 55132 24946 55188 25004
rect 55132 24894 55134 24946
rect 55186 24894 55188 24946
rect 55132 24882 55188 24894
rect 54908 23826 55076 23828
rect 54908 23774 55022 23826
rect 55074 23774 55076 23826
rect 54908 23772 55076 23774
rect 54908 22258 54964 23772
rect 55020 23762 55076 23772
rect 54908 22206 54910 22258
rect 54962 22206 54964 22258
rect 54908 22194 54964 22206
rect 54796 20178 54852 20188
rect 55132 20578 55188 20590
rect 55132 20526 55134 20578
rect 55186 20526 55188 20578
rect 55020 20130 55076 20142
rect 55020 20078 55022 20130
rect 55074 20078 55076 20130
rect 55020 19572 55076 20078
rect 55020 19506 55076 19516
rect 55132 18900 55188 20526
rect 55020 18844 55188 18900
rect 54684 18620 54852 18676
rect 54684 18450 54740 18462
rect 54684 18398 54686 18450
rect 54738 18398 54740 18450
rect 54684 18228 54740 18398
rect 54684 18162 54740 18172
rect 54460 17780 54516 17790
rect 54460 17686 54516 17724
rect 54684 17108 54740 17118
rect 54348 17052 54516 17108
rect 54348 16884 54404 16894
rect 54348 16790 54404 16828
rect 54348 16100 54404 16110
rect 54348 16006 54404 16044
rect 54460 15988 54516 17052
rect 54684 17014 54740 17052
rect 54684 16772 54740 16782
rect 54684 16098 54740 16716
rect 54684 16046 54686 16098
rect 54738 16046 54740 16098
rect 54684 16034 54740 16046
rect 54460 15540 54516 15932
rect 54796 15764 54852 18620
rect 54908 18564 54964 18574
rect 54908 18470 54964 18508
rect 55020 18340 55076 18844
rect 54460 15474 54516 15484
rect 54684 15708 54852 15764
rect 54908 18284 55076 18340
rect 55132 18676 55188 18686
rect 54908 15764 54964 18284
rect 55020 17892 55076 17902
rect 55020 16996 55076 17836
rect 55020 16930 55076 16940
rect 55132 16882 55188 18620
rect 55132 16830 55134 16882
rect 55186 16830 55188 16882
rect 55132 16818 55188 16830
rect 54012 14588 54292 14644
rect 54348 14644 54404 14654
rect 53788 14418 53844 14430
rect 53788 14366 53790 14418
rect 53842 14366 53844 14418
rect 53788 13860 53844 14366
rect 53788 13794 53844 13804
rect 53564 13122 53620 13132
rect 53452 12964 53508 12974
rect 53452 12290 53508 12908
rect 53564 12404 53620 12414
rect 54012 12404 54068 14588
rect 54348 14550 54404 14588
rect 54684 14644 54740 15708
rect 54908 15698 54964 15708
rect 54796 15540 54852 15550
rect 55132 15540 55188 15550
rect 54852 15538 55188 15540
rect 54852 15486 55134 15538
rect 55186 15486 55188 15538
rect 54852 15484 55188 15486
rect 54796 15446 54852 15484
rect 55132 15474 55188 15484
rect 55244 15148 55300 26852
rect 55468 26404 55524 30604
rect 56700 30324 56756 30828
rect 56700 30210 56756 30268
rect 56700 30158 56702 30210
rect 56754 30158 56756 30210
rect 56700 30146 56756 30158
rect 55580 29428 55636 29438
rect 55580 29334 55636 29372
rect 55916 28642 55972 28654
rect 55916 28590 55918 28642
rect 55970 28590 55972 28642
rect 55692 28530 55748 28542
rect 55692 28478 55694 28530
rect 55746 28478 55748 28530
rect 55692 27860 55748 28478
rect 55916 28532 55972 28590
rect 55916 28466 55972 28476
rect 55692 27794 55748 27804
rect 56252 28418 56308 28430
rect 56252 28366 56254 28418
rect 56306 28366 56308 28418
rect 56252 27860 56308 28366
rect 56252 27794 56308 27804
rect 56700 28418 56756 28430
rect 56700 28366 56702 28418
rect 56754 28366 56756 28418
rect 56700 27746 56756 28366
rect 56700 27694 56702 27746
rect 56754 27694 56756 27746
rect 56700 26964 56756 27694
rect 56700 26516 56756 26908
rect 56700 26450 56756 26460
rect 55468 26338 55524 26348
rect 55580 26292 55636 26302
rect 55580 25618 55636 26236
rect 55580 25566 55582 25618
rect 55634 25566 55636 25618
rect 55580 25554 55636 25566
rect 56924 25844 56980 33854
rect 57148 33570 57204 33966
rect 57148 33518 57150 33570
rect 57202 33518 57204 33570
rect 57148 33506 57204 33518
rect 57596 33460 57652 34750
rect 57932 34804 57988 34814
rect 57932 34710 57988 34748
rect 58940 34580 58996 36430
rect 60620 36370 60676 36382
rect 60620 36318 60622 36370
rect 60674 36318 60676 36370
rect 59172 36092 59436 36102
rect 59228 36036 59276 36092
rect 59332 36036 59380 36092
rect 59172 36026 59436 36036
rect 60284 35586 60340 35598
rect 60284 35534 60286 35586
rect 60338 35534 60340 35586
rect 60284 34804 60340 35534
rect 60620 35252 60676 36318
rect 60620 35186 60676 35196
rect 60284 34738 60340 34748
rect 60620 34916 60676 34926
rect 58940 34514 58996 34524
rect 59172 34524 59436 34534
rect 58828 34468 58884 34478
rect 59228 34468 59276 34524
rect 59332 34468 59380 34524
rect 59172 34458 59436 34468
rect 58156 34356 58212 34366
rect 57596 33394 57652 33404
rect 57820 34354 58212 34356
rect 57820 34302 58158 34354
rect 58210 34302 58212 34354
rect 57820 34300 58212 34302
rect 57148 33236 57204 33246
rect 57148 33012 57204 33180
rect 57260 33234 57316 33246
rect 57260 33182 57262 33234
rect 57314 33182 57316 33234
rect 57260 33124 57316 33182
rect 57596 33124 57652 33134
rect 57260 33122 57652 33124
rect 57260 33070 57598 33122
rect 57650 33070 57652 33122
rect 57260 33068 57652 33070
rect 57148 32956 57428 33012
rect 57372 32788 57428 32956
rect 57372 32694 57428 32732
rect 57596 32452 57652 33068
rect 57596 32386 57652 32396
rect 57820 31556 57876 34300
rect 58156 34290 58212 34300
rect 58828 34242 58884 34412
rect 58828 34190 58830 34242
rect 58882 34190 58884 34242
rect 58044 34132 58100 34142
rect 58100 34076 58212 34132
rect 58044 34038 58100 34076
rect 58044 33348 58100 33358
rect 58044 33254 58100 33292
rect 58156 33346 58212 34076
rect 58828 34020 58884 34190
rect 60060 34244 60116 34254
rect 60620 34244 60676 34860
rect 60732 34580 60788 39200
rect 62636 36484 62692 36494
rect 62636 36390 62692 36428
rect 63196 35924 63252 39200
rect 63196 35858 63252 35868
rect 64092 36706 64148 36718
rect 64092 36654 64094 36706
rect 64146 36654 64148 36706
rect 63868 35812 63924 35822
rect 63868 35718 63924 35756
rect 60956 35698 61012 35710
rect 60956 35646 60958 35698
rect 61010 35646 61012 35698
rect 60956 34916 61012 35646
rect 60956 34850 61012 34860
rect 61068 35476 61124 35486
rect 60732 34524 60900 34580
rect 60732 34244 60788 34254
rect 60620 34188 60732 34244
rect 60060 34150 60116 34188
rect 58828 33572 58884 33964
rect 58156 33294 58158 33346
rect 58210 33294 58212 33346
rect 58156 33282 58212 33294
rect 58380 33516 58828 33572
rect 58380 33346 58436 33516
rect 58828 33478 58884 33516
rect 59052 34130 59108 34142
rect 59052 34078 59054 34130
rect 59106 34078 59108 34130
rect 58380 33294 58382 33346
rect 58434 33294 58436 33346
rect 58380 33282 58436 33294
rect 59052 33348 59108 34078
rect 60396 34130 60452 34142
rect 60396 34078 60398 34130
rect 60450 34078 60452 34130
rect 59052 33254 59108 33292
rect 59276 33572 59332 33582
rect 59276 33346 59332 33516
rect 59276 33294 59278 33346
rect 59330 33294 59332 33346
rect 59276 33282 59332 33294
rect 59948 33236 60004 33246
rect 59948 33234 60228 33236
rect 59948 33182 59950 33234
rect 60002 33182 60228 33234
rect 59948 33180 60228 33182
rect 59948 33170 60004 33180
rect 59172 32956 59436 32966
rect 59228 32900 59276 32956
rect 59332 32900 59380 32956
rect 59172 32890 59436 32900
rect 58156 32788 58212 32798
rect 58156 32562 58212 32732
rect 59500 32788 59556 32798
rect 59836 32788 59892 32798
rect 59556 32732 59668 32788
rect 59500 32722 59556 32732
rect 58156 32510 58158 32562
rect 58210 32510 58212 32562
rect 58156 32498 58212 32510
rect 57596 31500 57876 31556
rect 58492 32452 58548 32462
rect 57596 30884 57652 31500
rect 57820 30994 57876 31006
rect 57820 30942 57822 30994
rect 57874 30942 57876 30994
rect 57820 30884 57876 30942
rect 57596 30882 57764 30884
rect 57596 30830 57598 30882
rect 57650 30830 57764 30882
rect 57596 30828 57764 30830
rect 57820 30828 58324 30884
rect 57596 30818 57652 30828
rect 57372 30770 57428 30782
rect 57372 30718 57374 30770
rect 57426 30718 57428 30770
rect 57372 30212 57428 30718
rect 57708 30772 57764 30828
rect 57708 30716 58100 30772
rect 57148 29986 57204 29998
rect 57148 29934 57150 29986
rect 57202 29934 57204 29986
rect 57148 29764 57204 29934
rect 57148 29698 57204 29708
rect 57148 28980 57204 28990
rect 57036 28418 57092 28430
rect 57036 28366 57038 28418
rect 57090 28366 57092 28418
rect 57036 27972 57092 28366
rect 57036 27906 57092 27916
rect 57148 26964 57204 28924
rect 57148 26898 57204 26908
rect 57148 26740 57204 26750
rect 57036 26684 57148 26740
rect 57036 26514 57092 26684
rect 57148 26674 57204 26684
rect 57036 26462 57038 26514
rect 57090 26462 57092 26514
rect 57036 26450 57092 26462
rect 57260 26402 57316 26414
rect 57260 26350 57262 26402
rect 57314 26350 57316 26402
rect 57260 26068 57316 26350
rect 57372 26292 57428 30156
rect 57820 30098 57876 30110
rect 57820 30046 57822 30098
rect 57874 30046 57876 30098
rect 57820 29764 57876 30046
rect 57484 29204 57540 29214
rect 57484 28866 57540 29148
rect 57484 28814 57486 28866
rect 57538 28814 57540 28866
rect 57484 28802 57540 28814
rect 57596 28530 57652 28542
rect 57596 28478 57598 28530
rect 57650 28478 57652 28530
rect 57484 28418 57540 28430
rect 57484 28366 57486 28418
rect 57538 28366 57540 28418
rect 57484 27972 57540 28366
rect 57596 28420 57652 28478
rect 57596 28354 57652 28364
rect 57484 27906 57540 27916
rect 57372 26290 57540 26292
rect 57372 26238 57374 26290
rect 57426 26238 57540 26290
rect 57372 26236 57540 26238
rect 57372 26226 57428 26236
rect 57260 26012 57428 26068
rect 56252 25506 56308 25518
rect 56252 25454 56254 25506
rect 56306 25454 56308 25506
rect 56252 24836 56308 25454
rect 56924 25506 56980 25788
rect 56924 25454 56926 25506
rect 56978 25454 56980 25506
rect 56924 25442 56980 25454
rect 57148 25394 57204 25406
rect 57148 25342 57150 25394
rect 57202 25342 57204 25394
rect 57148 24836 57204 25342
rect 56252 24770 56308 24780
rect 57036 24780 57204 24836
rect 57372 25284 57428 26012
rect 55356 24724 55412 24734
rect 55356 23268 55412 24668
rect 55468 24722 55524 24734
rect 55468 24670 55470 24722
rect 55522 24670 55524 24722
rect 55468 23940 55524 24670
rect 56588 24724 56644 24734
rect 56588 24630 56644 24668
rect 56028 24612 56084 24622
rect 56028 24610 56420 24612
rect 56028 24558 56030 24610
rect 56082 24558 56420 24610
rect 56028 24556 56420 24558
rect 56028 24546 56084 24556
rect 56364 24388 56420 24556
rect 56252 24052 56308 24062
rect 56252 23958 56308 23996
rect 55468 23874 55524 23884
rect 55468 23268 55524 23278
rect 55356 23266 55524 23268
rect 55356 23214 55470 23266
rect 55522 23214 55524 23266
rect 55356 23212 55524 23214
rect 55356 20692 55412 23212
rect 55468 23202 55524 23212
rect 56028 23154 56084 23166
rect 56028 23102 56030 23154
rect 56082 23102 56084 23154
rect 56028 23044 56084 23102
rect 56028 22978 56084 22988
rect 56140 22484 56196 22494
rect 56140 22390 56196 22428
rect 56364 22036 56420 24332
rect 57036 24052 57092 24780
rect 57260 24724 57316 24734
rect 57148 24668 57260 24724
rect 57148 24610 57204 24668
rect 57260 24658 57316 24668
rect 57148 24558 57150 24610
rect 57202 24558 57204 24610
rect 57148 24546 57204 24558
rect 57372 24276 57428 25228
rect 57036 23986 57092 23996
rect 57148 24220 57428 24276
rect 57148 23266 57204 24220
rect 57484 23940 57540 26236
rect 57820 25284 57876 29708
rect 58044 29426 58100 30716
rect 58268 30770 58324 30828
rect 58268 30718 58270 30770
rect 58322 30718 58324 30770
rect 58156 30324 58212 30334
rect 58156 30210 58212 30268
rect 58156 30158 58158 30210
rect 58210 30158 58212 30210
rect 58156 30146 58212 30158
rect 58044 29374 58046 29426
rect 58098 29374 58100 29426
rect 58044 29362 58100 29374
rect 58156 29428 58212 29438
rect 58044 28756 58100 28766
rect 58156 28756 58212 29372
rect 58268 29426 58324 30718
rect 58492 30770 58548 32396
rect 59388 32452 59444 32462
rect 59388 32450 59556 32452
rect 59388 32398 59390 32450
rect 59442 32398 59556 32450
rect 59388 32396 59556 32398
rect 59388 32386 59444 32396
rect 58716 31554 58772 31566
rect 58716 31502 58718 31554
rect 58770 31502 58772 31554
rect 58716 30996 58772 31502
rect 59172 31388 59436 31398
rect 59228 31332 59276 31388
rect 59332 31332 59380 31388
rect 59172 31322 59436 31332
rect 58492 30718 58494 30770
rect 58546 30718 58548 30770
rect 58492 30706 58548 30718
rect 58604 30882 58660 30894
rect 58604 30830 58606 30882
rect 58658 30830 58660 30882
rect 58604 30660 58660 30830
rect 58604 30594 58660 30604
rect 58716 30324 58772 30940
rect 58716 30258 58772 30268
rect 59052 30994 59108 31006
rect 59052 30942 59054 30994
rect 59106 30942 59108 30994
rect 58940 30212 58996 30222
rect 58940 30118 58996 30156
rect 58828 30100 58884 30110
rect 58828 30006 58884 30044
rect 58268 29374 58270 29426
rect 58322 29374 58324 29426
rect 58268 29362 58324 29374
rect 59052 29988 59108 30942
rect 59388 30996 59444 31006
rect 59500 30996 59556 32396
rect 59612 32116 59668 32732
rect 59836 32694 59892 32732
rect 59948 32674 60004 32686
rect 59948 32622 59950 32674
rect 60002 32622 60004 32674
rect 59724 32340 59780 32350
rect 59724 32338 59892 32340
rect 59724 32286 59726 32338
rect 59778 32286 59892 32338
rect 59724 32284 59892 32286
rect 59724 32274 59780 32284
rect 59612 31892 59668 32060
rect 59724 31892 59780 31902
rect 59612 31890 59780 31892
rect 59612 31838 59726 31890
rect 59778 31838 59780 31890
rect 59612 31836 59780 31838
rect 59724 31826 59780 31836
rect 59388 30994 59556 30996
rect 59388 30942 59390 30994
rect 59442 30942 59556 30994
rect 59388 30940 59556 30942
rect 59388 30436 59444 30940
rect 59724 30882 59780 30894
rect 59724 30830 59726 30882
rect 59778 30830 59780 30882
rect 59500 30772 59556 30782
rect 59500 30770 59668 30772
rect 59500 30718 59502 30770
rect 59554 30718 59668 30770
rect 59500 30716 59668 30718
rect 59500 30706 59556 30716
rect 59500 30436 59556 30446
rect 59388 30380 59500 30436
rect 59500 30370 59556 30380
rect 59500 30212 59556 30222
rect 59500 29988 59556 30156
rect 59052 29932 59556 29988
rect 58044 28754 58212 28756
rect 58044 28702 58046 28754
rect 58098 28702 58212 28754
rect 58044 28700 58212 28702
rect 58268 29202 58324 29214
rect 58268 29150 58270 29202
rect 58322 29150 58324 29202
rect 58044 28690 58100 28700
rect 57932 28644 57988 28654
rect 57932 28550 57988 28588
rect 58268 28642 58324 29150
rect 59052 28868 59108 29932
rect 59172 29820 59436 29830
rect 59228 29764 59276 29820
rect 59332 29764 59380 29820
rect 59172 29754 59436 29764
rect 59052 28802 59108 28812
rect 59276 29540 59332 29550
rect 58268 28590 58270 28642
rect 58322 28590 58324 28642
rect 58268 28532 58324 28590
rect 58492 28756 58548 28766
rect 58492 28642 58548 28700
rect 58940 28754 58996 28766
rect 58940 28702 58942 28754
rect 58994 28702 58996 28754
rect 58492 28590 58494 28642
rect 58546 28590 58548 28642
rect 58492 28578 58548 28590
rect 58716 28644 58772 28654
rect 58772 28588 58884 28644
rect 58716 28550 58772 28588
rect 58268 28466 58324 28476
rect 58828 27972 58884 28588
rect 58940 28420 58996 28702
rect 59276 28644 59332 29484
rect 58940 28354 58996 28364
rect 59052 28532 59108 28542
rect 58828 27916 58996 27972
rect 58716 27860 58772 27870
rect 58716 27858 58884 27860
rect 58716 27806 58718 27858
rect 58770 27806 58884 27858
rect 58716 27804 58884 27806
rect 58716 27794 58772 27804
rect 58828 27298 58884 27804
rect 58828 27246 58830 27298
rect 58882 27246 58884 27298
rect 58828 27234 58884 27246
rect 58940 27186 58996 27916
rect 59052 27858 59108 28476
rect 59276 28530 59332 28588
rect 59276 28478 59278 28530
rect 59330 28478 59332 28530
rect 59276 28466 59332 28478
rect 59388 29426 59444 29438
rect 59612 29428 59668 30716
rect 59724 30660 59780 30830
rect 59836 30772 59892 32284
rect 59948 31780 60004 32622
rect 59948 31714 60004 31724
rect 60060 31668 60116 31678
rect 60060 31218 60116 31612
rect 60060 31166 60062 31218
rect 60114 31166 60116 31218
rect 60060 31154 60116 31166
rect 59948 30996 60004 31006
rect 59948 30902 60004 30940
rect 59836 30716 60116 30772
rect 59724 30594 59780 30604
rect 59836 30436 59892 30446
rect 59724 30100 59780 30110
rect 59724 29650 59780 30044
rect 59724 29598 59726 29650
rect 59778 29598 59780 29650
rect 59724 29586 59780 29598
rect 59388 29374 59390 29426
rect 59442 29374 59444 29426
rect 59388 28420 59444 29374
rect 59388 28354 59444 28364
rect 59500 29372 59668 29428
rect 59172 28252 59436 28262
rect 59228 28196 59276 28252
rect 59332 28196 59380 28252
rect 59172 28186 59436 28196
rect 59052 27806 59054 27858
rect 59106 27806 59108 27858
rect 59052 27794 59108 27806
rect 59276 27746 59332 27758
rect 59276 27694 59278 27746
rect 59330 27694 59332 27746
rect 58940 27134 58942 27186
rect 58994 27134 58996 27186
rect 58940 26740 58996 27134
rect 58940 26674 58996 26684
rect 59052 27412 59108 27422
rect 58604 26516 58660 26526
rect 58604 26422 58660 26460
rect 58940 26402 58996 26414
rect 58940 26350 58942 26402
rect 58994 26350 58996 26402
rect 58940 26292 58996 26350
rect 58828 26068 58884 26078
rect 58716 26066 58884 26068
rect 58716 26014 58830 26066
rect 58882 26014 58884 26066
rect 58716 26012 58884 26014
rect 58380 25284 58436 25294
rect 57820 25218 57876 25228
rect 58268 25282 58436 25284
rect 58268 25230 58382 25282
rect 58434 25230 58436 25282
rect 58268 25228 58436 25230
rect 57932 24836 57988 24846
rect 57932 24742 57988 24780
rect 57820 24722 57876 24734
rect 57820 24670 57822 24722
rect 57874 24670 57876 24722
rect 57820 24612 57876 24670
rect 57820 24546 57876 24556
rect 58156 24722 58212 24734
rect 58156 24670 58158 24722
rect 58210 24670 58212 24722
rect 57820 24276 57876 24286
rect 57596 23940 57652 23950
rect 57484 23938 57652 23940
rect 57484 23886 57598 23938
rect 57650 23886 57652 23938
rect 57484 23884 57652 23886
rect 57596 23874 57652 23884
rect 57372 23828 57428 23838
rect 57372 23734 57428 23772
rect 57148 23214 57150 23266
rect 57202 23214 57204 23266
rect 57148 23202 57204 23214
rect 57708 23714 57764 23726
rect 57708 23662 57710 23714
rect 57762 23662 57764 23714
rect 57708 23156 57764 23662
rect 57708 23090 57764 23100
rect 57820 23714 57876 24220
rect 58044 24052 58100 24062
rect 57820 23662 57822 23714
rect 57874 23662 57876 23714
rect 57036 22708 57092 22718
rect 56812 22484 56868 22494
rect 56588 22036 56644 22046
rect 56364 21980 56588 22036
rect 56588 20802 56644 21980
rect 56812 21588 56868 22428
rect 56812 20914 56868 21532
rect 56812 20862 56814 20914
rect 56866 20862 56868 20914
rect 56812 20850 56868 20862
rect 56588 20750 56590 20802
rect 56642 20750 56644 20802
rect 56588 20738 56644 20750
rect 55580 20692 55636 20702
rect 55356 20690 55636 20692
rect 55356 20638 55582 20690
rect 55634 20638 55636 20690
rect 55356 20636 55636 20638
rect 55580 20626 55636 20636
rect 56812 20692 56868 20702
rect 56700 20244 56756 20254
rect 55468 19906 55524 19918
rect 55468 19854 55470 19906
rect 55522 19854 55524 19906
rect 55468 19572 55524 19854
rect 56028 19908 56084 19918
rect 56028 19814 56084 19852
rect 55468 19506 55524 19516
rect 55580 19348 55636 19358
rect 55468 19346 55636 19348
rect 55468 19294 55582 19346
rect 55634 19294 55636 19346
rect 55468 19292 55636 19294
rect 55468 18564 55524 19292
rect 55580 19282 55636 19292
rect 56700 19236 56756 20188
rect 56364 19234 56756 19236
rect 56364 19182 56702 19234
rect 56754 19182 56756 19234
rect 56364 19180 56756 19182
rect 56140 19010 56196 19022
rect 56140 18958 56142 19010
rect 56194 18958 56196 19010
rect 56140 18676 56196 18958
rect 55468 18498 55524 18508
rect 55580 18620 56196 18676
rect 55580 18562 55636 18620
rect 55580 18510 55582 18562
rect 55634 18510 55636 18562
rect 55356 18450 55412 18462
rect 55356 18398 55358 18450
rect 55410 18398 55412 18450
rect 55356 16772 55412 18398
rect 55468 17554 55524 17566
rect 55468 17502 55470 17554
rect 55522 17502 55524 17554
rect 55468 17106 55524 17502
rect 55580 17556 55636 18510
rect 55692 18452 55748 18462
rect 55692 18358 55748 18396
rect 55804 18450 55860 18462
rect 55804 18398 55806 18450
rect 55858 18398 55860 18450
rect 55804 18340 55860 18398
rect 56028 18450 56084 18462
rect 56028 18398 56030 18450
rect 56082 18398 56084 18450
rect 56028 18340 56084 18398
rect 56028 18284 56196 18340
rect 55804 18228 55860 18284
rect 55804 18172 56084 18228
rect 55916 17892 55972 17902
rect 55804 17836 55916 17892
rect 55580 17500 55748 17556
rect 55468 17054 55470 17106
rect 55522 17054 55524 17106
rect 55468 17042 55524 17054
rect 55468 16884 55524 16894
rect 55468 16790 55524 16828
rect 55356 16706 55412 16716
rect 55468 16548 55524 16558
rect 55524 16492 55636 16548
rect 55468 16482 55524 16492
rect 55468 15428 55524 15438
rect 55468 15334 55524 15372
rect 54684 14530 54740 14588
rect 54684 14478 54686 14530
rect 54738 14478 54740 14530
rect 54684 14466 54740 14478
rect 55132 15092 55300 15148
rect 55580 15148 55636 16492
rect 55692 15988 55748 17500
rect 55804 16994 55860 17836
rect 55916 17826 55972 17836
rect 55804 16942 55806 16994
rect 55858 16942 55860 16994
rect 55804 16930 55860 16942
rect 55916 17666 55972 17678
rect 55916 17614 55918 17666
rect 55970 17614 55972 17666
rect 55916 16210 55972 17614
rect 56028 16884 56084 18172
rect 56028 16818 56084 16828
rect 56140 16660 56196 18284
rect 56364 17108 56420 19180
rect 56700 19170 56756 19180
rect 56812 19122 56868 20636
rect 57036 20132 57092 22652
rect 57484 22146 57540 22158
rect 57484 22094 57486 22146
rect 57538 22094 57540 22146
rect 57036 20076 57204 20132
rect 56812 19070 56814 19122
rect 56866 19070 56868 19122
rect 56812 18900 56868 19070
rect 57036 19906 57092 19918
rect 57036 19854 57038 19906
rect 57090 19854 57092 19906
rect 56588 18844 56868 18900
rect 56924 19010 56980 19022
rect 56924 18958 56926 19010
rect 56978 18958 56980 19010
rect 56476 18450 56532 18462
rect 56476 18398 56478 18450
rect 56530 18398 56532 18450
rect 56476 18116 56532 18398
rect 56476 18050 56532 18060
rect 56588 17892 56644 18844
rect 56812 18564 56868 18574
rect 56924 18564 56980 18958
rect 57036 18676 57092 19854
rect 57036 18610 57092 18620
rect 56812 18562 56980 18564
rect 56812 18510 56814 18562
rect 56866 18510 56980 18562
rect 56812 18508 56980 18510
rect 56812 18498 56868 18508
rect 56700 18450 56756 18462
rect 56700 18398 56702 18450
rect 56754 18398 56756 18450
rect 56700 18340 56756 18398
rect 56700 18274 56756 18284
rect 56588 17836 57092 17892
rect 56924 17666 56980 17678
rect 56924 17614 56926 17666
rect 56978 17614 56980 17666
rect 56364 17052 56756 17108
rect 56588 16884 56644 16894
rect 56588 16790 56644 16828
rect 55916 16158 55918 16210
rect 55970 16158 55972 16210
rect 55916 16146 55972 16158
rect 56028 16604 56196 16660
rect 56028 16212 56084 16604
rect 56028 16156 56308 16212
rect 55692 15932 55972 15988
rect 55580 15092 55748 15148
rect 54460 13860 54516 13870
rect 53564 12402 54068 12404
rect 53564 12350 53566 12402
rect 53618 12350 54068 12402
rect 53564 12348 54068 12350
rect 54236 13804 54460 13860
rect 53564 12338 53620 12348
rect 53452 12238 53454 12290
rect 53506 12238 53508 12290
rect 53452 12226 53508 12238
rect 54236 12290 54292 13804
rect 54460 13766 54516 13804
rect 54908 13748 54964 13758
rect 54908 13654 54964 13692
rect 54236 12238 54238 12290
rect 54290 12238 54292 12290
rect 54236 12226 54292 12238
rect 54348 13524 54404 13534
rect 53788 11956 53844 11966
rect 53788 11282 53844 11900
rect 54236 11844 54292 11854
rect 53788 11230 53790 11282
rect 53842 11230 53844 11282
rect 53676 10500 53732 10510
rect 53452 9940 53508 9950
rect 53452 9846 53508 9884
rect 53228 9762 53284 9772
rect 52892 9538 52948 9548
rect 53228 9044 53284 9054
rect 53004 8988 53228 9044
rect 53004 5236 53060 8988
rect 53228 8950 53284 8988
rect 53676 8596 53732 10444
rect 53788 10498 53844 11230
rect 53900 11394 53956 11406
rect 53900 11342 53902 11394
rect 53954 11342 53956 11394
rect 53900 11172 53956 11342
rect 53900 11106 53956 11116
rect 53788 10446 53790 10498
rect 53842 10446 53844 10498
rect 53788 10434 53844 10446
rect 54012 9826 54068 9838
rect 54012 9774 54014 9826
rect 54066 9774 54068 9826
rect 54012 9044 54068 9774
rect 54012 8978 54068 8988
rect 53676 8530 53732 8540
rect 54236 8372 54292 11788
rect 54348 10834 54404 13468
rect 55132 12628 55188 15092
rect 55244 14530 55300 14542
rect 55244 14478 55246 14530
rect 55298 14478 55300 14530
rect 55244 14196 55300 14478
rect 55580 14308 55636 14318
rect 55244 14130 55300 14140
rect 55468 14306 55636 14308
rect 55468 14254 55582 14306
rect 55634 14254 55636 14306
rect 55468 14252 55636 14254
rect 55468 14084 55524 14252
rect 55580 14242 55636 14252
rect 55244 13746 55300 13758
rect 55244 13694 55246 13746
rect 55298 13694 55300 13746
rect 55244 13188 55300 13694
rect 55244 13122 55300 13132
rect 55468 13186 55524 14028
rect 55580 13972 55636 13982
rect 55580 13878 55636 13916
rect 55468 13134 55470 13186
rect 55522 13134 55524 13186
rect 55468 13122 55524 13134
rect 55356 12964 55412 12974
rect 55356 12870 55412 12908
rect 55132 12572 55300 12628
rect 54908 12178 54964 12190
rect 54908 12126 54910 12178
rect 54962 12126 54964 12178
rect 54572 11956 54628 11966
rect 54460 11172 54516 11182
rect 54460 11078 54516 11116
rect 54348 10782 54350 10834
rect 54402 10782 54404 10834
rect 54348 10276 54404 10782
rect 54348 10210 54404 10220
rect 54236 8306 54292 8316
rect 53116 7364 53172 7374
rect 53116 7362 53396 7364
rect 53116 7310 53118 7362
rect 53170 7310 53396 7362
rect 53116 7308 53396 7310
rect 53116 7298 53172 7308
rect 53340 6578 53396 7308
rect 53340 6526 53342 6578
rect 53394 6526 53396 6578
rect 53340 6514 53396 6526
rect 53676 6580 53732 6590
rect 53676 6486 53732 6524
rect 54348 6580 54404 6590
rect 54348 6486 54404 6524
rect 54572 5348 54628 11900
rect 54908 11844 54964 12126
rect 54908 11778 54964 11788
rect 55132 11844 55188 11854
rect 55020 11396 55076 11406
rect 54908 11394 55076 11396
rect 54908 11342 55022 11394
rect 55074 11342 55076 11394
rect 54908 11340 55076 11342
rect 54796 11172 54852 11182
rect 54684 11170 54852 11172
rect 54684 11118 54798 11170
rect 54850 11118 54852 11170
rect 54684 11116 54852 11118
rect 54684 9940 54740 11116
rect 54796 11106 54852 11116
rect 54796 10836 54852 10846
rect 54908 10836 54964 11340
rect 55020 11330 55076 11340
rect 54796 10834 54964 10836
rect 54796 10782 54798 10834
rect 54850 10782 54964 10834
rect 54796 10780 54964 10782
rect 54796 10770 54852 10780
rect 55132 10612 55188 11788
rect 55020 10556 55188 10612
rect 54796 9940 54852 9950
rect 54684 9938 54852 9940
rect 54684 9886 54798 9938
rect 54850 9886 54852 9938
rect 54684 9884 54852 9886
rect 54796 9874 54852 9884
rect 55020 7812 55076 10556
rect 55132 10386 55188 10398
rect 55132 10334 55134 10386
rect 55186 10334 55188 10386
rect 55132 10276 55188 10334
rect 55132 8148 55188 10220
rect 55244 8260 55300 12572
rect 55692 9380 55748 15092
rect 55916 14196 55972 15932
rect 56140 15986 56196 15998
rect 56140 15934 56142 15986
rect 56194 15934 56196 15986
rect 56028 15316 56084 15326
rect 56028 15222 56084 15260
rect 56140 14980 56196 15934
rect 56140 14914 56196 14924
rect 56140 14644 56196 14654
rect 56252 14644 56308 16156
rect 56588 15764 56644 15774
rect 56588 15538 56644 15708
rect 56588 15486 56590 15538
rect 56642 15486 56644 15538
rect 56588 15474 56644 15486
rect 56700 15316 56756 17052
rect 56924 17106 56980 17614
rect 56924 17054 56926 17106
rect 56978 17054 56980 17106
rect 56924 17042 56980 17054
rect 55916 14130 55972 14140
rect 56028 14642 56308 14644
rect 56028 14590 56142 14642
rect 56194 14590 56308 14642
rect 56028 14588 56308 14590
rect 56588 15260 56756 15316
rect 56812 16994 56868 17006
rect 56812 16942 56814 16994
rect 56866 16942 56868 16994
rect 56812 15316 56868 16942
rect 56924 16436 56980 16446
rect 56924 15876 56980 16380
rect 57036 16100 57092 17836
rect 57148 17778 57204 20076
rect 57260 19236 57316 19246
rect 57260 19234 57428 19236
rect 57260 19182 57262 19234
rect 57314 19182 57428 19234
rect 57260 19180 57428 19182
rect 57260 19170 57316 19180
rect 57260 18452 57316 18462
rect 57260 18358 57316 18396
rect 57148 17726 57150 17778
rect 57202 17726 57204 17778
rect 57148 17714 57204 17726
rect 57260 18004 57316 18014
rect 57260 16436 57316 17948
rect 57260 16370 57316 16380
rect 57260 16100 57316 16110
rect 57036 16098 57316 16100
rect 57036 16046 57262 16098
rect 57314 16046 57316 16098
rect 57036 16044 57316 16046
rect 57260 16034 57316 16044
rect 57260 15876 57316 15886
rect 56924 15820 57260 15876
rect 56924 15540 56980 15550
rect 56924 15446 56980 15484
rect 57260 15538 57316 15820
rect 57260 15486 57262 15538
rect 57314 15486 57316 15538
rect 57260 15474 57316 15486
rect 55916 13860 55972 13870
rect 55804 13188 55860 13198
rect 55804 13074 55860 13132
rect 55804 13022 55806 13074
rect 55858 13022 55860 13074
rect 55804 13010 55860 13022
rect 55804 12404 55860 12414
rect 55916 12404 55972 13804
rect 56028 13300 56084 14588
rect 56140 14578 56196 14588
rect 56588 14532 56644 15260
rect 56812 15250 56868 15260
rect 57372 15428 57428 19180
rect 57484 17108 57540 22094
rect 57596 21812 57652 21822
rect 57596 21698 57652 21756
rect 57596 21646 57598 21698
rect 57650 21646 57652 21698
rect 57596 21634 57652 21646
rect 57820 21140 57876 23662
rect 57932 23716 57988 23726
rect 57932 23622 57988 23660
rect 58044 22482 58100 23996
rect 58044 22430 58046 22482
rect 58098 22430 58100 22482
rect 58044 22418 58100 22430
rect 58156 23154 58212 24670
rect 58268 24612 58324 25228
rect 58380 25218 58436 25228
rect 58716 24948 58772 26012
rect 58828 26002 58884 26012
rect 58940 25618 58996 26236
rect 58940 25566 58942 25618
rect 58994 25566 58996 25618
rect 58940 25554 58996 25566
rect 59052 25284 59108 27356
rect 59276 27074 59332 27694
rect 59388 27188 59444 27198
rect 59500 27188 59556 29372
rect 59612 29204 59668 29214
rect 59612 29110 59668 29148
rect 59612 28980 59668 28990
rect 59612 28866 59668 28924
rect 59612 28814 59614 28866
rect 59666 28814 59668 28866
rect 59612 28802 59668 28814
rect 59612 28644 59668 28654
rect 59612 27970 59668 28588
rect 59836 28420 59892 30380
rect 60060 29986 60116 30716
rect 60060 29934 60062 29986
rect 60114 29934 60116 29986
rect 60060 29922 60116 29934
rect 60172 30100 60228 33180
rect 60396 31892 60452 34078
rect 60732 34130 60788 34188
rect 60732 34078 60734 34130
rect 60786 34078 60788 34130
rect 60732 32562 60788 34078
rect 60844 33572 60900 34524
rect 60844 33506 60900 33516
rect 61068 33346 61124 35420
rect 64092 35140 64148 36654
rect 65436 35924 65492 35934
rect 65436 35830 65492 35868
rect 64428 35812 64484 35822
rect 64428 35698 64484 35756
rect 64428 35646 64430 35698
rect 64482 35646 64484 35698
rect 64428 35634 64484 35646
rect 65660 35252 65716 39200
rect 65884 36484 65940 36494
rect 65884 36258 65940 36428
rect 66556 36484 66612 36494
rect 66556 36390 66612 36428
rect 65884 36206 65886 36258
rect 65938 36206 65940 36258
rect 65884 35700 65940 36206
rect 67452 36258 67508 36270
rect 67452 36206 67454 36258
rect 67506 36206 67508 36258
rect 65884 35634 65940 35644
rect 67340 35810 67396 35822
rect 67340 35758 67342 35810
rect 67394 35758 67396 35810
rect 65660 35186 65716 35196
rect 64092 35074 64148 35084
rect 64764 34914 64820 34926
rect 64764 34862 64766 34914
rect 64818 34862 64820 34914
rect 61068 33294 61070 33346
rect 61122 33294 61124 33346
rect 61068 33282 61124 33294
rect 61292 34802 61348 34814
rect 61292 34750 61294 34802
rect 61346 34750 61348 34802
rect 61292 32788 61348 34750
rect 63532 34690 63588 34702
rect 63532 34638 63534 34690
rect 63586 34638 63588 34690
rect 63532 34356 63588 34638
rect 63532 34290 63588 34300
rect 64764 34132 64820 34862
rect 65548 34804 65604 34814
rect 65324 34802 65604 34804
rect 65324 34750 65550 34802
rect 65602 34750 65604 34802
rect 65324 34748 65604 34750
rect 65324 34354 65380 34748
rect 65548 34738 65604 34748
rect 65324 34302 65326 34354
rect 65378 34302 65380 34354
rect 65324 34290 65380 34302
rect 66444 34244 66500 34254
rect 66444 34150 66500 34188
rect 67340 34244 67396 35758
rect 67452 35364 67508 36206
rect 67452 35298 67508 35308
rect 67676 35698 67732 35710
rect 67676 35646 67678 35698
rect 67730 35646 67732 35698
rect 67676 35308 67732 35646
rect 67676 35252 67844 35308
rect 67340 34178 67396 34188
rect 67676 35026 67732 35038
rect 67676 34974 67678 35026
rect 67730 34974 67732 35026
rect 61516 34020 61572 34030
rect 63644 34020 63700 34030
rect 61516 34018 61684 34020
rect 61516 33966 61518 34018
rect 61570 33966 61684 34018
rect 61516 33964 61684 33966
rect 61516 33954 61572 33964
rect 61292 32722 61348 32732
rect 60732 32510 60734 32562
rect 60786 32510 60788 32562
rect 60732 32498 60788 32510
rect 61516 32452 61572 32462
rect 60956 32450 61572 32452
rect 60956 32398 61518 32450
rect 61570 32398 61572 32450
rect 60956 32396 61572 32398
rect 60956 32002 61012 32396
rect 61516 32386 61572 32396
rect 60956 31950 60958 32002
rect 61010 31950 61012 32002
rect 60956 31938 61012 31950
rect 60396 31826 60452 31836
rect 61628 31890 61684 33964
rect 63644 33926 63700 33964
rect 61964 33572 62020 33582
rect 61964 33478 62020 33516
rect 63644 32450 63700 32462
rect 63644 32398 63646 32450
rect 63698 32398 63700 32450
rect 63644 32116 63700 32398
rect 63644 32050 63700 32060
rect 64428 32452 64484 32462
rect 61628 31838 61630 31890
rect 61682 31838 61684 31890
rect 61628 31826 61684 31838
rect 60844 31780 60900 31790
rect 60620 31668 60676 31678
rect 60620 31574 60676 31612
rect 60844 31666 60900 31724
rect 61516 31780 61572 31790
rect 60844 31614 60846 31666
rect 60898 31614 60900 31666
rect 60844 31602 60900 31614
rect 61292 31666 61348 31678
rect 61292 31614 61294 31666
rect 61346 31614 61348 31666
rect 60396 30996 60452 31006
rect 59948 29428 60004 29438
rect 59948 29334 60004 29372
rect 60172 28980 60228 30044
rect 60284 30548 60340 30558
rect 60284 29876 60340 30492
rect 60396 29988 60452 30940
rect 61068 30660 61124 30670
rect 60508 30212 60564 30222
rect 60508 30118 60564 30156
rect 60956 30212 61012 30250
rect 60956 30146 61012 30156
rect 60396 29922 60452 29932
rect 60732 30098 60788 30110
rect 60732 30046 60734 30098
rect 60786 30046 60788 30098
rect 60284 29652 60340 29820
rect 60396 29652 60452 29662
rect 60284 29650 60676 29652
rect 60284 29598 60398 29650
rect 60450 29598 60676 29650
rect 60284 29596 60676 29598
rect 60396 29586 60452 29596
rect 60172 28914 60228 28924
rect 59948 28868 60004 28878
rect 59948 28774 60004 28812
rect 59948 28644 60004 28654
rect 59948 28642 60564 28644
rect 59948 28590 59950 28642
rect 60002 28590 60564 28642
rect 59948 28588 60564 28590
rect 59948 28578 60004 28588
rect 60284 28420 60340 28430
rect 59836 28364 60004 28420
rect 59612 27918 59614 27970
rect 59666 27918 59668 27970
rect 59612 27906 59668 27918
rect 59388 27186 59556 27188
rect 59388 27134 59390 27186
rect 59442 27134 59556 27186
rect 59388 27132 59556 27134
rect 59612 27244 59892 27300
rect 59388 27122 59444 27132
rect 59276 27022 59278 27074
rect 59330 27022 59332 27074
rect 59276 26908 59332 27022
rect 59612 26962 59668 27244
rect 59612 26910 59614 26962
rect 59666 26910 59668 26962
rect 59276 26852 59556 26908
rect 59612 26898 59668 26910
rect 59724 27074 59780 27086
rect 59724 27022 59726 27074
rect 59778 27022 59780 27074
rect 59172 26684 59436 26694
rect 59228 26628 59276 26684
rect 59332 26628 59380 26684
rect 59172 26618 59436 26628
rect 59164 26404 59220 26414
rect 59500 26404 59556 26852
rect 59612 26516 59668 26526
rect 59724 26516 59780 27022
rect 59612 26514 59780 26516
rect 59612 26462 59614 26514
rect 59666 26462 59780 26514
rect 59612 26460 59780 26462
rect 59612 26450 59668 26460
rect 59164 26402 59556 26404
rect 59164 26350 59166 26402
rect 59218 26350 59502 26402
rect 59554 26350 59556 26402
rect 59164 26348 59556 26350
rect 59164 26338 59220 26348
rect 59500 26338 59556 26348
rect 59724 26292 59780 26302
rect 59836 26292 59892 27244
rect 59948 26908 60004 28364
rect 60172 27858 60228 27870
rect 60172 27806 60174 27858
rect 60226 27806 60228 27858
rect 60172 27188 60228 27806
rect 60172 27122 60228 27132
rect 60284 27076 60340 28364
rect 60508 28420 60564 28588
rect 60508 28082 60564 28364
rect 60508 28030 60510 28082
rect 60562 28030 60564 28082
rect 60508 28018 60564 28030
rect 60620 27860 60676 29596
rect 60732 28756 60788 30046
rect 60844 29540 60900 29550
rect 60844 29446 60900 29484
rect 60956 29426 61012 29438
rect 60956 29374 60958 29426
rect 61010 29374 61012 29426
rect 60956 28868 61012 29374
rect 60956 28802 61012 28812
rect 60732 28700 60900 28756
rect 60284 26908 60340 27020
rect 60508 27804 60676 27860
rect 60732 28418 60788 28430
rect 60732 28366 60734 28418
rect 60786 28366 60788 28418
rect 60732 27858 60788 28366
rect 60844 28308 60900 28700
rect 60844 28242 60900 28252
rect 60732 27806 60734 27858
rect 60786 27806 60788 27858
rect 59948 26852 60116 26908
rect 60284 26852 60452 26908
rect 59948 26516 60004 26526
rect 59948 26422 60004 26460
rect 59780 26236 59892 26292
rect 59724 26198 59780 26236
rect 59612 25506 59668 25518
rect 59612 25454 59614 25506
rect 59666 25454 59668 25506
rect 58380 24892 58772 24948
rect 58940 25228 59108 25284
rect 59388 25284 59444 25294
rect 59444 25228 59556 25284
rect 58380 24834 58436 24892
rect 58380 24782 58382 24834
rect 58434 24782 58436 24834
rect 58380 24770 58436 24782
rect 58716 24724 58772 24734
rect 58268 24556 58660 24612
rect 58156 23102 58158 23154
rect 58210 23102 58212 23154
rect 58156 23044 58212 23102
rect 58380 24052 58436 24062
rect 58380 23154 58436 23996
rect 58492 23716 58548 23726
rect 58492 23622 58548 23660
rect 58604 23714 58660 24556
rect 58716 24050 58772 24668
rect 58828 24610 58884 24622
rect 58828 24558 58830 24610
rect 58882 24558 58884 24610
rect 58828 24276 58884 24558
rect 58828 24210 58884 24220
rect 58716 23998 58718 24050
rect 58770 23998 58772 24050
rect 58716 23986 58772 23998
rect 58828 23940 58884 23950
rect 58940 23940 58996 25228
rect 59388 25218 59444 25228
rect 59172 25116 59436 25126
rect 59228 25060 59276 25116
rect 59332 25060 59380 25116
rect 59172 25050 59436 25060
rect 59276 24948 59332 24958
rect 59500 24948 59556 25228
rect 59612 25060 59668 25454
rect 59612 24994 59668 25004
rect 59836 25508 59892 25518
rect 60060 25508 60116 26852
rect 59836 25506 60116 25508
rect 59836 25454 59838 25506
rect 59890 25454 60116 25506
rect 59836 25452 60116 25454
rect 59276 24946 59556 24948
rect 59276 24894 59278 24946
rect 59330 24894 59556 24946
rect 59276 24892 59556 24894
rect 59276 24882 59332 24892
rect 58828 23938 58996 23940
rect 58828 23886 58830 23938
rect 58882 23886 58996 23938
rect 58828 23884 58996 23886
rect 58828 23874 58884 23884
rect 59052 23828 59108 23838
rect 59052 23734 59108 23772
rect 59388 23826 59444 23838
rect 59388 23774 59390 23826
rect 59442 23774 59444 23826
rect 58604 23662 58606 23714
rect 58658 23662 58660 23714
rect 58380 23102 58382 23154
rect 58434 23102 58436 23154
rect 58380 23090 58436 23102
rect 58156 21586 58212 22988
rect 58492 23042 58548 23054
rect 58492 22990 58494 23042
rect 58546 22990 58548 23042
rect 58268 22370 58324 22382
rect 58268 22318 58270 22370
rect 58322 22318 58324 22370
rect 58268 22036 58324 22318
rect 58268 21970 58324 21980
rect 58492 21812 58548 22990
rect 58156 21534 58158 21586
rect 58210 21534 58212 21586
rect 58156 21522 58212 21534
rect 58268 21756 58548 21812
rect 57708 21084 57876 21140
rect 57484 17042 57540 17052
rect 57596 17668 57652 17678
rect 57596 16994 57652 17612
rect 57596 16942 57598 16994
rect 57650 16942 57652 16994
rect 57596 16930 57652 16942
rect 57484 16884 57540 16894
rect 57484 16212 57540 16828
rect 57484 16146 57540 16156
rect 57148 15204 57204 15214
rect 56812 15092 56868 15102
rect 56252 14530 56644 14532
rect 56252 14478 56590 14530
rect 56642 14478 56644 14530
rect 56252 14476 56644 14478
rect 56140 13972 56196 13982
rect 56252 13972 56308 14476
rect 56588 14466 56644 14476
rect 56700 14532 56756 14542
rect 56700 14438 56756 14476
rect 56140 13970 56308 13972
rect 56140 13918 56142 13970
rect 56194 13918 56308 13970
rect 56140 13916 56308 13918
rect 56364 14196 56420 14206
rect 56140 13906 56196 13916
rect 56028 13234 56084 13244
rect 56252 13186 56308 13198
rect 56252 13134 56254 13186
rect 56306 13134 56308 13186
rect 56252 13074 56308 13134
rect 56252 13022 56254 13074
rect 56306 13022 56308 13074
rect 56252 13010 56308 13022
rect 55804 12402 55972 12404
rect 55804 12350 55806 12402
rect 55858 12350 55972 12402
rect 55804 12348 55972 12350
rect 55804 12338 55860 12348
rect 56364 12180 56420 14140
rect 56812 13972 56868 15036
rect 57036 14644 57092 14654
rect 57036 14530 57092 14588
rect 57036 14478 57038 14530
rect 57090 14478 57092 14530
rect 57036 14466 57092 14478
rect 56924 14420 56980 14430
rect 56924 14326 56980 14364
rect 56364 12114 56420 12124
rect 56476 13748 56532 13758
rect 56476 11956 56532 13692
rect 56028 11900 56532 11956
rect 56700 13746 56756 13758
rect 56700 13694 56702 13746
rect 56754 13694 56756 13746
rect 56700 12962 56756 13694
rect 56700 12910 56702 12962
rect 56754 12910 56756 12962
rect 56700 11956 56756 12910
rect 56812 12962 56868 13916
rect 56812 12910 56814 12962
rect 56866 12910 56868 12962
rect 56812 12898 56868 12910
rect 56924 13636 56980 13646
rect 56924 12964 56980 13580
rect 57036 13076 57092 13086
rect 57036 12982 57092 13020
rect 56812 12404 56868 12414
rect 56924 12404 56980 12908
rect 57148 12962 57204 15148
rect 57260 14868 57316 14878
rect 57260 14754 57316 14812
rect 57260 14702 57262 14754
rect 57314 14702 57316 14754
rect 57260 14690 57316 14702
rect 57372 14756 57428 15372
rect 57596 15426 57652 15438
rect 57596 15374 57598 15426
rect 57650 15374 57652 15426
rect 57596 15204 57652 15374
rect 57596 15138 57652 15148
rect 57372 14690 57428 14700
rect 57372 14530 57428 14542
rect 57372 14478 57374 14530
rect 57426 14478 57428 14530
rect 57372 13076 57428 14478
rect 57596 14420 57652 14430
rect 57596 14326 57652 14364
rect 57372 13010 57428 13020
rect 57148 12910 57150 12962
rect 57202 12910 57204 12962
rect 57148 12898 57204 12910
rect 56812 12402 56980 12404
rect 56812 12350 56814 12402
rect 56866 12350 56980 12402
rect 56812 12348 56980 12350
rect 57036 12852 57092 12862
rect 56812 12338 56868 12348
rect 56924 12068 56980 12078
rect 56028 11506 56084 11900
rect 56700 11890 56756 11900
rect 56812 12012 56924 12068
rect 56028 11454 56030 11506
rect 56082 11454 56084 11506
rect 56028 11442 56084 11454
rect 56812 11396 56868 12012
rect 56924 12002 56980 12012
rect 57036 11844 57092 12796
rect 57372 12404 57428 12414
rect 57372 12310 57428 12348
rect 57260 12292 57316 12302
rect 57036 11778 57092 11788
rect 57148 12236 57260 12292
rect 57148 11620 57204 12236
rect 57260 12226 57316 12236
rect 57708 11844 57764 21084
rect 58044 20804 58100 20814
rect 58268 20804 58324 21756
rect 58380 21588 58436 21598
rect 58380 21494 58436 21532
rect 58492 21474 58548 21486
rect 58492 21422 58494 21474
rect 58546 21422 58548 21474
rect 58044 20802 58212 20804
rect 58044 20750 58046 20802
rect 58098 20750 58212 20802
rect 58044 20748 58212 20750
rect 58268 20748 58436 20804
rect 58044 20738 58100 20748
rect 58044 19908 58100 19918
rect 57820 19236 57876 19246
rect 57820 19142 57876 19180
rect 58044 18676 58100 19852
rect 58156 19460 58212 20748
rect 58268 20578 58324 20590
rect 58268 20526 58270 20578
rect 58322 20526 58324 20578
rect 58268 20132 58324 20526
rect 58268 20066 58324 20076
rect 58268 19460 58324 19470
rect 58156 19458 58324 19460
rect 58156 19406 58270 19458
rect 58322 19406 58324 19458
rect 58156 19404 58324 19406
rect 58268 19394 58324 19404
rect 58380 19124 58436 20748
rect 58268 19068 58436 19124
rect 58044 18620 58212 18676
rect 58044 18452 58100 18462
rect 58044 18358 58100 18396
rect 57820 18340 57876 18350
rect 57820 17778 57876 18284
rect 57820 17726 57822 17778
rect 57874 17726 57876 17778
rect 57820 17714 57876 17726
rect 58156 17892 58212 18620
rect 57932 17668 57988 17678
rect 58156 17668 58212 17836
rect 57932 17666 58212 17668
rect 57932 17614 57934 17666
rect 57986 17614 58212 17666
rect 57932 17612 58212 17614
rect 57932 17602 57988 17612
rect 57820 17442 57876 17454
rect 57820 17390 57822 17442
rect 57874 17390 57876 17442
rect 57820 15204 57876 17390
rect 58156 17442 58212 17454
rect 58156 17390 58158 17442
rect 58210 17390 58212 17442
rect 57820 15138 57876 15148
rect 57932 17108 57988 17118
rect 57932 16212 57988 17052
rect 57932 16098 57988 16156
rect 57932 16046 57934 16098
rect 57986 16046 57988 16098
rect 57932 15148 57988 16046
rect 58044 15764 58100 15774
rect 58044 15538 58100 15708
rect 58044 15486 58046 15538
rect 58098 15486 58100 15538
rect 58044 15474 58100 15486
rect 57932 15092 58100 15148
rect 57932 14530 57988 14542
rect 57932 14478 57934 14530
rect 57986 14478 57988 14530
rect 57820 13412 57876 13422
rect 57820 12962 57876 13356
rect 57932 13300 57988 14478
rect 58044 13972 58100 15092
rect 58156 15092 58212 17390
rect 58156 15026 58212 15036
rect 58268 14084 58324 19068
rect 58380 17556 58436 17566
rect 58380 17332 58436 17500
rect 58492 17332 58548 21422
rect 58604 20356 58660 23662
rect 59388 23716 59444 23774
rect 59500 23826 59556 24892
rect 59500 23774 59502 23826
rect 59554 23774 59556 23826
rect 59500 23762 59556 23774
rect 59612 24836 59668 24846
rect 59388 23650 59444 23660
rect 59172 23548 59436 23558
rect 59228 23492 59276 23548
rect 59332 23492 59380 23548
rect 59172 23482 59436 23492
rect 59612 23380 59668 24780
rect 59724 24724 59780 24734
rect 59724 24630 59780 24668
rect 59836 24612 59892 25452
rect 59276 23324 59668 23380
rect 59724 23714 59780 23726
rect 59724 23662 59726 23714
rect 59778 23662 59780 23714
rect 59276 22260 59332 23324
rect 59724 23266 59780 23662
rect 59724 23214 59726 23266
rect 59778 23214 59780 23266
rect 59724 23202 59780 23214
rect 59500 23156 59556 23166
rect 59500 23062 59556 23100
rect 59836 23044 59892 24556
rect 59948 25060 60004 25070
rect 59948 24388 60004 25004
rect 59948 24322 60004 24332
rect 60060 24834 60116 24846
rect 60060 24782 60062 24834
rect 60114 24782 60116 24834
rect 60060 24164 60116 24782
rect 60396 24836 60452 26852
rect 60396 24770 60452 24780
rect 60396 24610 60452 24622
rect 60396 24558 60398 24610
rect 60450 24558 60452 24610
rect 60060 24108 60340 24164
rect 59724 22988 59892 23044
rect 59948 23940 60004 23950
rect 59052 22258 59332 22260
rect 59052 22206 59278 22258
rect 59330 22206 59332 22258
rect 59052 22204 59332 22206
rect 59052 21812 59108 22204
rect 59276 22194 59332 22204
rect 59500 22372 59556 22382
rect 59172 21980 59436 21990
rect 59228 21924 59276 21980
rect 59332 21924 59380 21980
rect 59172 21914 59436 21924
rect 59052 21746 59108 21756
rect 59500 21700 59556 22316
rect 59164 21698 59556 21700
rect 59164 21646 59502 21698
rect 59554 21646 59556 21698
rect 59164 21644 59556 21646
rect 59052 20916 59108 20926
rect 59164 20916 59220 21644
rect 59500 21634 59556 21644
rect 59612 22260 59668 22270
rect 59052 20914 59220 20916
rect 59052 20862 59054 20914
rect 59106 20862 59220 20914
rect 59052 20860 59220 20862
rect 59388 20916 59444 20926
rect 59612 20916 59668 22204
rect 59724 21810 59780 22988
rect 59948 22708 60004 23884
rect 59948 22642 60004 22652
rect 60060 23604 60116 23614
rect 60060 22484 60116 23548
rect 60284 23380 60340 24108
rect 60396 24052 60452 24558
rect 60396 23986 60452 23996
rect 60396 23380 60452 23390
rect 60284 23378 60452 23380
rect 60284 23326 60398 23378
rect 60450 23326 60452 23378
rect 60284 23324 60452 23326
rect 60508 23380 60564 27804
rect 60620 27188 60676 27198
rect 60620 27094 60676 27132
rect 60732 26516 60788 27806
rect 60732 26450 60788 26460
rect 60956 24610 61012 24622
rect 60956 24558 60958 24610
rect 61010 24558 61012 24610
rect 60620 23716 60676 23726
rect 60956 23716 61012 24558
rect 60676 23660 61012 23716
rect 60620 23622 60676 23660
rect 60620 23380 60676 23390
rect 60508 23324 60620 23380
rect 60396 23314 60452 23324
rect 60620 23286 60676 23324
rect 60732 23156 60788 23660
rect 61068 23604 61124 30604
rect 61292 30322 61348 31614
rect 61516 31666 61572 31724
rect 61516 31614 61518 31666
rect 61570 31614 61572 31666
rect 61516 31602 61572 31614
rect 61292 30270 61294 30322
rect 61346 30270 61348 30322
rect 61292 30258 61348 30270
rect 61180 30210 61236 30222
rect 61180 30158 61182 30210
rect 61234 30158 61236 30210
rect 61180 29876 61236 30158
rect 62636 30212 62692 30222
rect 61404 30098 61460 30110
rect 61404 30046 61406 30098
rect 61458 30046 61460 30098
rect 61404 29988 61460 30046
rect 61740 30100 61796 30110
rect 61740 30006 61796 30044
rect 62076 29988 62132 29998
rect 61404 29922 61460 29932
rect 61964 29986 62132 29988
rect 61964 29934 62078 29986
rect 62130 29934 62132 29986
rect 61964 29932 62132 29934
rect 61180 29810 61236 29820
rect 61180 29428 61236 29438
rect 61180 27860 61236 29372
rect 61516 28754 61572 28766
rect 61516 28702 61518 28754
rect 61570 28702 61572 28754
rect 61404 28644 61460 28654
rect 61292 28532 61348 28542
rect 61292 28082 61348 28476
rect 61292 28030 61294 28082
rect 61346 28030 61348 28082
rect 61292 28018 61348 28030
rect 61404 28082 61460 28588
rect 61404 28030 61406 28082
rect 61458 28030 61460 28082
rect 61404 28018 61460 28030
rect 61516 28308 61572 28702
rect 61628 28642 61684 28654
rect 61628 28590 61630 28642
rect 61682 28590 61684 28642
rect 61628 28420 61684 28590
rect 61628 28354 61684 28364
rect 61964 28308 62020 29932
rect 62076 29922 62132 29932
rect 62636 29650 62692 30156
rect 62636 29598 62638 29650
rect 62690 29598 62692 29650
rect 62636 29586 62692 29598
rect 62748 29540 62804 29550
rect 62076 29428 62132 29438
rect 62076 28644 62132 29372
rect 62188 29428 62244 29438
rect 62412 29428 62468 29438
rect 62188 29426 62356 29428
rect 62188 29374 62190 29426
rect 62242 29374 62356 29426
rect 62188 29372 62356 29374
rect 62188 29362 62244 29372
rect 62076 28550 62132 28588
rect 62300 28642 62356 29372
rect 62412 29334 62468 29372
rect 62748 29426 62804 29484
rect 62748 29374 62750 29426
rect 62802 29374 62804 29426
rect 62748 29362 62804 29374
rect 62972 29426 63028 29438
rect 62972 29374 62974 29426
rect 63026 29374 63028 29426
rect 62300 28590 62302 28642
rect 62354 28590 62356 28642
rect 62300 28578 62356 28590
rect 62636 28530 62692 28542
rect 62636 28478 62638 28530
rect 62690 28478 62692 28530
rect 62524 28420 62580 28430
rect 62076 28308 62132 28318
rect 61964 28252 62076 28308
rect 61180 27766 61236 27804
rect 61404 27412 61460 27422
rect 61516 27412 61572 28252
rect 62076 28242 62132 28252
rect 61460 27356 61572 27412
rect 62076 27858 62132 27870
rect 62076 27806 62078 27858
rect 62130 27806 62132 27858
rect 61404 27346 61460 27356
rect 62076 27186 62132 27806
rect 62524 27858 62580 28364
rect 62636 28308 62692 28478
rect 62972 28532 63028 29374
rect 62972 28466 63028 28476
rect 62636 28242 62692 28252
rect 62524 27806 62526 27858
rect 62578 27806 62580 27858
rect 62524 27794 62580 27806
rect 63420 27858 63476 27870
rect 63420 27806 63422 27858
rect 63474 27806 63476 27858
rect 62300 27634 62356 27646
rect 62300 27582 62302 27634
rect 62354 27582 62356 27634
rect 62300 27300 62356 27582
rect 62300 27234 62356 27244
rect 63420 27300 63476 27806
rect 63420 27234 63476 27244
rect 63532 27636 63588 27646
rect 62076 27134 62078 27186
rect 62130 27134 62132 27186
rect 61628 27076 61684 27114
rect 61628 27010 61684 27020
rect 61292 26964 61348 27002
rect 62076 26964 62132 27134
rect 62412 27188 62468 27198
rect 62076 26908 62356 26964
rect 61292 26898 61348 26908
rect 61628 26852 61684 26862
rect 61292 26516 61348 26526
rect 61292 23940 61348 26460
rect 61628 26514 61684 26796
rect 61628 26462 61630 26514
rect 61682 26462 61684 26514
rect 61628 26450 61684 26462
rect 61964 26404 62020 26414
rect 61964 26402 62244 26404
rect 61964 26350 61966 26402
rect 62018 26350 62244 26402
rect 61964 26348 62244 26350
rect 61964 26338 62020 26348
rect 62188 26292 62244 26348
rect 62188 24722 62244 26236
rect 62188 24670 62190 24722
rect 62242 24670 62244 24722
rect 61852 24612 61908 24622
rect 61628 24388 61684 24398
rect 61404 24164 61460 24202
rect 61404 24098 61460 24108
rect 61292 23874 61348 23884
rect 61628 23938 61684 24332
rect 61628 23886 61630 23938
rect 61682 23886 61684 23938
rect 61628 23874 61684 23886
rect 61852 24050 61908 24556
rect 61852 23998 61854 24050
rect 61906 23998 61908 24050
rect 61068 23548 61236 23604
rect 61180 23268 61236 23548
rect 61740 23380 61796 23390
rect 61740 23286 61796 23324
rect 61180 23174 61236 23212
rect 60732 23062 60788 23100
rect 60956 23154 61012 23166
rect 60956 23102 60958 23154
rect 61010 23102 61012 23154
rect 60172 23044 60228 23054
rect 60172 22950 60228 22988
rect 60060 22428 60228 22484
rect 60060 22260 60116 22270
rect 59724 21758 59726 21810
rect 59778 21758 59780 21810
rect 59724 21746 59780 21758
rect 59836 21812 59892 21822
rect 59836 21718 59892 21756
rect 60060 21810 60116 22204
rect 60060 21758 60062 21810
rect 60114 21758 60116 21810
rect 60060 21746 60116 21758
rect 59948 21586 60004 21598
rect 59948 21534 59950 21586
rect 60002 21534 60004 21586
rect 59948 21476 60004 21534
rect 59948 21410 60004 21420
rect 59388 20914 59668 20916
rect 59388 20862 59390 20914
rect 59442 20862 59668 20914
rect 59388 20860 59668 20862
rect 59724 21028 59780 21038
rect 59052 20850 59108 20860
rect 59388 20850 59444 20860
rect 59172 20412 59436 20422
rect 59228 20356 59276 20412
rect 59332 20356 59380 20412
rect 59724 20356 59780 20972
rect 59172 20346 59436 20356
rect 58604 20290 58660 20300
rect 59612 20300 59724 20356
rect 59164 20132 59220 20142
rect 59164 20038 59220 20076
rect 59388 20020 59444 20030
rect 58604 19234 58660 19246
rect 58604 19182 58606 19234
rect 58658 19182 58660 19234
rect 58604 18676 58660 19182
rect 59276 19236 59332 19246
rect 59276 19142 59332 19180
rect 59388 19124 59444 19964
rect 59388 19030 59444 19068
rect 59172 18844 59436 18854
rect 59228 18788 59276 18844
rect 59332 18788 59380 18844
rect 59172 18778 59436 18788
rect 58604 18610 58660 18620
rect 58940 18676 58996 18686
rect 58828 18452 58884 18462
rect 58716 18004 58772 18014
rect 58716 17666 58772 17948
rect 58828 17778 58884 18396
rect 58828 17726 58830 17778
rect 58882 17726 58884 17778
rect 58828 17714 58884 17726
rect 58716 17614 58718 17666
rect 58770 17614 58772 17666
rect 58716 17602 58772 17614
rect 58940 17666 58996 18620
rect 58940 17614 58942 17666
rect 58994 17614 58996 17666
rect 58940 17602 58996 17614
rect 59388 17668 59444 17678
rect 59388 17574 59444 17612
rect 59164 17444 59220 17454
rect 59164 17442 59556 17444
rect 59164 17390 59166 17442
rect 59218 17390 59556 17442
rect 59164 17388 59556 17390
rect 59164 17378 59220 17388
rect 58604 17332 58660 17342
rect 58492 17276 58604 17332
rect 58380 17266 58436 17276
rect 58604 17266 58660 17276
rect 58772 17332 58828 17342
rect 58828 17276 58996 17332
rect 58772 17266 58828 17276
rect 58492 16884 58548 16894
rect 58492 16790 58548 16828
rect 58380 16436 58436 16446
rect 58380 16210 58436 16380
rect 58380 16158 58382 16210
rect 58434 16158 58436 16210
rect 58380 14308 58436 16158
rect 58940 16210 58996 17276
rect 59172 17276 59436 17286
rect 59228 17220 59276 17276
rect 59332 17220 59380 17276
rect 59172 17210 59436 17220
rect 58940 16158 58942 16210
rect 58994 16158 58996 16210
rect 58940 15876 58996 16158
rect 58940 15810 58996 15820
rect 59052 16884 59108 16894
rect 59052 15540 59108 16828
rect 59388 16212 59444 16222
rect 59388 16118 59444 16156
rect 59172 15708 59436 15718
rect 59228 15652 59276 15708
rect 59332 15652 59380 15708
rect 59172 15642 59436 15652
rect 59500 15540 59556 17388
rect 59052 15484 59220 15540
rect 58380 14242 58436 14252
rect 58492 15428 58548 15438
rect 58268 14018 58324 14028
rect 58044 13916 58212 13972
rect 58044 13748 58100 13758
rect 58044 13654 58100 13692
rect 57932 13244 58100 13300
rect 57820 12910 57822 12962
rect 57874 12910 57876 12962
rect 57820 12898 57876 12910
rect 57932 12852 57988 12862
rect 57932 12758 57988 12796
rect 58044 12404 58100 13244
rect 58156 12628 58212 13916
rect 58380 13746 58436 13758
rect 58380 13694 58382 13746
rect 58434 13694 58436 13746
rect 58380 13636 58436 13694
rect 58380 13570 58436 13580
rect 58156 12562 58212 12572
rect 58380 13300 58436 13310
rect 58380 12964 58436 13244
rect 58492 13074 58548 15372
rect 58828 14756 58884 14766
rect 58492 13022 58494 13074
rect 58546 13022 58548 13074
rect 58492 13010 58548 13022
rect 58604 14532 58660 14542
rect 58156 12404 58212 12414
rect 58044 12402 58212 12404
rect 58044 12350 58158 12402
rect 58210 12350 58212 12402
rect 58044 12348 58212 12350
rect 58156 12338 58212 12348
rect 58380 12402 58436 12908
rect 58380 12350 58382 12402
rect 58434 12350 58436 12402
rect 58380 12338 58436 12350
rect 57932 12292 57988 12302
rect 57932 12178 57988 12236
rect 57932 12126 57934 12178
rect 57986 12126 57988 12178
rect 57932 12114 57988 12126
rect 58044 12180 58100 12190
rect 58044 11956 58100 12124
rect 58268 12180 58324 12190
rect 58268 12086 58324 12124
rect 56700 11340 56868 11396
rect 56924 11564 57204 11620
rect 57260 11788 57764 11844
rect 57820 11900 58044 11956
rect 56700 10948 56756 11340
rect 55804 10892 56756 10948
rect 55804 10610 55860 10892
rect 56700 10834 56756 10892
rect 56700 10782 56702 10834
rect 56754 10782 56756 10834
rect 56700 10770 56756 10782
rect 56812 11170 56868 11182
rect 56812 11118 56814 11170
rect 56866 11118 56868 11170
rect 56812 11060 56868 11118
rect 55916 10724 55972 10734
rect 55916 10630 55972 10668
rect 55804 10558 55806 10610
rect 55858 10558 55860 10610
rect 55804 9940 55860 10558
rect 56812 10276 56868 11004
rect 56812 10210 56868 10220
rect 56924 10724 56980 11564
rect 55804 9874 55860 9884
rect 56924 9938 56980 10668
rect 57260 10052 57316 11788
rect 57820 11732 57876 11900
rect 58044 11890 58100 11900
rect 57372 11676 57876 11732
rect 57372 11506 57428 11676
rect 57372 11454 57374 11506
rect 57426 11454 57428 11506
rect 57372 11442 57428 11454
rect 57708 11396 57764 11406
rect 58380 11396 58436 11406
rect 57708 11394 58436 11396
rect 57708 11342 57710 11394
rect 57762 11342 58382 11394
rect 58434 11342 58436 11394
rect 57708 11340 58436 11342
rect 57708 11330 57764 11340
rect 58380 11330 58436 11340
rect 57932 11172 57988 11182
rect 57932 11170 58548 11172
rect 57932 11118 57934 11170
rect 57986 11118 58548 11170
rect 57932 11116 58548 11118
rect 57932 11106 57988 11116
rect 56924 9886 56926 9938
rect 56978 9886 56980 9938
rect 56924 9874 56980 9886
rect 57036 9996 57316 10052
rect 57932 10610 57988 10622
rect 57932 10558 57934 10610
rect 57986 10558 57988 10610
rect 55692 9324 56084 9380
rect 56028 9268 56084 9324
rect 56028 9266 56868 9268
rect 56028 9214 56030 9266
rect 56082 9214 56868 9266
rect 56028 9212 56868 9214
rect 56028 9202 56084 9212
rect 55244 8204 55412 8260
rect 55132 8036 55188 8092
rect 55244 8036 55300 8046
rect 55132 8034 55300 8036
rect 55132 7982 55246 8034
rect 55298 7982 55300 8034
rect 55132 7980 55300 7982
rect 55244 7970 55300 7980
rect 54684 7756 55300 7812
rect 54684 6914 54740 7756
rect 55244 7362 55300 7756
rect 55244 7310 55246 7362
rect 55298 7310 55300 7362
rect 55244 7298 55300 7310
rect 54684 6862 54686 6914
rect 54738 6862 54740 6914
rect 54684 6850 54740 6862
rect 55244 6580 55300 6590
rect 55020 5794 55076 5806
rect 55020 5742 55022 5794
rect 55074 5742 55076 5794
rect 55020 5682 55076 5742
rect 55020 5630 55022 5682
rect 55074 5630 55076 5682
rect 55020 5618 55076 5630
rect 54572 5346 55188 5348
rect 54572 5294 54574 5346
rect 54626 5294 55188 5346
rect 54572 5292 55188 5294
rect 54572 5282 54628 5292
rect 53004 5122 53060 5180
rect 53004 5070 53006 5122
rect 53058 5070 53060 5122
rect 53004 5058 53060 5070
rect 53564 5124 53620 5134
rect 53564 5030 53620 5068
rect 54236 5124 54292 5134
rect 54236 5030 54292 5068
rect 53340 4900 53396 4910
rect 53116 4898 53396 4900
rect 53116 4846 53342 4898
rect 53394 4846 53396 4898
rect 53116 4844 53396 4846
rect 53004 4452 53060 4462
rect 53116 4452 53172 4844
rect 53340 4834 53396 4844
rect 53004 4450 53172 4452
rect 53004 4398 53006 4450
rect 53058 4398 53172 4450
rect 53004 4396 53172 4398
rect 53004 4386 53060 4396
rect 55132 4226 55188 5292
rect 55244 5010 55300 6524
rect 55356 6132 55412 8204
rect 55804 8148 55860 8158
rect 55580 7586 55636 7598
rect 55580 7534 55582 7586
rect 55634 7534 55636 7586
rect 55468 6692 55524 6702
rect 55468 6598 55524 6636
rect 55580 6580 55636 7534
rect 55804 7474 55860 8092
rect 55804 7422 55806 7474
rect 55858 7422 55860 7474
rect 55804 7410 55860 7422
rect 56028 7476 56084 7486
rect 56028 6692 56084 7420
rect 56028 6598 56084 6636
rect 55580 6514 55636 6524
rect 55356 6038 55412 6076
rect 55692 6356 55748 6366
rect 55692 6130 55748 6300
rect 55692 6078 55694 6130
rect 55746 6078 55748 6130
rect 55244 4958 55246 5010
rect 55298 4958 55300 5010
rect 55244 4946 55300 4958
rect 55356 5682 55412 5694
rect 55356 5630 55358 5682
rect 55410 5630 55412 5682
rect 55356 5348 55412 5630
rect 55356 5122 55412 5292
rect 55356 5070 55358 5122
rect 55410 5070 55412 5122
rect 55356 4676 55412 5070
rect 55692 5124 55748 6078
rect 56028 6132 56084 6142
rect 56028 6018 56084 6076
rect 56028 5966 56030 6018
rect 56082 5966 56084 6018
rect 56028 5954 56084 5966
rect 56252 5460 56308 9212
rect 56812 9042 56868 9212
rect 56812 8990 56814 9042
rect 56866 8990 56868 9042
rect 56812 8978 56868 8990
rect 56700 8260 56756 8270
rect 56700 8166 56756 8204
rect 56588 6132 56644 6142
rect 56588 6038 56644 6076
rect 55692 5058 55748 5068
rect 55804 5404 56308 5460
rect 55356 4610 55412 4620
rect 55132 4174 55134 4226
rect 55186 4174 55188 4226
rect 55132 4162 55188 4174
rect 55804 4338 55860 5404
rect 56028 5236 56084 5246
rect 55916 5124 55972 5134
rect 55916 5030 55972 5068
rect 55804 4286 55806 4338
rect 55858 4286 55860 4338
rect 55804 3668 55860 4286
rect 56028 4450 56084 5180
rect 56252 5010 56308 5404
rect 56252 4958 56254 5010
rect 56306 4958 56308 5010
rect 56252 4946 56308 4958
rect 56924 5906 56980 5918
rect 56924 5854 56926 5906
rect 56978 5854 56980 5906
rect 56028 4398 56030 4450
rect 56082 4398 56084 4450
rect 56028 4340 56084 4398
rect 56924 4452 56980 5854
rect 56924 4386 56980 4396
rect 56588 4340 56644 4350
rect 56028 4338 56644 4340
rect 56028 4286 56590 4338
rect 56642 4286 56644 4338
rect 56028 4284 56644 4286
rect 56588 4274 56644 4284
rect 57036 4228 57092 9996
rect 57932 9940 57988 10558
rect 58492 10500 58548 11116
rect 58604 10836 58660 14476
rect 58828 14530 58884 14700
rect 58828 14478 58830 14530
rect 58882 14478 58884 14530
rect 58828 14466 58884 14478
rect 59164 14308 59220 15484
rect 59276 15428 59332 15438
rect 59276 15334 59332 15372
rect 59276 14756 59332 14766
rect 59276 14642 59332 14700
rect 59276 14590 59278 14642
rect 59330 14590 59332 14642
rect 59276 14578 59332 14590
rect 59500 14532 59556 15484
rect 59612 15202 59668 20300
rect 59724 20290 59780 20300
rect 59948 20018 60004 20030
rect 59948 19966 59950 20018
rect 60002 19966 60004 20018
rect 59948 18116 60004 19966
rect 60172 19236 60228 22428
rect 60508 22370 60564 22382
rect 60508 22318 60510 22370
rect 60562 22318 60564 22370
rect 60508 21812 60564 22318
rect 60844 22260 60900 22270
rect 60956 22260 61012 23102
rect 61292 23156 61348 23166
rect 61292 23062 61348 23100
rect 61852 22370 61908 23998
rect 62188 23268 62244 24670
rect 62300 24612 62356 26908
rect 62412 25620 62468 27132
rect 62748 27076 62804 27086
rect 62748 27074 63140 27076
rect 62748 27022 62750 27074
rect 62802 27022 63140 27074
rect 62748 27020 63140 27022
rect 62748 27010 62804 27020
rect 63084 26514 63140 27020
rect 63532 26908 63588 27580
rect 63084 26462 63086 26514
rect 63138 26462 63140 26514
rect 63084 26450 63140 26462
rect 63420 26852 63588 26908
rect 63308 26402 63364 26414
rect 63308 26350 63310 26402
rect 63362 26350 63364 26402
rect 63308 26292 63364 26350
rect 63420 26402 63476 26852
rect 63420 26350 63422 26402
rect 63474 26350 63476 26402
rect 63420 26338 63476 26350
rect 63308 26226 63364 26236
rect 62412 25554 62468 25564
rect 63084 25732 63140 25742
rect 62300 24546 62356 24556
rect 62748 24612 62804 24622
rect 62748 24518 62804 24556
rect 62524 23940 62580 23950
rect 62524 23938 63028 23940
rect 62524 23886 62526 23938
rect 62578 23886 63028 23938
rect 62524 23884 63028 23886
rect 62524 23874 62580 23884
rect 62972 23378 63028 23884
rect 62972 23326 62974 23378
rect 63026 23326 63028 23378
rect 62972 23314 63028 23326
rect 62300 23268 62356 23278
rect 62188 23212 62300 23268
rect 62300 23202 62356 23212
rect 61964 23156 62020 23166
rect 61964 23044 62020 23100
rect 62636 23156 62692 23166
rect 63084 23156 63140 25676
rect 63420 25508 63476 25518
rect 63420 25506 63812 25508
rect 63420 25454 63422 25506
rect 63474 25454 63812 25506
rect 63420 25452 63812 25454
rect 63420 25442 63476 25452
rect 63644 24724 63700 24734
rect 63644 24630 63700 24668
rect 63196 23268 63252 23278
rect 63196 23174 63252 23212
rect 62636 23062 62692 23100
rect 62972 23100 63140 23156
rect 63308 23156 63364 23166
rect 62188 23044 62244 23054
rect 61964 23042 62244 23044
rect 61964 22990 62190 23042
rect 62242 22990 62244 23042
rect 61964 22988 62244 22990
rect 62188 22978 62244 22988
rect 61852 22318 61854 22370
rect 61906 22318 61908 22370
rect 61852 22306 61908 22318
rect 62300 22594 62356 22606
rect 62300 22542 62302 22594
rect 62354 22542 62356 22594
rect 60844 22258 61012 22260
rect 60844 22206 60846 22258
rect 60898 22206 61012 22258
rect 60844 22204 61012 22206
rect 60844 22194 60900 22204
rect 60508 21746 60564 21756
rect 61068 22146 61124 22158
rect 61068 22094 61070 22146
rect 61122 22094 61124 22146
rect 60620 21476 60676 21486
rect 60956 21476 61012 21486
rect 60508 21364 60564 21374
rect 60508 20468 60564 21308
rect 60508 20402 60564 20412
rect 60620 20244 60676 21420
rect 60844 21474 61012 21476
rect 60844 21422 60958 21474
rect 61010 21422 61012 21474
rect 60844 21420 61012 21422
rect 60732 20692 60788 20702
rect 60844 20692 60900 21420
rect 60956 21410 61012 21420
rect 61068 20916 61124 22094
rect 62300 22148 62356 22542
rect 62300 22082 62356 22092
rect 61068 20850 61124 20860
rect 61404 20804 61460 20814
rect 62076 20804 62132 20814
rect 61404 20802 62132 20804
rect 61404 20750 61406 20802
rect 61458 20750 62078 20802
rect 62130 20750 62132 20802
rect 61404 20748 62132 20750
rect 61404 20738 61460 20748
rect 62076 20738 62132 20748
rect 62412 20804 62468 20814
rect 62412 20710 62468 20748
rect 62860 20804 62916 20814
rect 62860 20710 62916 20748
rect 60788 20636 60900 20692
rect 60732 20626 60788 20636
rect 60956 20580 61012 20590
rect 60956 20486 61012 20524
rect 61628 20580 61684 20590
rect 61628 20486 61684 20524
rect 62076 20468 62132 20478
rect 60620 20178 60676 20188
rect 61628 20244 61684 20254
rect 61180 20132 61236 20142
rect 61180 20038 61236 20076
rect 60844 20020 60900 20030
rect 60844 19926 60900 19964
rect 61068 19796 61124 19806
rect 61068 19346 61124 19740
rect 61068 19294 61070 19346
rect 61122 19294 61124 19346
rect 61068 19282 61124 19294
rect 60172 19170 60228 19180
rect 61404 19122 61460 19134
rect 61404 19070 61406 19122
rect 61458 19070 61460 19122
rect 60732 18562 60788 18574
rect 60732 18510 60734 18562
rect 60786 18510 60788 18562
rect 60508 18450 60564 18462
rect 60508 18398 60510 18450
rect 60562 18398 60564 18450
rect 59948 17106 60004 18060
rect 59948 17054 59950 17106
rect 60002 17054 60004 17106
rect 59948 17042 60004 17054
rect 60060 18338 60116 18350
rect 60060 18286 60062 18338
rect 60114 18286 60116 18338
rect 60060 18228 60116 18286
rect 60508 18340 60564 18398
rect 60732 18452 60788 18510
rect 61068 18508 61348 18564
rect 61068 18452 61124 18508
rect 60732 18396 61124 18452
rect 61180 18340 61236 18350
rect 60508 18338 61236 18340
rect 60508 18286 61182 18338
rect 61234 18286 61236 18338
rect 60508 18284 61236 18286
rect 61180 18274 61236 18284
rect 60060 17108 60116 18172
rect 60620 18116 60676 18126
rect 60620 17666 60676 18060
rect 61292 17778 61348 18508
rect 61404 18452 61460 19070
rect 61404 18386 61460 18396
rect 61292 17726 61294 17778
rect 61346 17726 61348 17778
rect 61292 17714 61348 17726
rect 61516 18226 61572 18238
rect 61516 18174 61518 18226
rect 61570 18174 61572 18226
rect 60620 17614 60622 17666
rect 60674 17614 60676 17666
rect 60620 17602 60676 17614
rect 60956 17668 61012 17678
rect 60060 17042 60116 17052
rect 59724 16884 59780 16894
rect 60172 16884 60228 16894
rect 59724 16882 60228 16884
rect 59724 16830 59726 16882
rect 59778 16830 60174 16882
rect 60226 16830 60228 16882
rect 59724 16828 60228 16830
rect 59724 16818 59780 16828
rect 59612 15150 59614 15202
rect 59666 15150 59668 15202
rect 59612 15138 59668 15150
rect 59724 15314 59780 15326
rect 59724 15262 59726 15314
rect 59778 15262 59780 15314
rect 59612 14532 59668 14542
rect 59500 14476 59612 14532
rect 59612 14438 59668 14476
rect 58940 14252 59220 14308
rect 59276 14308 59332 14346
rect 58828 13746 58884 13758
rect 58828 13694 58830 13746
rect 58882 13694 58884 13746
rect 58828 12292 58884 13694
rect 58828 12226 58884 12236
rect 58940 12180 58996 14252
rect 59276 14242 59332 14252
rect 59388 14308 59444 14318
rect 59388 14306 59556 14308
rect 59388 14254 59390 14306
rect 59442 14254 59556 14306
rect 59388 14252 59556 14254
rect 59388 14242 59444 14252
rect 59172 14140 59436 14150
rect 59228 14084 59276 14140
rect 59332 14084 59380 14140
rect 59172 14074 59436 14084
rect 59276 12964 59332 12974
rect 59500 12964 59556 14252
rect 59724 13970 59780 15262
rect 59836 15148 59892 16828
rect 60172 16818 60228 16828
rect 60844 16884 60900 16894
rect 60396 15652 60452 15662
rect 60284 15314 60340 15326
rect 60284 15262 60286 15314
rect 60338 15262 60340 15314
rect 59836 15092 60004 15148
rect 59724 13918 59726 13970
rect 59778 13918 59780 13970
rect 59724 13906 59780 13918
rect 59836 14418 59892 14430
rect 59836 14366 59838 14418
rect 59890 14366 59892 14418
rect 59276 12962 59556 12964
rect 59276 12910 59278 12962
rect 59330 12910 59556 12962
rect 59276 12908 59556 12910
rect 59276 12898 59332 12908
rect 59052 12738 59108 12750
rect 59052 12686 59054 12738
rect 59106 12686 59108 12738
rect 59052 12404 59108 12686
rect 59172 12572 59436 12582
rect 59228 12516 59276 12572
rect 59332 12516 59380 12572
rect 59172 12506 59436 12516
rect 59500 12516 59556 12908
rect 59724 13412 59780 13422
rect 59724 13074 59780 13356
rect 59724 13022 59726 13074
rect 59778 13022 59780 13074
rect 59724 12852 59780 13022
rect 59724 12786 59780 12796
rect 59500 12460 59780 12516
rect 59052 12338 59108 12348
rect 59388 12292 59444 12302
rect 59276 12236 59388 12292
rect 59052 12180 59108 12190
rect 58940 12178 59108 12180
rect 58940 12126 59054 12178
rect 59106 12126 59108 12178
rect 58940 12124 59108 12126
rect 59052 11508 59108 12124
rect 59052 11442 59108 11452
rect 58716 11394 58772 11406
rect 58716 11342 58718 11394
rect 58770 11342 58772 11394
rect 58716 11060 58772 11342
rect 59276 11172 59332 12236
rect 59388 12198 59444 12236
rect 58716 10994 58772 11004
rect 58828 11116 59332 11172
rect 59388 11394 59444 11406
rect 59388 11342 59390 11394
rect 59442 11342 59444 11394
rect 59388 11172 59444 11342
rect 59500 11284 59556 11294
rect 59500 11190 59556 11228
rect 58604 10780 58772 10836
rect 58604 10500 58660 10510
rect 58492 10498 58660 10500
rect 58492 10446 58606 10498
rect 58658 10446 58660 10498
rect 58492 10444 58660 10446
rect 58604 10434 58660 10444
rect 57708 9884 57932 9940
rect 57484 9604 57540 9614
rect 57484 9602 57652 9604
rect 57484 9550 57486 9602
rect 57538 9550 57652 9602
rect 57484 9548 57652 9550
rect 57484 9538 57540 9548
rect 57596 9154 57652 9548
rect 57596 9102 57598 9154
rect 57650 9102 57652 9154
rect 57596 9090 57652 9102
rect 57148 8148 57204 8158
rect 57148 8054 57204 8092
rect 57708 7140 57764 9884
rect 57932 9874 57988 9884
rect 57820 9714 57876 9726
rect 57820 9662 57822 9714
rect 57874 9662 57876 9714
rect 57820 8482 57876 9662
rect 57820 8430 57822 8482
rect 57874 8430 57876 8482
rect 57820 8418 57876 8430
rect 58380 8932 58436 8942
rect 58156 8372 58212 8382
rect 58156 8278 58212 8316
rect 58380 8260 58436 8876
rect 58716 8372 58772 10780
rect 58380 8146 58436 8204
rect 58380 8094 58382 8146
rect 58434 8094 58436 8146
rect 58380 8082 58436 8094
rect 58604 8316 58772 8372
rect 57484 7084 57764 7140
rect 57260 6692 57316 6702
rect 57260 6598 57316 6636
rect 57372 6580 57428 6590
rect 57148 6468 57204 6478
rect 57148 5236 57204 6412
rect 57372 6132 57428 6524
rect 57148 5122 57204 5180
rect 57148 5070 57150 5122
rect 57202 5070 57204 5122
rect 57148 5058 57204 5070
rect 57260 6076 57428 6132
rect 57260 5010 57316 6076
rect 57484 5908 57540 7084
rect 58268 6690 58324 6702
rect 58268 6638 58270 6690
rect 58322 6638 58324 6690
rect 58044 6580 58100 6590
rect 58044 6486 58100 6524
rect 57596 6468 57652 6478
rect 58268 6468 58324 6638
rect 57596 6466 57988 6468
rect 57596 6414 57598 6466
rect 57650 6414 57988 6466
rect 57596 6412 57988 6414
rect 57596 6402 57652 6412
rect 57932 6020 57988 6412
rect 58268 6244 58324 6412
rect 58268 6178 58324 6188
rect 58156 6020 58212 6030
rect 57932 6018 58212 6020
rect 57932 5966 58158 6018
rect 58210 5966 58212 6018
rect 57932 5964 58212 5966
rect 58156 5954 58212 5964
rect 57484 5814 57540 5852
rect 57820 5124 57876 5134
rect 57820 5030 57876 5068
rect 58156 5124 58212 5134
rect 58604 5124 58660 8316
rect 58716 8148 58772 8158
rect 58716 8054 58772 8092
rect 58828 6916 58884 11116
rect 59388 11106 59444 11116
rect 59172 11004 59436 11014
rect 59228 10948 59276 11004
rect 59332 10948 59380 11004
rect 59172 10938 59436 10948
rect 59172 9436 59436 9446
rect 59228 9380 59276 9436
rect 59332 9380 59380 9436
rect 59172 9370 59436 9380
rect 59724 8930 59780 12460
rect 59836 12292 59892 14366
rect 59836 12226 59892 12236
rect 59724 8878 59726 8930
rect 59778 8878 59780 8930
rect 59724 8372 59780 8878
rect 59724 8306 59780 8316
rect 59836 8596 59892 8606
rect 59172 7868 59436 7878
rect 59228 7812 59276 7868
rect 59332 7812 59380 7868
rect 59172 7802 59436 7812
rect 59500 6916 59556 6926
rect 58828 6914 59556 6916
rect 58828 6862 58830 6914
rect 58882 6862 59502 6914
rect 59554 6862 59556 6914
rect 58828 6860 59556 6862
rect 58828 6850 58884 6860
rect 59500 6850 59556 6860
rect 59164 6692 59220 6702
rect 59164 6598 59220 6636
rect 59724 6468 59780 6478
rect 59724 6374 59780 6412
rect 59172 6300 59436 6310
rect 59228 6244 59276 6300
rect 59332 6244 59380 6300
rect 59172 6234 59436 6244
rect 59836 5460 59892 8540
rect 59948 6020 60004 15092
rect 60172 12404 60228 12414
rect 60284 12404 60340 15262
rect 60172 12402 60340 12404
rect 60172 12350 60174 12402
rect 60226 12350 60340 12402
rect 60172 12348 60340 12350
rect 60396 15316 60452 15596
rect 60396 12404 60452 15260
rect 60732 14868 60788 14878
rect 60732 13860 60788 14812
rect 60732 13766 60788 13804
rect 60172 12338 60228 12348
rect 60396 12310 60452 12348
rect 60844 12962 60900 16828
rect 60956 16770 61012 17612
rect 61516 17556 61572 18174
rect 61516 17490 61572 17500
rect 60956 16718 60958 16770
rect 61010 16718 61012 16770
rect 60956 16706 61012 16718
rect 61628 15148 61684 20188
rect 61852 19796 61908 19806
rect 61852 19460 61908 19740
rect 61852 19234 61908 19404
rect 61852 19182 61854 19234
rect 61906 19182 61908 19234
rect 61852 19170 61908 19182
rect 61964 18450 62020 18462
rect 61964 18398 61966 18450
rect 62018 18398 62020 18450
rect 61964 18228 62020 18398
rect 61964 18162 62020 18172
rect 60844 12910 60846 12962
rect 60898 12910 60900 12962
rect 60396 12180 60452 12190
rect 60396 11284 60452 12124
rect 60732 11508 60788 11518
rect 60732 11414 60788 11452
rect 60396 10500 60452 11228
rect 60732 10500 60788 10510
rect 60396 10498 60788 10500
rect 60396 10446 60734 10498
rect 60786 10446 60788 10498
rect 60396 10444 60788 10446
rect 60732 10434 60788 10444
rect 60844 9604 60900 12910
rect 60732 9548 60900 9604
rect 60956 15092 61684 15148
rect 60620 8596 60676 8606
rect 60060 6916 60116 6926
rect 60060 6914 60340 6916
rect 60060 6862 60062 6914
rect 60114 6862 60340 6914
rect 60060 6860 60340 6862
rect 60060 6850 60116 6860
rect 59948 5954 60004 5964
rect 60284 5794 60340 6860
rect 60620 6466 60676 8540
rect 60620 6414 60622 6466
rect 60674 6414 60676 6466
rect 60284 5742 60286 5794
rect 60338 5742 60340 5794
rect 60284 5730 60340 5742
rect 60508 5908 60564 5918
rect 59388 5236 59444 5246
rect 59836 5236 59892 5404
rect 59948 5236 60004 5246
rect 59836 5234 60004 5236
rect 59836 5182 59950 5234
rect 60002 5182 60004 5234
rect 59836 5180 60004 5182
rect 59388 5142 59444 5180
rect 59948 5170 60004 5180
rect 58828 5124 58884 5134
rect 58604 5068 58772 5124
rect 58156 5030 58212 5068
rect 57260 4958 57262 5010
rect 57314 4958 57316 5010
rect 57260 4946 57316 4958
rect 58716 5012 58772 5068
rect 58828 5030 58884 5068
rect 58716 4946 58772 4956
rect 59500 5012 59556 5022
rect 58604 4900 58660 4910
rect 57596 4898 58660 4900
rect 57596 4846 58606 4898
rect 58658 4846 58660 4898
rect 57596 4844 58660 4846
rect 57596 4564 57652 4844
rect 58604 4834 58660 4844
rect 59172 4732 59436 4742
rect 59228 4676 59276 4732
rect 59332 4676 59380 4732
rect 59172 4666 59436 4676
rect 57372 4508 57652 4564
rect 57372 4450 57428 4508
rect 57372 4398 57374 4450
rect 57426 4398 57428 4450
rect 57372 4386 57428 4398
rect 55804 3602 55860 3612
rect 56924 4172 57092 4228
rect 59500 4226 59556 4956
rect 60508 5010 60564 5852
rect 60620 5796 60676 6414
rect 60620 5730 60676 5740
rect 60732 5236 60788 9548
rect 60844 8932 60900 8942
rect 60844 8838 60900 8876
rect 60844 5906 60900 5918
rect 60844 5854 60846 5906
rect 60898 5854 60900 5906
rect 60844 5796 60900 5854
rect 60844 5730 60900 5740
rect 60732 5122 60788 5180
rect 60732 5070 60734 5122
rect 60786 5070 60788 5122
rect 60732 5058 60788 5070
rect 60508 4958 60510 5010
rect 60562 4958 60564 5010
rect 60508 4340 60564 4958
rect 60620 4340 60676 4350
rect 60508 4338 60676 4340
rect 60508 4286 60622 4338
rect 60674 4286 60676 4338
rect 60508 4284 60676 4286
rect 60620 4274 60676 4284
rect 59500 4174 59502 4226
rect 59554 4174 59556 4226
rect 52556 3442 52836 3444
rect 52556 3390 52558 3442
rect 52610 3390 52836 3442
rect 52556 3388 52836 3390
rect 56028 3444 56084 3482
rect 56252 3444 56308 3454
rect 56028 3442 56308 3444
rect 56028 3390 56030 3442
rect 56082 3390 56254 3442
rect 56306 3390 56308 3442
rect 56028 3388 56308 3390
rect 52556 3378 52612 3388
rect 56028 800 56084 3388
rect 56252 3378 56308 3388
rect 56588 3444 56644 3454
rect 56924 3444 56980 4172
rect 59500 4162 59556 4174
rect 57036 3668 57092 3678
rect 57036 3574 57092 3612
rect 56588 3442 56980 3444
rect 56588 3390 56590 3442
rect 56642 3390 56980 3442
rect 56588 3388 56980 3390
rect 60060 3444 60116 3482
rect 60284 3444 60340 3454
rect 60060 3442 60340 3444
rect 60060 3390 60062 3442
rect 60114 3390 60286 3442
rect 60338 3390 60340 3442
rect 60060 3388 60340 3390
rect 56588 3378 56644 3388
rect 59172 3164 59436 3174
rect 59228 3108 59276 3164
rect 59332 3108 59380 3164
rect 59172 3098 59436 3108
rect 60060 800 60116 3388
rect 60284 3378 60340 3388
rect 60620 3444 60676 3454
rect 60956 3444 61012 15092
rect 61292 14420 61348 14430
rect 61292 13746 61348 14364
rect 61964 13860 62020 13870
rect 61292 13694 61294 13746
rect 61346 13694 61348 13746
rect 61292 13682 61348 13694
rect 61628 13858 62020 13860
rect 61628 13806 61966 13858
rect 62018 13806 62020 13858
rect 61628 13804 62020 13806
rect 61628 13074 61684 13804
rect 61964 13794 62020 13804
rect 61628 13022 61630 13074
rect 61682 13022 61684 13074
rect 61628 13010 61684 13022
rect 61068 12404 61124 12414
rect 61068 12310 61124 12348
rect 61740 12404 61796 12414
rect 61740 12310 61796 12348
rect 62076 12180 62132 20412
rect 62188 20020 62244 20030
rect 62188 19796 62244 19964
rect 62300 19796 62356 19806
rect 62188 19740 62300 19796
rect 62188 18562 62244 19740
rect 62300 19730 62356 19740
rect 62188 18510 62190 18562
rect 62242 18510 62244 18562
rect 62188 18498 62244 18510
rect 62300 19572 62356 19582
rect 62188 13746 62244 13758
rect 62188 13694 62190 13746
rect 62242 13694 62244 13746
rect 62188 12404 62244 13694
rect 62188 12338 62244 12348
rect 61516 12178 62132 12180
rect 61516 12126 62078 12178
rect 62130 12126 62132 12178
rect 61516 12124 62132 12126
rect 61516 11508 61572 12124
rect 62076 12114 62132 12124
rect 61292 11506 61572 11508
rect 61292 11454 61518 11506
rect 61570 11454 61572 11506
rect 61292 11452 61572 11454
rect 61068 11172 61124 11182
rect 61068 11078 61124 11116
rect 61068 9940 61124 9950
rect 61068 9826 61124 9884
rect 61068 9774 61070 9826
rect 61122 9774 61124 9826
rect 61068 9762 61124 9774
rect 61292 9268 61348 11452
rect 61516 11442 61572 11452
rect 61740 10722 61796 10734
rect 61740 10670 61742 10722
rect 61794 10670 61796 10722
rect 61740 9940 61796 10670
rect 61964 10610 62020 10622
rect 61964 10558 61966 10610
rect 62018 10558 62020 10610
rect 61852 9940 61908 9950
rect 61740 9938 61908 9940
rect 61740 9886 61854 9938
rect 61906 9886 61908 9938
rect 61740 9884 61908 9886
rect 61852 9874 61908 9884
rect 61292 9174 61348 9212
rect 61964 9266 62020 10558
rect 61964 9214 61966 9266
rect 62018 9214 62020 9266
rect 61964 9202 62020 9214
rect 62300 9268 62356 19516
rect 62412 18452 62468 18462
rect 62412 17780 62468 18396
rect 62860 18452 62916 18462
rect 62860 18358 62916 18396
rect 62412 12290 62468 17724
rect 62860 15876 62916 15886
rect 62412 12238 62414 12290
rect 62466 12238 62468 12290
rect 62412 12068 62468 12238
rect 62412 12002 62468 12012
rect 62748 14420 62804 14430
rect 62300 9212 62468 9268
rect 62300 9044 62356 9054
rect 62300 8950 62356 8988
rect 61964 6916 62020 6926
rect 61964 6802 62020 6860
rect 61964 6750 61966 6802
rect 62018 6750 62020 6802
rect 61964 6738 62020 6750
rect 61740 6466 61796 6478
rect 61740 6414 61742 6466
rect 61794 6414 61796 6466
rect 61740 6244 61796 6414
rect 61292 6188 61740 6244
rect 61180 5124 61236 5134
rect 61292 5124 61348 6188
rect 61740 6178 61796 6188
rect 61740 6020 61796 6030
rect 61516 6018 61796 6020
rect 61516 5966 61742 6018
rect 61794 5966 61796 6018
rect 61516 5964 61796 5966
rect 61236 5068 61348 5124
rect 61404 5794 61460 5806
rect 61404 5742 61406 5794
rect 61458 5742 61460 5794
rect 61404 5348 61460 5742
rect 61404 5124 61460 5292
rect 61180 5030 61236 5068
rect 61404 5058 61460 5068
rect 61404 4452 61460 4462
rect 61516 4452 61572 5964
rect 61740 5954 61796 5964
rect 62076 5908 62132 5918
rect 62076 5906 62244 5908
rect 62076 5854 62078 5906
rect 62130 5854 62244 5906
rect 62076 5852 62244 5854
rect 62076 5842 62132 5852
rect 61628 5460 61684 5470
rect 61628 5122 61684 5404
rect 62188 5346 62244 5852
rect 62188 5294 62190 5346
rect 62242 5294 62244 5346
rect 62188 5282 62244 5294
rect 61628 5070 61630 5122
rect 61682 5070 61684 5122
rect 61628 5058 61684 5070
rect 61404 4450 61572 4452
rect 61404 4398 61406 4450
rect 61458 4398 61572 4450
rect 61404 4396 61572 4398
rect 61404 4386 61460 4396
rect 62412 3668 62468 9212
rect 62524 9156 62580 9166
rect 62524 9062 62580 9100
rect 62636 7474 62692 7486
rect 62636 7422 62638 7474
rect 62690 7422 62692 7474
rect 62636 6130 62692 7422
rect 62636 6078 62638 6130
rect 62690 6078 62692 6130
rect 62636 6066 62692 6078
rect 62748 5908 62804 14364
rect 62860 13860 62916 15820
rect 62972 15428 63028 23100
rect 63308 23062 63364 23100
rect 63756 23044 63812 25452
rect 64092 25396 64148 25406
rect 63868 25394 64148 25396
rect 63868 25342 64094 25394
rect 64146 25342 64148 25394
rect 63868 25340 64148 25342
rect 63868 24946 63924 25340
rect 64092 25330 64148 25340
rect 63868 24894 63870 24946
rect 63922 24894 63924 24946
rect 63868 24882 63924 24894
rect 64204 23714 64260 23726
rect 64204 23662 64206 23714
rect 64258 23662 64260 23714
rect 64204 23604 64260 23662
rect 64204 23538 64260 23548
rect 63756 22596 63812 22988
rect 63756 22540 63924 22596
rect 63084 22372 63140 22382
rect 63084 22278 63140 22316
rect 63868 21812 63924 22540
rect 64428 22036 64484 32396
rect 64652 31892 64708 31902
rect 64540 31836 64652 31892
rect 64540 29988 64596 31836
rect 64652 31826 64708 31836
rect 64764 30996 64820 34076
rect 65100 34130 65156 34142
rect 65100 34078 65102 34130
rect 65154 34078 65156 34130
rect 65100 33572 65156 34078
rect 65660 34132 65716 34142
rect 65660 34038 65716 34076
rect 65100 33506 65156 33516
rect 66444 33572 66500 33582
rect 66444 33478 66500 33516
rect 66780 33348 66836 33358
rect 65996 33124 66052 33134
rect 65996 31948 66052 33068
rect 66668 32562 66724 32574
rect 66668 32510 66670 32562
rect 66722 32510 66724 32562
rect 66220 32452 66276 32462
rect 66220 32358 66276 32396
rect 66668 32452 66724 32510
rect 66668 32386 66724 32396
rect 64876 31892 64932 31902
rect 64876 31666 64932 31836
rect 65772 31892 66052 31948
rect 64876 31614 64878 31666
rect 64930 31614 64932 31666
rect 64876 31602 64932 31614
rect 65212 31666 65268 31678
rect 65212 31614 65214 31666
rect 65266 31614 65268 31666
rect 64652 30994 64820 30996
rect 64652 30942 64766 30994
rect 64818 30942 64820 30994
rect 64652 30940 64820 30942
rect 64652 30210 64708 30940
rect 64764 30930 64820 30940
rect 65212 31556 65268 31614
rect 64652 30158 64654 30210
rect 64706 30158 64708 30210
rect 64652 30100 64708 30158
rect 64652 30044 65156 30100
rect 64540 29932 64820 29988
rect 64764 29538 64820 29932
rect 64764 29486 64766 29538
rect 64818 29486 64820 29538
rect 64764 29474 64820 29486
rect 64988 29652 65044 29662
rect 64876 26290 64932 26302
rect 64876 26238 64878 26290
rect 64930 26238 64932 26290
rect 64540 26180 64596 26190
rect 64876 26180 64932 26238
rect 64540 26178 64932 26180
rect 64540 26126 64542 26178
rect 64594 26126 64932 26178
rect 64540 26124 64932 26126
rect 64540 25956 64596 26124
rect 64540 25890 64596 25900
rect 64764 25172 64820 25182
rect 64764 24052 64820 25116
rect 64876 24724 64932 24734
rect 64876 24630 64932 24668
rect 64764 23958 64820 23996
rect 64876 22930 64932 22942
rect 64876 22878 64878 22930
rect 64930 22878 64932 22930
rect 64876 22596 64932 22878
rect 64428 21980 64708 22036
rect 64540 21812 64596 21822
rect 63868 21810 64596 21812
rect 63868 21758 64542 21810
rect 64594 21758 64596 21810
rect 63868 21756 64596 21758
rect 63868 21586 63924 21756
rect 63868 21534 63870 21586
rect 63922 21534 63924 21586
rect 63868 21522 63924 21534
rect 63084 21474 63140 21486
rect 63084 21422 63086 21474
rect 63138 21422 63140 21474
rect 63084 20580 63140 21422
rect 63756 20802 63812 20814
rect 63756 20750 63758 20802
rect 63810 20750 63812 20802
rect 63084 20514 63140 20524
rect 63196 20690 63252 20702
rect 63196 20638 63198 20690
rect 63250 20638 63252 20690
rect 63196 19796 63252 20638
rect 63196 19730 63252 19740
rect 63308 20356 63364 20366
rect 63084 18562 63140 18574
rect 63084 18510 63086 18562
rect 63138 18510 63140 18562
rect 63084 16994 63140 18510
rect 63308 17444 63364 20300
rect 63756 20132 63812 20750
rect 64428 20802 64484 21756
rect 64540 21746 64596 21756
rect 64428 20750 64430 20802
rect 64482 20750 64484 20802
rect 64428 20738 64484 20750
rect 63980 20692 64036 20702
rect 64316 20692 64372 20702
rect 63980 20690 64316 20692
rect 63980 20638 63982 20690
rect 64034 20638 64316 20690
rect 63980 20636 64316 20638
rect 63980 20626 64036 20636
rect 64316 20626 64372 20636
rect 63756 20066 63812 20076
rect 64540 20132 64596 20142
rect 64540 20038 64596 20076
rect 63868 19906 63924 19918
rect 63868 19854 63870 19906
rect 63922 19854 63924 19906
rect 63868 19684 63924 19854
rect 63868 19618 63924 19628
rect 63868 18452 63924 18462
rect 63532 18340 63588 18350
rect 63420 17778 63476 17790
rect 63420 17726 63422 17778
rect 63474 17726 63476 17778
rect 63420 17556 63476 17726
rect 63420 17490 63476 17500
rect 63308 17378 63364 17388
rect 63084 16942 63086 16994
rect 63138 16942 63140 16994
rect 63084 16930 63140 16942
rect 63532 16660 63588 18284
rect 63868 17890 63924 18396
rect 63868 17838 63870 17890
rect 63922 17838 63924 17890
rect 63868 17826 63924 17838
rect 64652 18340 64708 21980
rect 64876 21698 64932 22540
rect 64876 21646 64878 21698
rect 64930 21646 64932 21698
rect 64876 21634 64932 21646
rect 64988 20132 65044 29596
rect 65100 29650 65156 30044
rect 65100 29598 65102 29650
rect 65154 29598 65156 29650
rect 65100 29586 65156 29598
rect 65212 29428 65268 31500
rect 65548 31554 65604 31566
rect 65548 31502 65550 31554
rect 65602 31502 65604 31554
rect 65436 31108 65492 31118
rect 65548 31108 65604 31502
rect 65436 31106 65604 31108
rect 65436 31054 65438 31106
rect 65490 31054 65604 31106
rect 65436 31052 65604 31054
rect 65436 31042 65492 31052
rect 65324 30098 65380 30110
rect 65324 30046 65326 30098
rect 65378 30046 65380 30098
rect 65324 29652 65380 30046
rect 65436 29652 65492 29662
rect 65324 29650 65492 29652
rect 65324 29598 65438 29650
rect 65490 29598 65492 29650
rect 65324 29596 65492 29598
rect 65436 29586 65492 29596
rect 65772 29652 65828 31892
rect 65884 31668 65940 31678
rect 65884 31666 66276 31668
rect 65884 31614 65886 31666
rect 65938 31614 66276 31666
rect 65884 31612 66276 31614
rect 65884 31602 65940 31612
rect 66220 29988 66276 31612
rect 66332 31556 66388 31566
rect 66332 31462 66388 31500
rect 66668 30212 66724 30222
rect 66556 29988 66612 29998
rect 66220 29932 66388 29988
rect 65772 29586 65828 29596
rect 65100 29372 65268 29428
rect 65772 29428 65828 29438
rect 66220 29428 66276 29438
rect 65772 29426 66276 29428
rect 65772 29374 65774 29426
rect 65826 29374 66222 29426
rect 66274 29374 66276 29426
rect 65772 29372 66276 29374
rect 65100 23378 65156 29372
rect 65772 29362 65828 29372
rect 66220 29362 66276 29372
rect 65212 29204 65268 29214
rect 65212 26290 65268 29148
rect 66332 28866 66388 29932
rect 66556 29204 66612 29932
rect 66556 29110 66612 29148
rect 66332 28814 66334 28866
rect 66386 28814 66388 28866
rect 66332 28802 66388 28814
rect 66668 28866 66724 30156
rect 66668 28814 66670 28866
rect 66722 28814 66724 28866
rect 65884 28644 65940 28654
rect 65324 26964 65380 26974
rect 65884 26908 65940 28588
rect 66220 27300 66276 27310
rect 66220 27206 66276 27244
rect 66332 27074 66388 27086
rect 66332 27022 66334 27074
rect 66386 27022 66388 27074
rect 66332 26908 66388 27022
rect 65324 26514 65380 26908
rect 65324 26462 65326 26514
rect 65378 26462 65380 26514
rect 65324 26450 65380 26462
rect 65772 26852 65940 26908
rect 66108 26852 66388 26908
rect 66556 26964 66612 26974
rect 66556 26870 66612 26908
rect 65436 26404 65492 26414
rect 65436 26310 65492 26348
rect 65212 26238 65214 26290
rect 65266 26238 65268 26290
rect 65212 26226 65268 26238
rect 65212 25508 65268 25518
rect 65212 24722 65268 25452
rect 65212 24670 65214 24722
rect 65266 24670 65268 24722
rect 65212 24658 65268 24670
rect 65436 24834 65492 24846
rect 65436 24782 65438 24834
rect 65490 24782 65492 24834
rect 65436 23604 65492 24782
rect 65772 23716 65828 26852
rect 66108 26514 66164 26852
rect 66108 26462 66110 26514
rect 66162 26462 66164 26514
rect 66108 26450 66164 26462
rect 65884 26290 65940 26302
rect 65884 26238 65886 26290
rect 65938 26238 65940 26290
rect 65884 23828 65940 26238
rect 65996 26290 66052 26302
rect 65996 26238 65998 26290
rect 66050 26238 66052 26290
rect 65996 25396 66052 26238
rect 66220 26290 66276 26302
rect 66220 26238 66222 26290
rect 66274 26238 66276 26290
rect 66220 25844 66276 26238
rect 66444 26292 66500 26302
rect 66668 26292 66724 28814
rect 66780 26516 66836 33292
rect 67676 33348 67732 34974
rect 67676 33282 67732 33292
rect 67004 33234 67060 33246
rect 67340 33236 67396 33246
rect 67004 33182 67006 33234
rect 67058 33182 67060 33234
rect 67004 33124 67060 33182
rect 67004 33058 67060 33068
rect 67116 33234 67396 33236
rect 67116 33182 67342 33234
rect 67394 33182 67396 33234
rect 67116 33180 67396 33182
rect 66892 32676 66948 32686
rect 67116 32676 67172 33180
rect 67340 33170 67396 33180
rect 67788 32786 67844 35252
rect 68124 35140 68180 39200
rect 68832 36876 69096 36886
rect 68888 36820 68936 36876
rect 68992 36820 69040 36876
rect 68832 36810 69096 36820
rect 68348 36708 68404 36718
rect 70588 36708 70644 39200
rect 71820 36708 71876 36718
rect 70588 36706 71876 36708
rect 70588 36654 71822 36706
rect 71874 36654 71876 36706
rect 70588 36652 71876 36654
rect 68348 35698 68404 36652
rect 71820 36642 71876 36652
rect 73052 36708 73108 39200
rect 73948 38388 74004 38398
rect 73052 36642 73108 36652
rect 73724 36932 73780 36942
rect 70812 36482 70868 36494
rect 70812 36430 70814 36482
rect 70866 36430 70868 36482
rect 70476 36260 70532 36270
rect 70476 36166 70532 36204
rect 70812 36260 70868 36430
rect 70812 36194 70868 36204
rect 72380 36372 72436 36382
rect 68348 35646 68350 35698
rect 68402 35646 68404 35698
rect 68348 35308 68404 35646
rect 71260 35810 71316 35822
rect 71260 35758 71262 35810
rect 71314 35758 71316 35810
rect 69356 35586 69412 35598
rect 69356 35534 69358 35586
rect 69410 35534 69412 35586
rect 68832 35308 69096 35318
rect 68348 35252 68628 35308
rect 68124 35074 68180 35084
rect 68572 35026 68628 35252
rect 68888 35252 68936 35308
rect 68992 35252 69040 35308
rect 68832 35242 69096 35252
rect 69356 35140 69412 35534
rect 71260 35308 71316 35758
rect 69356 35074 69412 35084
rect 70700 35252 71316 35308
rect 71596 35698 71652 35710
rect 71596 35646 71598 35698
rect 71650 35646 71652 35698
rect 68572 34974 68574 35026
rect 68626 34974 68628 35026
rect 68572 34962 68628 34974
rect 70140 34914 70196 34926
rect 70140 34862 70142 34914
rect 70194 34862 70196 34914
rect 70028 34244 70084 34254
rect 70028 34150 70084 34188
rect 69692 34132 69748 34142
rect 69692 34038 69748 34076
rect 68572 34020 68628 34030
rect 67788 32734 67790 32786
rect 67842 32734 67844 32786
rect 67788 32722 67844 32734
rect 67900 34018 68628 34020
rect 67900 33966 68574 34018
rect 68626 33966 68628 34018
rect 67900 33964 68628 33966
rect 66892 32674 67284 32676
rect 66892 32622 66894 32674
rect 66946 32622 67284 32674
rect 66892 32620 67284 32622
rect 66892 32610 66948 32620
rect 67228 29876 67284 32620
rect 67452 32564 67508 32574
rect 67900 32564 67956 33964
rect 68572 33954 68628 33964
rect 69356 34020 69412 34030
rect 68832 33740 69096 33750
rect 68888 33684 68936 33740
rect 68992 33684 69040 33740
rect 68832 33674 69096 33684
rect 69356 33124 69412 33964
rect 70140 33908 70196 34862
rect 70476 34132 70532 34142
rect 70476 34038 70532 34076
rect 70028 33852 70196 33908
rect 70028 33346 70084 33852
rect 70700 33460 70756 35252
rect 70924 34802 70980 34814
rect 70924 34750 70926 34802
rect 70978 34750 70980 34802
rect 70924 34468 70980 34750
rect 70924 34402 70980 34412
rect 71036 34242 71092 34254
rect 71036 34190 71038 34242
rect 71090 34190 71092 34242
rect 70812 34132 70868 34142
rect 70812 34038 70868 34076
rect 71036 34020 71092 34190
rect 71036 33954 71092 33964
rect 71372 34242 71428 34254
rect 71372 34190 71374 34242
rect 71426 34190 71428 34242
rect 70812 33460 70868 33470
rect 70700 33458 70868 33460
rect 70700 33406 70814 33458
rect 70866 33406 70868 33458
rect 70700 33404 70868 33406
rect 70812 33394 70868 33404
rect 70028 33294 70030 33346
rect 70082 33294 70084 33346
rect 69356 33058 69412 33068
rect 69692 33124 69748 33134
rect 67452 32562 67956 32564
rect 67452 32510 67454 32562
rect 67506 32510 67956 32562
rect 67452 32508 67956 32510
rect 67452 32498 67508 32508
rect 67564 30882 67620 30894
rect 67564 30830 67566 30882
rect 67618 30830 67620 30882
rect 67564 30212 67620 30830
rect 67564 30146 67620 30156
rect 67564 29988 67620 29998
rect 67564 29894 67620 29932
rect 66892 29538 66948 29550
rect 66892 29486 66894 29538
rect 66946 29486 66948 29538
rect 66892 29316 66948 29486
rect 66892 26908 66948 29260
rect 67228 29538 67284 29820
rect 67228 29486 67230 29538
rect 67282 29486 67284 29538
rect 67116 28644 67172 28654
rect 67116 28550 67172 28588
rect 67228 28530 67284 29486
rect 67228 28478 67230 28530
rect 67282 28478 67284 28530
rect 67228 28466 67284 28478
rect 67004 27748 67060 27758
rect 67004 27074 67060 27692
rect 67564 27076 67620 27086
rect 67004 27022 67006 27074
rect 67058 27022 67060 27074
rect 67004 27010 67060 27022
rect 67452 27074 67620 27076
rect 67452 27022 67566 27074
rect 67618 27022 67620 27074
rect 67452 27020 67620 27022
rect 66892 26852 67060 26908
rect 66780 26460 66948 26516
rect 66780 26292 66836 26302
rect 66444 26290 66836 26292
rect 66444 26238 66446 26290
rect 66498 26238 66782 26290
rect 66834 26238 66836 26290
rect 66444 26236 66836 26238
rect 66444 26226 66500 26236
rect 66780 26226 66836 26236
rect 66220 25788 66612 25844
rect 66220 25618 66276 25630
rect 66220 25566 66222 25618
rect 66274 25566 66276 25618
rect 66220 25508 66276 25566
rect 66220 25442 66276 25452
rect 65996 25330 66052 25340
rect 65996 25172 66052 25182
rect 65996 24834 66052 25116
rect 65996 24782 65998 24834
rect 66050 24782 66052 24834
rect 65996 24770 66052 24782
rect 65884 23772 66388 23828
rect 65772 23660 65940 23716
rect 65492 23548 65828 23604
rect 65436 23538 65492 23548
rect 65100 23326 65102 23378
rect 65154 23326 65156 23378
rect 65100 22930 65156 23326
rect 65660 23380 65716 23390
rect 65100 22878 65102 22930
rect 65154 22878 65156 22930
rect 65100 22866 65156 22878
rect 65548 23268 65604 23278
rect 65100 22372 65156 22382
rect 65100 22370 65268 22372
rect 65100 22318 65102 22370
rect 65154 22318 65268 22370
rect 65100 22316 65268 22318
rect 65100 22306 65156 22316
rect 65100 20692 65156 20702
rect 65100 20598 65156 20636
rect 65100 20132 65156 20142
rect 64988 20130 65156 20132
rect 64988 20078 65102 20130
rect 65154 20078 65156 20130
rect 64988 20076 65156 20078
rect 64876 20020 64932 20030
rect 64876 19926 64932 19964
rect 64988 19684 65044 20076
rect 65100 20066 65156 20076
rect 64988 19618 65044 19628
rect 65212 19012 65268 22316
rect 65324 22370 65380 22382
rect 65324 22318 65326 22370
rect 65378 22318 65380 22370
rect 65324 21810 65380 22318
rect 65324 21758 65326 21810
rect 65378 21758 65380 21810
rect 65324 21746 65380 21758
rect 65548 21698 65604 23212
rect 65660 22932 65716 23324
rect 65660 22866 65716 22876
rect 65772 22484 65828 23548
rect 65772 22390 65828 22428
rect 65548 21646 65550 21698
rect 65602 21646 65604 21698
rect 65548 21634 65604 21646
rect 65324 21588 65380 21598
rect 65324 21494 65380 21532
rect 65548 20132 65604 20142
rect 65212 18946 65268 18956
rect 65436 20130 65604 20132
rect 65436 20078 65550 20130
rect 65602 20078 65604 20130
rect 65436 20076 65604 20078
rect 65436 19796 65492 20076
rect 65548 20066 65604 20076
rect 65324 18450 65380 18462
rect 65324 18398 65326 18450
rect 65378 18398 65380 18450
rect 64988 18340 65044 18350
rect 65324 18340 65380 18398
rect 64204 17668 64260 17678
rect 64204 17574 64260 17612
rect 64652 17666 64708 18284
rect 64652 17614 64654 17666
rect 64706 17614 64708 17666
rect 64652 17602 64708 17614
rect 64876 18338 65380 18340
rect 64876 18286 64990 18338
rect 65042 18286 65380 18338
rect 64876 18284 65380 18286
rect 63532 16594 63588 16604
rect 63644 17444 63700 17454
rect 62972 15362 63028 15372
rect 63308 15764 63364 15774
rect 63308 15204 63364 15708
rect 63308 13970 63364 15148
rect 63532 14868 63588 14878
rect 63532 14306 63588 14812
rect 63532 14254 63534 14306
rect 63586 14254 63588 14306
rect 63532 14196 63588 14254
rect 63532 14130 63588 14140
rect 63644 14532 63700 17388
rect 63868 16884 63924 16894
rect 63868 16790 63924 16828
rect 64876 16772 64932 18284
rect 64988 18274 65044 18284
rect 65324 18228 65380 18284
rect 65324 18162 65380 18172
rect 64988 17556 65044 17566
rect 65436 17556 65492 19740
rect 65660 18564 65716 18574
rect 65660 18338 65716 18508
rect 65660 18286 65662 18338
rect 65714 18286 65716 18338
rect 65660 18274 65716 18286
rect 65884 18340 65940 23660
rect 66220 23604 66276 23614
rect 65996 23154 66052 23166
rect 65996 23102 65998 23154
rect 66050 23102 66052 23154
rect 65996 23044 66052 23102
rect 65996 22978 66052 22988
rect 66220 22820 66276 23548
rect 65884 18274 65940 18284
rect 65996 22764 66276 22820
rect 65996 18116 66052 22764
rect 66220 21812 66276 21822
rect 66220 21698 66276 21756
rect 66220 21646 66222 21698
rect 66274 21646 66276 21698
rect 66220 21634 66276 21646
rect 65884 18060 66052 18116
rect 66108 20018 66164 20030
rect 66108 19966 66110 20018
rect 66162 19966 66164 20018
rect 65548 17668 65604 17678
rect 65548 17666 65828 17668
rect 65548 17614 65550 17666
rect 65602 17614 65828 17666
rect 65548 17612 65828 17614
rect 65548 17602 65604 17612
rect 64988 17554 65492 17556
rect 64988 17502 64990 17554
rect 65042 17502 65492 17554
rect 64988 17500 65492 17502
rect 64988 17490 65044 17500
rect 64876 16706 64932 16716
rect 65100 17108 65156 17118
rect 64988 15876 65044 15886
rect 64988 15782 65044 15820
rect 63868 15652 63924 15662
rect 63868 15538 63924 15596
rect 63868 15486 63870 15538
rect 63922 15486 63924 15538
rect 63868 15474 63924 15486
rect 64652 15428 64708 15438
rect 64652 15334 64708 15372
rect 64764 15314 64820 15326
rect 64764 15262 64766 15314
rect 64818 15262 64820 15314
rect 64764 15148 64820 15262
rect 65100 15148 65156 17052
rect 65548 16884 65604 16894
rect 65548 16100 65604 16828
rect 65324 16044 65604 16100
rect 64092 15092 64148 15102
rect 63308 13918 63310 13970
rect 63362 13918 63364 13970
rect 63308 13906 63364 13918
rect 63532 13972 63588 13982
rect 63532 13878 63588 13916
rect 63644 13970 63700 14476
rect 63980 14530 64036 14542
rect 63980 14478 63982 14530
rect 64034 14478 64036 14530
rect 63980 14420 64036 14478
rect 64092 14530 64148 15036
rect 64428 15092 64820 15148
rect 64876 15092 65156 15148
rect 65212 15426 65268 15438
rect 65212 15374 65214 15426
rect 65266 15374 65268 15426
rect 64428 14642 64484 15092
rect 64428 14590 64430 14642
rect 64482 14590 64484 14642
rect 64428 14578 64484 14590
rect 64540 14644 64596 14654
rect 64092 14478 64094 14530
rect 64146 14478 64148 14530
rect 64092 14466 64148 14478
rect 64540 14530 64596 14588
rect 64540 14478 64542 14530
rect 64594 14478 64596 14530
rect 64540 14466 64596 14478
rect 63980 14354 64036 14364
rect 64316 14306 64372 14318
rect 64316 14254 64318 14306
rect 64370 14254 64372 14306
rect 63644 13918 63646 13970
rect 63698 13918 63700 13970
rect 63644 13906 63700 13918
rect 63868 14084 63924 14094
rect 62860 13766 62916 13804
rect 63868 13858 63924 14028
rect 63868 13806 63870 13858
rect 63922 13806 63924 13858
rect 63868 13794 63924 13806
rect 63420 13748 63476 13758
rect 63420 13654 63476 13692
rect 64316 13748 64372 14254
rect 64876 14308 64932 15092
rect 65212 14644 65268 15374
rect 65324 14756 65380 16044
rect 65324 14690 65380 14700
rect 65436 15876 65492 15886
rect 65660 15876 65716 15886
rect 65436 15874 65716 15876
rect 65436 15822 65438 15874
rect 65490 15822 65662 15874
rect 65714 15822 65716 15874
rect 65436 15820 65716 15822
rect 64428 13748 64484 13758
rect 64316 13746 64484 13748
rect 64316 13694 64430 13746
rect 64482 13694 64484 13746
rect 64316 13692 64484 13694
rect 64204 13636 64260 13646
rect 62860 13076 62916 13086
rect 62860 12290 62916 13020
rect 63756 13076 63812 13086
rect 63756 12982 63812 13020
rect 64204 13074 64260 13580
rect 64204 13022 64206 13074
rect 64258 13022 64260 13074
rect 64204 13010 64260 13022
rect 63980 12740 64036 12750
rect 62860 12238 62862 12290
rect 62914 12238 62916 12290
rect 62860 12226 62916 12238
rect 63868 12628 63924 12638
rect 63420 12178 63476 12190
rect 63420 12126 63422 12178
rect 63474 12126 63476 12178
rect 63308 12068 63364 12078
rect 63420 12068 63476 12126
rect 63868 12180 63924 12572
rect 63868 12086 63924 12124
rect 63364 12012 63476 12068
rect 63308 12002 63364 12012
rect 63868 10500 63924 10510
rect 63868 10052 63924 10444
rect 63756 9996 63924 10052
rect 63084 9156 63140 9166
rect 63140 9100 63364 9156
rect 63084 9062 63140 9100
rect 63196 8372 63252 8382
rect 63084 8316 63196 8372
rect 62972 7586 63028 7598
rect 62972 7534 62974 7586
rect 63026 7534 63028 7586
rect 62972 6692 63028 7534
rect 62972 6626 63028 6636
rect 63084 6916 63140 8316
rect 63196 8306 63252 8316
rect 63308 8370 63364 9100
rect 63308 8318 63310 8370
rect 63362 8318 63364 8370
rect 63308 8306 63364 8318
rect 63532 9154 63588 9166
rect 63532 9102 63534 9154
rect 63586 9102 63588 9154
rect 62972 5908 63028 5918
rect 63084 5908 63140 6860
rect 63532 8148 63588 9102
rect 63756 9156 63812 9996
rect 63756 9042 63812 9100
rect 63756 8990 63758 9042
rect 63810 8990 63812 9042
rect 63756 8978 63812 8990
rect 63980 9938 64036 12684
rect 63980 9886 63982 9938
rect 64034 9886 64036 9938
rect 63980 9044 64036 9886
rect 63980 8978 64036 8988
rect 64316 8372 64372 13692
rect 64428 13682 64484 13692
rect 64540 13412 64596 13422
rect 64540 12402 64596 13356
rect 64876 12850 64932 14252
rect 65100 14588 65268 14644
rect 65100 13076 65156 14588
rect 65436 14420 65492 15820
rect 65660 15810 65716 15820
rect 65772 15652 65828 17612
rect 65884 17556 65940 18060
rect 65996 17780 66052 17790
rect 65996 17686 66052 17724
rect 65884 17500 66052 17556
rect 65884 16882 65940 16894
rect 65884 16830 65886 16882
rect 65938 16830 65940 16882
rect 65884 15764 65940 16830
rect 65884 15698 65940 15708
rect 65660 15596 65828 15652
rect 65324 14364 65492 14420
rect 65548 15426 65604 15438
rect 65548 15374 65550 15426
rect 65602 15374 65604 15426
rect 65324 13636 65380 14364
rect 65436 14196 65492 14206
rect 65436 13860 65492 14140
rect 65548 13972 65604 15374
rect 65660 14644 65716 15596
rect 65660 14578 65716 14588
rect 65996 14642 66052 17500
rect 66108 15092 66164 19966
rect 66332 19684 66388 23772
rect 66444 23826 66500 23838
rect 66444 23774 66446 23826
rect 66498 23774 66500 23826
rect 66444 22594 66500 23774
rect 66444 22542 66446 22594
rect 66498 22542 66500 22594
rect 66444 22530 66500 22542
rect 66556 21476 66612 25788
rect 66780 25396 66836 25406
rect 66892 25396 66948 26460
rect 66836 25340 66948 25396
rect 66780 25330 66836 25340
rect 66780 23714 66836 23726
rect 66780 23662 66782 23714
rect 66834 23662 66836 23714
rect 66780 23266 66836 23662
rect 66780 23214 66782 23266
rect 66834 23214 66836 23266
rect 66780 23202 66836 23214
rect 66892 23492 66948 23502
rect 66780 22596 66836 22606
rect 66892 22596 66948 23436
rect 67004 22820 67060 26852
rect 67452 25618 67508 27020
rect 67564 27010 67620 27020
rect 67452 25566 67454 25618
rect 67506 25566 67508 25618
rect 67452 25554 67508 25566
rect 67116 25506 67172 25518
rect 67116 25454 67118 25506
rect 67170 25454 67172 25506
rect 67116 23828 67172 25454
rect 67340 25508 67396 25518
rect 67340 25414 67396 25452
rect 67788 25394 67844 32508
rect 69244 32452 69300 32462
rect 69244 32358 69300 32396
rect 68832 32172 69096 32182
rect 68888 32116 68936 32172
rect 68992 32116 69040 32172
rect 68832 32106 69096 32116
rect 69692 31948 69748 33068
rect 69356 31892 69748 31948
rect 69804 32450 69860 32462
rect 69804 32398 69806 32450
rect 69858 32398 69860 32450
rect 69804 31948 69860 32398
rect 69804 31892 69972 31948
rect 69132 31666 69188 31678
rect 69132 31614 69134 31666
rect 69186 31614 69188 31666
rect 69132 31556 69188 31614
rect 69132 31490 69188 31500
rect 68124 30882 68180 30894
rect 68124 30830 68126 30882
rect 68178 30830 68180 30882
rect 68124 30212 68180 30830
rect 68832 30604 69096 30614
rect 68888 30548 68936 30604
rect 68992 30548 69040 30604
rect 68832 30538 69096 30548
rect 69132 30436 69188 30446
rect 68572 30324 68628 30334
rect 68572 30212 68628 30268
rect 68124 30210 68628 30212
rect 68124 30158 68574 30210
rect 68626 30158 68628 30210
rect 68124 30156 68628 30158
rect 68348 29986 68404 29998
rect 68348 29934 68350 29986
rect 68402 29934 68404 29986
rect 68348 29876 68404 29934
rect 68348 29810 68404 29820
rect 67900 29316 67956 29326
rect 67900 29222 67956 29260
rect 68460 26908 68516 30156
rect 68572 30146 68628 30156
rect 69132 30210 69188 30380
rect 69132 30158 69134 30210
rect 69186 30158 69188 30210
rect 69132 30146 69188 30158
rect 68832 29036 69096 29046
rect 68888 28980 68936 29036
rect 68992 28980 69040 29036
rect 68832 28970 69096 28980
rect 68572 27860 68628 27870
rect 68572 27766 68628 27804
rect 68684 27858 68740 27870
rect 68684 27806 68686 27858
rect 68738 27806 68740 27858
rect 68236 26852 68516 26908
rect 68684 26964 68740 27806
rect 68908 27860 68964 27870
rect 69132 27860 69188 27870
rect 68908 27858 69076 27860
rect 68908 27806 68910 27858
rect 68962 27806 69076 27858
rect 68908 27804 69076 27806
rect 68908 27794 68964 27804
rect 68796 27748 68852 27758
rect 68796 27654 68852 27692
rect 69020 27748 69076 27804
rect 69132 27858 69300 27860
rect 69132 27806 69134 27858
rect 69186 27806 69300 27858
rect 69132 27804 69300 27806
rect 69132 27794 69188 27804
rect 69020 27682 69076 27692
rect 68832 27468 69096 27478
rect 68888 27412 68936 27468
rect 68992 27412 69040 27468
rect 68832 27402 69096 27412
rect 69244 27300 69300 27804
rect 68684 26898 68740 26908
rect 69132 27244 69300 27300
rect 68124 26290 68180 26302
rect 68124 26238 68126 26290
rect 68178 26238 68180 26290
rect 68124 26068 68180 26238
rect 68124 26002 68180 26012
rect 67788 25342 67790 25394
rect 67842 25342 67844 25394
rect 67116 23762 67172 23772
rect 67564 25282 67620 25294
rect 67564 25230 67566 25282
rect 67618 25230 67620 25282
rect 67452 23268 67508 23278
rect 67340 23044 67396 23054
rect 67004 22764 67172 22820
rect 66780 22594 66948 22596
rect 66780 22542 66782 22594
rect 66834 22542 66948 22594
rect 66780 22540 66948 22542
rect 66780 22530 66836 22540
rect 67004 22484 67060 22494
rect 67004 22258 67060 22428
rect 67004 22206 67006 22258
rect 67058 22206 67060 22258
rect 67004 22194 67060 22206
rect 67116 22036 67172 22764
rect 67004 21980 67172 22036
rect 66892 21812 66948 21822
rect 66892 21718 66948 21756
rect 66668 21476 66724 21486
rect 66556 21420 66668 21476
rect 66668 20018 66724 21420
rect 67004 20804 67060 21980
rect 67116 21700 67172 21710
rect 67116 21606 67172 21644
rect 67228 21586 67284 21598
rect 67228 21534 67230 21586
rect 67282 21534 67284 21586
rect 67228 21476 67284 21534
rect 67228 21410 67284 21420
rect 67004 20738 67060 20748
rect 67228 20914 67284 20926
rect 67228 20862 67230 20914
rect 67282 20862 67284 20914
rect 66668 19966 66670 20018
rect 66722 19966 66724 20018
rect 66668 19954 66724 19966
rect 67116 20132 67172 20142
rect 66332 19628 66500 19684
rect 66444 19236 66500 19628
rect 66332 16996 66388 17006
rect 66220 16772 66276 16782
rect 66220 16210 66276 16716
rect 66220 16158 66222 16210
rect 66274 16158 66276 16210
rect 66220 16146 66276 16158
rect 66332 15314 66388 16940
rect 66444 16882 66500 19180
rect 67004 18900 67060 18910
rect 66780 18564 66836 18574
rect 66836 18508 66948 18564
rect 66780 18498 66836 18508
rect 66668 18450 66724 18462
rect 66668 18398 66670 18450
rect 66722 18398 66724 18450
rect 66556 17444 66612 17454
rect 66556 17350 66612 17388
rect 66668 17108 66724 18398
rect 66668 17042 66724 17052
rect 66444 16830 66446 16882
rect 66498 16830 66500 16882
rect 66444 16818 66500 16830
rect 66556 16884 66612 16894
rect 66780 16884 66836 16894
rect 66612 16882 66836 16884
rect 66612 16830 66782 16882
rect 66834 16830 66836 16882
rect 66612 16828 66836 16830
rect 66556 16818 66612 16828
rect 66780 16818 66836 16828
rect 66892 16660 66948 18508
rect 67004 17778 67060 18844
rect 67116 18338 67172 20076
rect 67228 20020 67284 20862
rect 67228 19954 67284 19964
rect 67116 18286 67118 18338
rect 67170 18286 67172 18338
rect 67116 18274 67172 18286
rect 67004 17726 67006 17778
rect 67058 17726 67060 17778
rect 67004 17714 67060 17726
rect 67340 16772 67396 22988
rect 67452 22258 67508 23212
rect 67452 22206 67454 22258
rect 67506 22206 67508 22258
rect 67452 22194 67508 22206
rect 67564 18900 67620 25230
rect 67788 25060 67844 25342
rect 68236 25284 68292 26852
rect 68572 26290 68628 26302
rect 68572 26238 68574 26290
rect 68626 26238 68628 26290
rect 68572 25732 68628 26238
rect 69132 26292 69188 27244
rect 69356 27188 69412 31892
rect 69804 31666 69860 31678
rect 69804 31614 69806 31666
rect 69858 31614 69860 31666
rect 69468 31556 69524 31566
rect 69804 31556 69860 31614
rect 69468 31554 69860 31556
rect 69468 31502 69470 31554
rect 69522 31502 69860 31554
rect 69468 31500 69860 31502
rect 69468 31490 69524 31500
rect 69804 31332 69860 31500
rect 69916 31556 69972 31892
rect 69916 31490 69972 31500
rect 70028 31556 70084 33294
rect 70700 32676 70756 32686
rect 71372 32676 71428 34190
rect 71596 32786 71652 35646
rect 71596 32734 71598 32786
rect 71650 32734 71652 32786
rect 71596 32722 71652 32734
rect 72380 32788 72436 36316
rect 73164 35698 73220 35710
rect 73164 35646 73166 35698
rect 73218 35646 73220 35698
rect 72492 35588 72548 35598
rect 73164 35588 73220 35646
rect 72492 35586 73220 35588
rect 72492 35534 72494 35586
rect 72546 35534 73220 35586
rect 72492 35532 73220 35534
rect 72492 35522 72548 35532
rect 73164 35308 73220 35532
rect 73164 35252 73556 35308
rect 73052 35026 73108 35038
rect 73052 34974 73054 35026
rect 73106 34974 73108 35026
rect 73052 34356 73108 34974
rect 73500 34468 73556 35252
rect 73724 35026 73780 36876
rect 73724 34974 73726 35026
rect 73778 34974 73780 35026
rect 73724 34962 73780 34974
rect 73500 34412 73892 34468
rect 73052 34300 73668 34356
rect 73052 34132 73108 34300
rect 73052 34066 73108 34076
rect 73164 34130 73220 34142
rect 73164 34078 73166 34130
rect 73218 34078 73220 34130
rect 72940 33460 72996 33470
rect 72940 33366 72996 33404
rect 73164 33236 73220 34078
rect 72380 32786 72772 32788
rect 72380 32734 72382 32786
rect 72434 32734 72772 32786
rect 72380 32732 72772 32734
rect 72380 32722 72436 32732
rect 70700 32674 71428 32676
rect 70700 32622 70702 32674
rect 70754 32622 71428 32674
rect 70700 32620 71428 32622
rect 70700 32610 70756 32620
rect 70476 32562 70532 32574
rect 70476 32510 70478 32562
rect 70530 32510 70532 32562
rect 70476 32452 70532 32510
rect 70476 32386 70532 32396
rect 70476 31778 70532 31790
rect 70476 31726 70478 31778
rect 70530 31726 70532 31778
rect 70140 31556 70196 31566
rect 70476 31556 70532 31726
rect 70028 31554 70532 31556
rect 70028 31502 70142 31554
rect 70194 31502 70532 31554
rect 70028 31500 70532 31502
rect 69804 31276 69972 31332
rect 69804 31106 69860 31118
rect 69804 31054 69806 31106
rect 69858 31054 69860 31106
rect 69804 30322 69860 31054
rect 69916 31108 69972 31276
rect 69916 31042 69972 31052
rect 69916 30436 69972 30446
rect 70028 30436 70084 31500
rect 70140 31490 70196 31500
rect 69972 30380 70084 30436
rect 70140 30994 70196 31006
rect 70140 30942 70142 30994
rect 70194 30942 70196 30994
rect 69916 30370 69972 30380
rect 69804 30270 69806 30322
rect 69858 30270 69860 30322
rect 69804 30258 69860 30270
rect 70140 29650 70196 30942
rect 70140 29598 70142 29650
rect 70194 29598 70196 29650
rect 70140 29586 70196 29598
rect 70700 29538 70756 29550
rect 70700 29486 70702 29538
rect 70754 29486 70756 29538
rect 69692 29316 69748 29326
rect 69692 28644 69748 29260
rect 70700 29316 70756 29486
rect 70924 29540 70980 32620
rect 72716 32562 72772 32732
rect 72716 32510 72718 32562
rect 72770 32510 72772 32562
rect 72716 32498 72772 32510
rect 71260 32340 71316 32350
rect 71260 32246 71316 32284
rect 71260 31668 71316 31678
rect 71036 31666 71316 31668
rect 71036 31614 71262 31666
rect 71314 31614 71316 31666
rect 71036 31612 71316 31614
rect 71036 31218 71092 31612
rect 71260 31602 71316 31612
rect 71036 31166 71038 31218
rect 71090 31166 71092 31218
rect 71036 31154 71092 31166
rect 71372 30994 71428 31006
rect 71372 30942 71374 30994
rect 71426 30942 71428 30994
rect 71372 30212 71428 30942
rect 72492 30882 72548 30894
rect 72492 30830 72494 30882
rect 72546 30830 72548 30882
rect 72492 30324 72548 30830
rect 72492 30268 72884 30324
rect 71372 30146 71428 30156
rect 72828 30210 72884 30268
rect 72828 30158 72830 30210
rect 72882 30158 72884 30210
rect 72716 30098 72772 30110
rect 72716 30046 72718 30098
rect 72770 30046 72772 30098
rect 71484 29988 71540 29998
rect 71036 29540 71092 29550
rect 70924 29484 71036 29540
rect 71036 29446 71092 29484
rect 70700 29250 70756 29260
rect 70476 29202 70532 29214
rect 70476 29150 70478 29202
rect 70530 29150 70532 29202
rect 70476 29092 70532 29150
rect 70476 29026 70532 29036
rect 69692 28578 69748 28588
rect 70140 27970 70196 27982
rect 70140 27918 70142 27970
rect 70194 27918 70196 27970
rect 69356 27094 69412 27132
rect 69468 27860 69524 27870
rect 69132 26226 69188 26236
rect 69244 27074 69300 27086
rect 69244 27022 69246 27074
rect 69298 27022 69300 27074
rect 68832 25900 69096 25910
rect 68888 25844 68936 25900
rect 68992 25844 69040 25900
rect 68832 25834 69096 25844
rect 69244 25732 69300 27022
rect 69356 26964 69412 26974
rect 69356 25844 69412 26908
rect 69468 26180 69524 27804
rect 70028 27636 70084 27646
rect 70028 27542 70084 27580
rect 70028 26964 70084 26974
rect 69692 26962 70084 26964
rect 69692 26910 70030 26962
rect 70082 26910 70084 26962
rect 69692 26908 70084 26910
rect 69468 26114 69524 26124
rect 69580 26292 69636 26302
rect 69356 25788 69524 25844
rect 68572 25666 68628 25676
rect 69132 25676 69300 25732
rect 68348 25508 68404 25518
rect 68348 25414 68404 25452
rect 68236 25218 68292 25228
rect 68572 25284 68628 25294
rect 68572 25190 68628 25228
rect 67788 25004 68740 25060
rect 68684 24834 68740 25004
rect 69132 24946 69188 25676
rect 69356 25620 69412 25630
rect 69244 25564 69356 25620
rect 69244 25506 69300 25564
rect 69356 25554 69412 25564
rect 69244 25454 69246 25506
rect 69298 25454 69300 25506
rect 69244 25442 69300 25454
rect 69356 25396 69412 25406
rect 69356 25302 69412 25340
rect 69132 24894 69134 24946
rect 69186 24894 69188 24946
rect 69132 24882 69188 24894
rect 68684 24782 68686 24834
rect 68738 24782 68740 24834
rect 68684 24770 68740 24782
rect 69020 24836 69076 24846
rect 69020 24722 69076 24780
rect 69020 24670 69022 24722
rect 69074 24670 69076 24722
rect 69020 24658 69076 24670
rect 69468 24722 69524 25788
rect 69580 25396 69636 26236
rect 69692 25618 69748 26908
rect 70028 26898 70084 26908
rect 70028 26628 70084 26638
rect 70028 26514 70084 26572
rect 70028 26462 70030 26514
rect 70082 26462 70084 26514
rect 70028 26450 70084 26462
rect 69916 26180 69972 26190
rect 69692 25566 69694 25618
rect 69746 25566 69748 25618
rect 69692 25554 69748 25566
rect 69804 25844 69860 25854
rect 69580 25330 69636 25340
rect 69804 24948 69860 25788
rect 69468 24670 69470 24722
rect 69522 24670 69524 24722
rect 69468 24658 69524 24670
rect 69580 24946 69860 24948
rect 69580 24894 69806 24946
rect 69858 24894 69860 24946
rect 69580 24892 69860 24894
rect 68832 24332 69096 24342
rect 68888 24276 68936 24332
rect 68992 24276 69040 24332
rect 68832 24266 69096 24276
rect 69580 24052 69636 24892
rect 69804 24882 69860 24892
rect 69468 23996 69636 24052
rect 69244 23714 69300 23726
rect 69244 23662 69246 23714
rect 69298 23662 69300 23714
rect 68908 23492 68964 23502
rect 68348 23156 68404 23166
rect 68348 22594 68404 23100
rect 68908 23042 68964 23436
rect 69244 23156 69300 23662
rect 69244 23090 69300 23100
rect 68908 22990 68910 23042
rect 68962 22990 68964 23042
rect 68908 22978 68964 22990
rect 68348 22542 68350 22594
rect 68402 22542 68404 22594
rect 68348 22530 68404 22542
rect 68460 22932 68516 22942
rect 68460 22258 68516 22876
rect 68832 22764 69096 22774
rect 68888 22708 68936 22764
rect 68992 22708 69040 22764
rect 68832 22698 69096 22708
rect 69356 22484 69412 22494
rect 69020 22482 69412 22484
rect 69020 22430 69358 22482
rect 69410 22430 69412 22482
rect 69020 22428 69412 22430
rect 69020 22370 69076 22428
rect 69356 22418 69412 22428
rect 69468 22484 69524 23996
rect 69916 23940 69972 26124
rect 70140 25284 70196 27918
rect 71372 27972 71428 27982
rect 71372 27878 71428 27916
rect 70364 27860 70420 27870
rect 70364 27766 70420 27804
rect 70700 27858 70756 27870
rect 70924 27860 70980 27870
rect 70700 27806 70702 27858
rect 70754 27806 70756 27858
rect 70140 25218 70196 25228
rect 70252 27748 70308 27758
rect 70028 23940 70084 23950
rect 70252 23940 70308 27692
rect 70364 27074 70420 27086
rect 70364 27022 70366 27074
rect 70418 27022 70420 27074
rect 70364 26628 70420 27022
rect 70364 26562 70420 26572
rect 69804 23938 70084 23940
rect 69804 23886 70030 23938
rect 70082 23886 70084 23938
rect 69804 23884 70084 23886
rect 69468 22418 69524 22428
rect 69580 23828 69636 23838
rect 69020 22318 69022 22370
rect 69074 22318 69076 22370
rect 69020 22306 69076 22318
rect 69356 22260 69412 22270
rect 68460 22206 68462 22258
rect 68514 22206 68516 22258
rect 68460 22194 68516 22206
rect 69244 22204 69356 22260
rect 68684 22146 68740 22158
rect 68684 22094 68686 22146
rect 68738 22094 68740 22146
rect 68684 21812 68740 22094
rect 68684 21746 68740 21756
rect 67564 18834 67620 18844
rect 67676 21700 67732 21710
rect 67564 18452 67620 18462
rect 67340 16706 67396 16716
rect 67452 18450 67620 18452
rect 67452 18398 67566 18450
rect 67618 18398 67620 18450
rect 67452 18396 67620 18398
rect 66668 16604 66948 16660
rect 66556 15986 66612 15998
rect 66556 15934 66558 15986
rect 66610 15934 66612 15986
rect 66556 15876 66612 15934
rect 66556 15810 66612 15820
rect 66332 15262 66334 15314
rect 66386 15262 66388 15314
rect 66332 15250 66388 15262
rect 66108 15026 66164 15036
rect 65996 14590 65998 14642
rect 66050 14590 66052 14642
rect 65996 14578 66052 14590
rect 66220 14756 66276 14766
rect 66108 14530 66164 14542
rect 66108 14478 66110 14530
rect 66162 14478 66164 14530
rect 65884 14418 65940 14430
rect 65884 14366 65886 14418
rect 65938 14366 65940 14418
rect 65548 13906 65604 13916
rect 65772 13972 65828 13982
rect 65436 13766 65492 13804
rect 65324 13580 65492 13636
rect 65436 13188 65492 13580
rect 65436 13132 65716 13188
rect 65324 13076 65380 13086
rect 65100 13074 65380 13076
rect 65100 13022 65326 13074
rect 65378 13022 65380 13074
rect 65100 13020 65380 13022
rect 65324 13010 65380 13020
rect 65548 12964 65604 12974
rect 65548 12870 65604 12908
rect 64876 12798 64878 12850
rect 64930 12798 64932 12850
rect 64876 12786 64932 12798
rect 64652 12740 64708 12750
rect 64652 12646 64708 12684
rect 65548 12740 65604 12750
rect 64540 12350 64542 12402
rect 64594 12350 64596 12402
rect 64540 11956 64596 12350
rect 65100 12516 65156 12526
rect 65100 12402 65156 12460
rect 65100 12350 65102 12402
rect 65154 12350 65156 12402
rect 65100 12338 65156 12350
rect 65548 12178 65604 12684
rect 65660 12516 65716 13132
rect 65660 12402 65716 12460
rect 65660 12350 65662 12402
rect 65714 12350 65716 12402
rect 65660 12338 65716 12350
rect 65548 12126 65550 12178
rect 65602 12126 65604 12178
rect 65548 12114 65604 12126
rect 65772 11956 65828 13916
rect 65884 12402 65940 14366
rect 66108 13970 66164 14478
rect 66108 13918 66110 13970
rect 66162 13918 66164 13970
rect 66108 13906 66164 13918
rect 66220 13858 66276 14700
rect 66220 13806 66222 13858
rect 66274 13806 66276 13858
rect 66220 13636 66276 13806
rect 66220 13570 66276 13580
rect 66556 13748 66612 13758
rect 66444 13188 66500 13198
rect 66220 13132 66444 13188
rect 66220 12962 66276 13132
rect 66444 13122 66500 13132
rect 66220 12910 66222 12962
rect 66274 12910 66276 12962
rect 66220 12898 66276 12910
rect 65884 12350 65886 12402
rect 65938 12350 65940 12402
rect 65884 12338 65940 12350
rect 64540 11890 64596 11900
rect 65548 11900 65828 11956
rect 66556 12290 66612 13692
rect 66668 13636 66724 16604
rect 66780 15426 66836 15438
rect 66780 15374 66782 15426
rect 66834 15374 66836 15426
rect 66780 13972 66836 15374
rect 67228 15314 67284 15326
rect 67228 15262 67230 15314
rect 67282 15262 67284 15314
rect 66892 15202 66948 15214
rect 66892 15150 66894 15202
rect 66946 15150 66948 15202
rect 66892 14530 66948 15150
rect 66892 14478 66894 14530
rect 66946 14478 66948 14530
rect 66892 14466 66948 14478
rect 66780 13906 66836 13916
rect 66892 13746 66948 13758
rect 66892 13694 66894 13746
rect 66946 13694 66948 13746
rect 66668 13580 66836 13636
rect 66668 13412 66724 13422
rect 66668 12962 66724 13356
rect 66668 12910 66670 12962
rect 66722 12910 66724 12962
rect 66668 12898 66724 12910
rect 66556 12238 66558 12290
rect 66610 12238 66612 12290
rect 65212 11732 65268 11742
rect 65212 11508 65268 11676
rect 65212 11442 65268 11452
rect 65436 11732 65492 11742
rect 64988 11396 65044 11406
rect 64988 11394 65156 11396
rect 64988 11342 64990 11394
rect 65042 11342 65156 11394
rect 64988 11340 65156 11342
rect 64988 11330 65044 11340
rect 64988 10724 65044 10734
rect 64988 10630 65044 10668
rect 64988 9716 65044 9726
rect 64988 9622 65044 9660
rect 65100 9044 65156 11340
rect 65436 11172 65492 11676
rect 65436 10722 65492 11116
rect 65436 10670 65438 10722
rect 65490 10670 65492 10722
rect 65436 10658 65492 10670
rect 64316 8306 64372 8316
rect 64876 9042 65156 9044
rect 64876 8990 65102 9042
rect 65154 8990 65156 9042
rect 64876 8988 65156 8990
rect 63196 6020 63252 6030
rect 63532 6020 63588 8092
rect 64092 6692 64148 6702
rect 64092 6598 64148 6636
rect 64876 6690 64932 8988
rect 65100 8978 65156 8988
rect 65436 9938 65492 9950
rect 65436 9886 65438 9938
rect 65490 9886 65492 9938
rect 65436 8372 65492 9886
rect 65548 8932 65604 11900
rect 65660 11284 65716 11294
rect 65660 11282 66500 11284
rect 65660 11230 65662 11282
rect 65714 11230 66500 11282
rect 65660 11228 66500 11230
rect 65660 11218 65716 11228
rect 66444 10834 66500 11228
rect 66444 10782 66446 10834
rect 66498 10782 66500 10834
rect 66444 10770 66500 10782
rect 65996 10612 66052 10622
rect 66556 10612 66612 12238
rect 66780 11732 66836 13580
rect 66892 13076 66948 13694
rect 67116 13524 67172 13534
rect 66892 12850 66948 13020
rect 66892 12798 66894 12850
rect 66946 12798 66948 12850
rect 66892 12786 66948 12798
rect 67004 13468 67116 13524
rect 66892 12180 66948 12190
rect 66892 12086 66948 12124
rect 66780 11666 66836 11676
rect 65996 10518 66052 10556
rect 66332 10556 66612 10612
rect 66780 10612 66836 10622
rect 65660 10500 65716 10510
rect 65660 10406 65716 10444
rect 65884 9716 65940 9726
rect 65884 9622 65940 9660
rect 66220 9604 66276 9614
rect 65996 9602 66276 9604
rect 65996 9550 66222 9602
rect 66274 9550 66276 9602
rect 65996 9548 66276 9550
rect 65996 9268 66052 9548
rect 66220 9538 66276 9548
rect 65772 9212 66052 9268
rect 65772 9154 65828 9212
rect 65772 9102 65774 9154
rect 65826 9102 65828 9154
rect 65772 9090 65828 9102
rect 66332 8932 66388 10556
rect 66780 10518 66836 10556
rect 65548 8876 65940 8932
rect 65660 8372 65716 8382
rect 65436 8316 65660 8372
rect 65660 8258 65716 8316
rect 65660 8206 65662 8258
rect 65714 8206 65716 8258
rect 65548 8148 65604 8158
rect 65548 8054 65604 8092
rect 64876 6638 64878 6690
rect 64930 6638 64932 6690
rect 63196 5926 63252 5964
rect 63308 6018 63588 6020
rect 63308 5966 63534 6018
rect 63586 5966 63588 6018
rect 63308 5964 63588 5966
rect 62524 5852 62916 5908
rect 62524 5346 62580 5852
rect 62524 5294 62526 5346
rect 62578 5294 62580 5346
rect 62524 5282 62580 5294
rect 62860 4788 62916 5852
rect 62972 5906 63140 5908
rect 62972 5854 62974 5906
rect 63026 5854 63140 5906
rect 62972 5852 63140 5854
rect 62972 5842 63028 5852
rect 62972 5124 63028 5134
rect 62972 5030 63028 5068
rect 63308 5012 63364 5964
rect 63532 5954 63588 5964
rect 63868 5124 63924 5134
rect 63868 5030 63924 5068
rect 63308 4918 63364 4956
rect 64764 5012 64820 5022
rect 64876 5012 64932 6638
rect 65324 7588 65380 7598
rect 65324 6692 65380 7532
rect 65660 7476 65716 8206
rect 65660 7410 65716 7420
rect 65324 6598 65380 6636
rect 65660 6580 65716 6590
rect 65716 6524 65828 6580
rect 65660 6486 65716 6524
rect 65660 6018 65716 6030
rect 65660 5966 65662 6018
rect 65714 5966 65716 6018
rect 65436 5908 65492 5918
rect 65436 5814 65492 5852
rect 64988 5236 65044 5246
rect 65660 5236 65716 5966
rect 65044 5180 65156 5236
rect 64988 5170 65044 5180
rect 65100 5122 65156 5180
rect 65660 5170 65716 5180
rect 65100 5070 65102 5122
rect 65154 5070 65156 5122
rect 65100 5058 65156 5070
rect 65772 5124 65828 6524
rect 65884 6132 65940 8876
rect 66220 8372 66276 8382
rect 66332 8372 66388 8876
rect 66556 9714 66612 9726
rect 66556 9662 66558 9714
rect 66610 9662 66612 9714
rect 66556 8482 66612 9662
rect 66556 8430 66558 8482
rect 66610 8430 66612 8482
rect 66556 8418 66612 8430
rect 66220 8370 66388 8372
rect 66220 8318 66222 8370
rect 66274 8318 66388 8370
rect 66220 8316 66388 8318
rect 66220 8306 66276 8316
rect 66220 6692 66276 6702
rect 66220 6598 66276 6636
rect 67004 6132 67060 13468
rect 67116 13458 67172 13468
rect 67228 13188 67284 15262
rect 67284 13132 67396 13188
rect 67228 13122 67284 13132
rect 67340 12628 67396 13132
rect 67452 12964 67508 18396
rect 67564 18386 67620 18396
rect 67676 17668 67732 21644
rect 68832 21196 69096 21206
rect 68888 21140 68936 21196
rect 68992 21140 69040 21196
rect 68832 21130 69096 21140
rect 68460 20356 68516 20366
rect 67900 19012 67956 19022
rect 68348 19012 68404 19022
rect 67676 17602 67732 17612
rect 67788 19010 68404 19012
rect 67788 18958 67902 19010
rect 67954 18958 68350 19010
rect 68402 18958 68404 19010
rect 67788 18956 68404 18958
rect 67564 17556 67620 17566
rect 67564 16994 67620 17500
rect 67564 16942 67566 16994
rect 67618 16942 67620 16994
rect 67564 16930 67620 16942
rect 67676 17444 67732 17454
rect 67564 16324 67620 16334
rect 67676 16324 67732 17388
rect 67564 16322 67732 16324
rect 67564 16270 67566 16322
rect 67618 16270 67732 16322
rect 67564 16268 67732 16270
rect 67564 16258 67620 16268
rect 67564 15652 67620 15662
rect 67564 15538 67620 15596
rect 67564 15486 67566 15538
rect 67618 15486 67620 15538
rect 67564 15474 67620 15486
rect 67788 13412 67844 18956
rect 67900 18946 67956 18956
rect 68348 18946 68404 18956
rect 68124 18452 68180 18462
rect 68124 18358 68180 18396
rect 67900 17442 67956 17454
rect 68348 17444 68404 17454
rect 67900 17390 67902 17442
rect 67954 17390 67956 17442
rect 67900 16996 67956 17390
rect 68236 17442 68404 17444
rect 68236 17390 68350 17442
rect 68402 17390 68404 17442
rect 68236 17388 68404 17390
rect 68236 16996 68292 17388
rect 68348 17378 68404 17388
rect 68460 17220 68516 20300
rect 69020 20356 69076 20366
rect 69020 20242 69076 20300
rect 69020 20190 69022 20242
rect 69074 20190 69076 20242
rect 68684 19908 68740 19918
rect 68460 17154 68516 17164
rect 68572 18338 68628 18350
rect 68572 18286 68574 18338
rect 68626 18286 68628 18338
rect 67956 16940 68292 16996
rect 67900 16930 67956 16940
rect 67900 15876 67956 15886
rect 67900 13746 67956 15820
rect 68236 15538 68292 16940
rect 68348 16884 68404 16894
rect 68572 16884 68628 18286
rect 68684 17332 68740 19852
rect 69020 19796 69076 20190
rect 69020 19730 69076 19740
rect 68832 19628 69096 19638
rect 68888 19572 68936 19628
rect 68992 19572 69040 19628
rect 68832 19562 69096 19572
rect 69244 19458 69300 22204
rect 69356 22166 69412 22204
rect 69468 22148 69524 22158
rect 69468 22054 69524 22092
rect 69580 21924 69636 23772
rect 69468 21868 69636 21924
rect 69692 23380 69748 23390
rect 69692 22370 69748 23324
rect 69692 22318 69694 22370
rect 69746 22318 69748 22370
rect 69468 20244 69524 21868
rect 69692 21812 69748 22318
rect 69580 21756 69748 21812
rect 69580 21476 69636 21756
rect 69580 21410 69636 21420
rect 69692 21588 69748 21598
rect 69356 20242 69524 20244
rect 69356 20190 69470 20242
rect 69522 20190 69524 20242
rect 69356 20188 69524 20190
rect 69356 20132 69412 20188
rect 69468 20178 69524 20188
rect 69356 20066 69412 20076
rect 69692 20130 69748 21532
rect 69692 20078 69694 20130
rect 69746 20078 69748 20130
rect 69692 20066 69748 20078
rect 69580 20020 69636 20030
rect 69580 19926 69636 19964
rect 69804 20018 69860 23884
rect 70028 23874 70084 23884
rect 70140 23884 70252 23940
rect 69916 23714 69972 23726
rect 69916 23662 69918 23714
rect 69970 23662 69972 23714
rect 69916 22932 69972 23662
rect 69916 22866 69972 22876
rect 69916 22258 69972 22270
rect 69916 22206 69918 22258
rect 69970 22206 69972 22258
rect 69916 22148 69972 22206
rect 69916 22082 69972 22092
rect 70028 20916 70084 20926
rect 70028 20822 70084 20860
rect 70140 20188 70196 23884
rect 70252 23874 70308 23884
rect 70476 26180 70532 26190
rect 70476 25172 70532 26124
rect 70700 25508 70756 27806
rect 70700 25442 70756 25452
rect 70812 27858 70980 27860
rect 70812 27806 70926 27858
rect 70978 27806 70980 27858
rect 70812 27804 70980 27806
rect 70812 26404 70868 27804
rect 70924 27794 70980 27804
rect 71148 27858 71204 27870
rect 71148 27806 71150 27858
rect 71202 27806 71204 27858
rect 71148 27748 71204 27806
rect 71260 27860 71316 27870
rect 71260 27766 71316 27804
rect 71148 27682 71204 27692
rect 70476 23548 70532 25116
rect 70812 24164 70868 26348
rect 71036 26404 71092 26414
rect 71036 26310 71092 26348
rect 71484 26290 71540 29932
rect 72044 29986 72100 29998
rect 72044 29934 72046 29986
rect 72098 29934 72100 29986
rect 72044 29092 72100 29934
rect 72268 29540 72324 29550
rect 72268 29446 72324 29484
rect 72716 29540 72772 30046
rect 72716 29474 72772 29484
rect 71932 28644 71988 28654
rect 71596 27860 71652 27870
rect 71596 27766 71652 27804
rect 71932 27524 71988 28588
rect 71484 26238 71486 26290
rect 71538 26238 71540 26290
rect 71484 26226 71540 26238
rect 71596 27468 71988 27524
rect 71596 25732 71652 27468
rect 72044 27412 72100 29036
rect 72492 29426 72548 29438
rect 72492 29374 72494 29426
rect 72546 29374 72548 29426
rect 72492 28644 72548 29374
rect 72716 29316 72772 29326
rect 72716 28754 72772 29260
rect 72828 29204 72884 30158
rect 72828 29138 72884 29148
rect 72716 28702 72718 28754
rect 72770 28702 72772 28754
rect 72716 28644 72772 28702
rect 73052 28644 73108 28654
rect 72716 28642 73108 28644
rect 72716 28590 73054 28642
rect 73106 28590 73108 28642
rect 72716 28588 73108 28590
rect 72492 28578 72548 28588
rect 73052 28578 73108 28588
rect 71484 25676 71652 25732
rect 71708 27356 72100 27412
rect 72380 28082 72436 28094
rect 72380 28030 72382 28082
rect 72434 28030 72436 28082
rect 70364 23492 70532 23548
rect 70700 24108 70868 24164
rect 71148 25620 71204 25630
rect 70364 23378 70420 23492
rect 70364 23326 70366 23378
rect 70418 23326 70420 23378
rect 70364 23044 70420 23326
rect 70364 22978 70420 22988
rect 70588 23156 70644 23166
rect 70476 22484 70532 22494
rect 69804 19966 69806 20018
rect 69858 19966 69860 20018
rect 69804 19796 69860 19966
rect 69244 19406 69246 19458
rect 69298 19406 69300 19458
rect 69244 19394 69300 19406
rect 69580 19740 69860 19796
rect 69916 20132 70196 20188
rect 70364 22370 70420 22382
rect 70364 22318 70366 22370
rect 70418 22318 70420 22370
rect 70364 22148 70420 22318
rect 69580 19348 69636 19740
rect 69468 19292 69636 19348
rect 69692 19348 69748 19358
rect 68908 19234 68964 19246
rect 69468 19236 69524 19292
rect 68908 19182 68910 19234
rect 68962 19182 68964 19234
rect 68908 19124 68964 19182
rect 68908 19058 68964 19068
rect 69244 19180 69524 19236
rect 69244 18452 69300 19180
rect 69580 19122 69636 19134
rect 69580 19070 69582 19122
rect 69634 19070 69636 19122
rect 69244 18386 69300 18396
rect 69356 19010 69412 19022
rect 69356 18958 69358 19010
rect 69410 18958 69412 19010
rect 69356 18450 69412 18958
rect 69580 18674 69636 19070
rect 69692 19122 69748 19292
rect 69916 19236 69972 20132
rect 69692 19070 69694 19122
rect 69746 19070 69748 19122
rect 69692 19058 69748 19070
rect 69804 19180 69972 19236
rect 70028 20018 70084 20030
rect 70028 19966 70030 20018
rect 70082 19966 70084 20018
rect 69804 19124 69860 19180
rect 69580 18622 69582 18674
rect 69634 18622 69636 18674
rect 69580 18610 69636 18622
rect 69692 18676 69748 18686
rect 69804 18676 69860 19068
rect 69916 19012 69972 19022
rect 69916 18918 69972 18956
rect 69692 18674 69860 18676
rect 69692 18622 69694 18674
rect 69746 18622 69860 18674
rect 69692 18620 69860 18622
rect 69692 18610 69748 18620
rect 69356 18398 69358 18450
rect 69410 18398 69412 18450
rect 68832 18060 69096 18070
rect 68888 18004 68936 18060
rect 68992 18004 69040 18060
rect 68832 17994 69096 18004
rect 68796 17892 68852 17902
rect 68796 17778 68852 17836
rect 68796 17726 68798 17778
rect 68850 17726 68852 17778
rect 68796 17714 68852 17726
rect 69356 17780 69412 18398
rect 69468 18450 69524 18462
rect 69468 18398 69470 18450
rect 69522 18398 69524 18450
rect 69468 17780 69524 18398
rect 69916 18452 69972 18462
rect 69916 18358 69972 18396
rect 70028 18340 70084 19966
rect 70364 19908 70420 22092
rect 70028 18274 70084 18284
rect 70140 19852 70420 19908
rect 70476 21698 70532 22428
rect 70476 21646 70478 21698
rect 70530 21646 70532 21698
rect 70476 19908 70532 21646
rect 70588 21364 70644 23100
rect 70700 22260 70756 24108
rect 70700 22194 70756 22204
rect 70812 23938 70868 23950
rect 70812 23886 70814 23938
rect 70866 23886 70868 23938
rect 70812 23044 70868 23886
rect 71036 23940 71092 23950
rect 71036 23846 71092 23884
rect 71148 23156 71204 25564
rect 70700 21924 70756 21934
rect 70700 21364 70756 21868
rect 70812 21586 70868 22988
rect 70812 21534 70814 21586
rect 70866 21534 70868 21586
rect 70812 21522 70868 21534
rect 70924 23154 71204 23156
rect 70924 23102 71150 23154
rect 71202 23102 71204 23154
rect 70924 23100 71204 23102
rect 70700 21308 70868 21364
rect 70588 21298 70644 21308
rect 70700 21140 70756 21150
rect 70588 20916 70644 20926
rect 70588 20130 70644 20860
rect 70588 20078 70590 20130
rect 70642 20078 70644 20130
rect 70588 20066 70644 20078
rect 70700 19908 70756 21084
rect 70812 20916 70868 21308
rect 70812 20850 70868 20860
rect 69580 17780 69636 17790
rect 69468 17778 69636 17780
rect 69468 17726 69582 17778
rect 69634 17726 69636 17778
rect 69468 17724 69636 17726
rect 69356 17714 69412 17724
rect 68908 17332 68964 17342
rect 68684 17276 68908 17332
rect 68908 16994 68964 17276
rect 68908 16942 68910 16994
rect 68962 16942 68964 16994
rect 68908 16930 68964 16942
rect 69468 17220 69524 17230
rect 68348 16882 68628 16884
rect 68348 16830 68350 16882
rect 68402 16830 68628 16882
rect 68348 16828 68628 16830
rect 69244 16882 69300 16894
rect 69244 16830 69246 16882
rect 69298 16830 69300 16882
rect 68348 15652 68404 16828
rect 68832 16492 69096 16502
rect 68888 16436 68936 16492
rect 68992 16436 69040 16492
rect 68832 16426 69096 16436
rect 69132 16324 69188 16334
rect 69132 16230 69188 16268
rect 68460 16100 68516 16110
rect 68460 16098 68740 16100
rect 68460 16046 68462 16098
rect 68514 16046 68740 16098
rect 68460 16044 68740 16046
rect 68460 16034 68516 16044
rect 68348 15586 68404 15596
rect 68236 15486 68238 15538
rect 68290 15486 68292 15538
rect 68236 15474 68292 15486
rect 68684 15538 68740 16044
rect 68684 15486 68686 15538
rect 68738 15486 68740 15538
rect 67900 13694 67902 13746
rect 67954 13694 67956 13746
rect 67900 13682 67956 13694
rect 68236 14420 68292 14430
rect 68236 13746 68292 14364
rect 68684 13860 68740 15486
rect 69132 15540 69188 15550
rect 69244 15540 69300 16830
rect 69132 15538 69300 15540
rect 69132 15486 69134 15538
rect 69186 15486 69300 15538
rect 69132 15484 69300 15486
rect 69132 15474 69188 15484
rect 68832 14924 69096 14934
rect 68888 14868 68936 14924
rect 68992 14868 69040 14924
rect 68832 14858 69096 14868
rect 68908 14642 68964 14654
rect 68908 14590 68910 14642
rect 68962 14590 68964 14642
rect 68908 14420 68964 14590
rect 68908 14354 68964 14364
rect 68684 13794 68740 13804
rect 68236 13694 68238 13746
rect 68290 13694 68292 13746
rect 68236 13682 68292 13694
rect 68460 13748 68516 13758
rect 67900 13412 67956 13422
rect 67788 13356 67900 13412
rect 67900 13346 67956 13356
rect 67452 12898 67508 12908
rect 67340 12572 67844 12628
rect 67228 11732 67284 11742
rect 67228 10834 67284 11676
rect 67228 10782 67230 10834
rect 67282 10782 67284 10834
rect 67228 10770 67284 10782
rect 67788 11506 67844 12572
rect 67788 11454 67790 11506
rect 67842 11454 67844 11506
rect 67788 10724 67844 11454
rect 67788 10658 67844 10668
rect 68124 11508 68180 11518
rect 68124 10834 68180 11452
rect 68124 10782 68126 10834
rect 68178 10782 68180 10834
rect 68124 10724 68180 10782
rect 68124 10658 68180 10668
rect 67900 8932 67956 8942
rect 67900 8838 67956 8876
rect 68460 8596 68516 13692
rect 68832 13356 69096 13366
rect 68888 13300 68936 13356
rect 68992 13300 69040 13356
rect 68832 13290 69096 13300
rect 69244 12180 69300 15484
rect 69244 12114 69300 12124
rect 68832 11788 69096 11798
rect 68888 11732 68936 11788
rect 68992 11732 69040 11788
rect 68832 11722 69096 11732
rect 69356 10724 69412 10734
rect 69356 10630 69412 10668
rect 69132 10610 69188 10622
rect 69132 10558 69134 10610
rect 69186 10558 69188 10610
rect 68572 10500 68628 10510
rect 68572 10406 68628 10444
rect 69132 10500 69188 10558
rect 69132 10434 69188 10444
rect 69244 10498 69300 10510
rect 69244 10446 69246 10498
rect 69298 10446 69300 10498
rect 68832 10220 69096 10230
rect 68888 10164 68936 10220
rect 68992 10164 69040 10220
rect 68832 10154 69096 10164
rect 68908 10052 68964 10062
rect 68796 9996 68908 10052
rect 68572 9828 68628 9838
rect 68572 9734 68628 9772
rect 68572 9268 68628 9278
rect 68796 9268 68852 9996
rect 68908 9986 68964 9996
rect 69244 9938 69300 10446
rect 69468 10052 69524 17164
rect 69580 16884 69636 17724
rect 69804 17668 69860 17678
rect 69580 16818 69636 16828
rect 69692 17612 69804 17668
rect 69580 16212 69636 16222
rect 69692 16212 69748 17612
rect 69804 17574 69860 17612
rect 69804 16996 69860 17006
rect 69804 16902 69860 16940
rect 69580 16210 69748 16212
rect 69580 16158 69582 16210
rect 69634 16158 69748 16210
rect 69580 16156 69748 16158
rect 69580 13524 69636 16156
rect 70028 15426 70084 15438
rect 70028 15374 70030 15426
rect 70082 15374 70084 15426
rect 69804 15314 69860 15326
rect 69804 15262 69806 15314
rect 69858 15262 69860 15314
rect 69804 15148 69860 15262
rect 69804 15092 69972 15148
rect 69580 13458 69636 13468
rect 69692 14532 69748 14542
rect 69692 12964 69748 14476
rect 69916 13972 69972 15092
rect 70028 14644 70084 15374
rect 70028 14578 70084 14588
rect 70140 14420 70196 19852
rect 70476 19842 70532 19852
rect 70588 19852 70756 19908
rect 70812 20018 70868 20030
rect 70812 19966 70814 20018
rect 70866 19966 70868 20018
rect 70252 19348 70308 19386
rect 70252 19282 70308 19292
rect 70364 19236 70420 19246
rect 70364 19234 70532 19236
rect 70364 19182 70366 19234
rect 70418 19182 70532 19234
rect 70364 19180 70532 19182
rect 70364 19170 70420 19180
rect 70252 19012 70308 19022
rect 70476 19012 70532 19180
rect 70252 18918 70308 18956
rect 70364 18956 70532 19012
rect 70588 19234 70644 19852
rect 70812 19796 70868 19966
rect 70812 19730 70868 19740
rect 70924 19348 70980 23100
rect 71148 23090 71204 23100
rect 71260 24836 71316 24846
rect 71036 22820 71092 22830
rect 71036 21924 71092 22764
rect 71036 21858 71092 21868
rect 71260 21588 71316 24780
rect 71372 23266 71428 23278
rect 71372 23214 71374 23266
rect 71426 23214 71428 23266
rect 71372 21700 71428 23214
rect 71484 23268 71540 25676
rect 71596 25508 71652 25518
rect 71708 25508 71764 27356
rect 72156 27076 72212 27086
rect 72156 26982 72212 27020
rect 71596 25506 71764 25508
rect 71596 25454 71598 25506
rect 71650 25454 71764 25506
rect 71596 25452 71764 25454
rect 71932 26068 71988 26078
rect 71932 25506 71988 26012
rect 72380 25956 72436 28030
rect 72604 28082 72660 28094
rect 73164 28084 73220 33180
rect 72604 28030 72606 28082
rect 72658 28030 72660 28082
rect 72604 27076 72660 28030
rect 72940 28028 73220 28084
rect 73276 33460 73332 33470
rect 73276 32340 73332 33404
rect 72828 27860 72884 27870
rect 72828 27766 72884 27804
rect 72604 27010 72660 27020
rect 72492 26402 72548 26414
rect 72492 26350 72494 26402
rect 72546 26350 72548 26402
rect 72492 26180 72548 26350
rect 72492 26114 72548 26124
rect 72828 26290 72884 26302
rect 72828 26238 72830 26290
rect 72882 26238 72884 26290
rect 72380 25890 72436 25900
rect 72156 25732 72212 25742
rect 72156 25620 72212 25676
rect 72156 25564 72324 25620
rect 71932 25454 71934 25506
rect 71986 25454 71988 25506
rect 71596 24724 71652 25452
rect 71596 24658 71652 24668
rect 71708 24610 71764 24622
rect 71708 24558 71710 24610
rect 71762 24558 71764 24610
rect 71708 24164 71764 24558
rect 71708 24098 71764 24108
rect 71820 24276 71876 24286
rect 71484 23202 71540 23212
rect 71596 23826 71652 23838
rect 71596 23774 71598 23826
rect 71650 23774 71652 23826
rect 71372 21634 71428 21644
rect 71484 23042 71540 23054
rect 71484 22990 71486 23042
rect 71538 22990 71540 23042
rect 70588 19182 70590 19234
rect 70642 19182 70644 19234
rect 70364 16996 70420 18956
rect 70588 18900 70644 19182
rect 70588 18834 70644 18844
rect 70700 19292 70980 19348
rect 71036 21586 71316 21588
rect 71036 21534 71262 21586
rect 71314 21534 71316 21586
rect 71036 21532 71316 21534
rect 70588 18674 70644 18686
rect 70588 18622 70590 18674
rect 70642 18622 70644 18674
rect 70476 18562 70532 18574
rect 70476 18510 70478 18562
rect 70530 18510 70532 18562
rect 70476 17332 70532 18510
rect 70588 18564 70644 18622
rect 70588 18498 70644 18508
rect 70476 17266 70532 17276
rect 70476 16996 70532 17006
rect 70364 16994 70532 16996
rect 70364 16942 70478 16994
rect 70530 16942 70532 16994
rect 70364 16940 70532 16942
rect 70364 14420 70420 14430
rect 70140 14364 70364 14420
rect 70028 13972 70084 13982
rect 69916 13970 70084 13972
rect 69916 13918 70030 13970
rect 70082 13918 70084 13970
rect 69916 13916 70084 13918
rect 70028 13906 70084 13916
rect 70364 13746 70420 14364
rect 70364 13694 70366 13746
rect 70418 13694 70420 13746
rect 70364 13682 70420 13694
rect 70476 13524 70532 16940
rect 70700 16996 70756 19292
rect 70812 19122 70868 19134
rect 70812 19070 70814 19122
rect 70866 19070 70868 19122
rect 70812 18676 70868 19070
rect 70812 18610 70868 18620
rect 70812 18450 70868 18462
rect 70812 18398 70814 18450
rect 70866 18398 70868 18450
rect 70812 18340 70868 18398
rect 70812 18274 70868 18284
rect 71036 18340 71092 21532
rect 71260 21522 71316 21532
rect 71372 21474 71428 21486
rect 71372 21422 71374 21474
rect 71426 21422 71428 21474
rect 71148 21364 71204 21374
rect 71148 20020 71204 21308
rect 71372 20802 71428 21422
rect 71372 20750 71374 20802
rect 71426 20750 71428 20802
rect 71372 20738 71428 20750
rect 71484 20692 71540 22990
rect 71596 22932 71652 23774
rect 71820 23604 71876 24220
rect 71820 23538 71876 23548
rect 71596 22866 71652 22876
rect 71484 20626 71540 20636
rect 71596 22314 71652 22326
rect 71596 22262 71598 22314
rect 71650 22262 71652 22314
rect 71596 22260 71652 22262
rect 71596 20244 71652 22204
rect 71932 22260 71988 25454
rect 72268 25506 72324 25564
rect 72268 25454 72270 25506
rect 72322 25454 72324 25506
rect 72156 25284 72212 25294
rect 72156 24946 72212 25228
rect 72268 25172 72324 25454
rect 72268 25106 72324 25116
rect 72380 25508 72436 25518
rect 72156 24894 72158 24946
rect 72210 24894 72212 24946
rect 72156 24882 72212 24894
rect 72268 24834 72324 24846
rect 72268 24782 72270 24834
rect 72322 24782 72324 24834
rect 72268 24276 72324 24782
rect 72268 24210 72324 24220
rect 72268 24052 72324 24062
rect 72380 24052 72436 25452
rect 72716 25508 72772 25518
rect 72604 24724 72660 24734
rect 72604 24630 72660 24668
rect 72268 24050 72436 24052
rect 72268 23998 72270 24050
rect 72322 23998 72436 24050
rect 72268 23996 72436 23998
rect 72268 23986 72324 23996
rect 72156 23940 72212 23950
rect 72044 23938 72212 23940
rect 72044 23886 72158 23938
rect 72210 23886 72212 23938
rect 72044 23884 72212 23886
rect 72044 23828 72100 23884
rect 72156 23874 72212 23884
rect 72604 23940 72660 23950
rect 72044 23762 72100 23772
rect 72268 23828 72324 23838
rect 72156 23604 72212 23614
rect 72156 23380 72212 23548
rect 72268 23492 72324 23772
rect 72492 23716 72548 23726
rect 72604 23716 72660 23884
rect 72716 23938 72772 25452
rect 72716 23886 72718 23938
rect 72770 23886 72772 23938
rect 72716 23874 72772 23886
rect 72828 23828 72884 26238
rect 72828 23762 72884 23772
rect 72492 23714 72660 23716
rect 72492 23662 72494 23714
rect 72546 23662 72660 23714
rect 72492 23660 72660 23662
rect 72492 23650 72548 23660
rect 72268 23426 72324 23436
rect 72380 23604 72436 23614
rect 72156 23314 72212 23324
rect 72268 22932 72324 22942
rect 72268 22708 72324 22876
rect 72268 22370 72324 22652
rect 72268 22318 72270 22370
rect 72322 22318 72324 22370
rect 72268 22306 72324 22318
rect 71932 22194 71988 22204
rect 72380 22148 72436 23548
rect 72940 23548 72996 28028
rect 73276 27972 73332 32284
rect 73388 31890 73444 31902
rect 73388 31838 73390 31890
rect 73442 31838 73444 31890
rect 73388 30324 73444 31838
rect 73388 30322 73556 30324
rect 73388 30270 73390 30322
rect 73442 30270 73556 30322
rect 73388 30268 73556 30270
rect 73388 30258 73444 30268
rect 73276 27970 73444 27972
rect 73276 27918 73278 27970
rect 73330 27918 73444 27970
rect 73276 27916 73444 27918
rect 73276 27906 73332 27916
rect 73164 27858 73220 27870
rect 73164 27806 73166 27858
rect 73218 27806 73220 27858
rect 73164 27188 73220 27806
rect 73052 27132 73220 27188
rect 73052 24836 73108 27132
rect 73164 26962 73220 26974
rect 73164 26910 73166 26962
rect 73218 26910 73220 26962
rect 73164 26514 73220 26910
rect 73164 26462 73166 26514
rect 73218 26462 73220 26514
rect 73164 26450 73220 26462
rect 73164 26290 73220 26302
rect 73164 26238 73166 26290
rect 73218 26238 73220 26290
rect 73164 25620 73220 26238
rect 73164 25554 73220 25564
rect 73052 24770 73108 24780
rect 73276 25284 73332 25294
rect 73052 24164 73108 24174
rect 73052 23938 73108 24108
rect 73052 23886 73054 23938
rect 73106 23886 73108 23938
rect 73052 23874 73108 23886
rect 72940 23492 73108 23548
rect 72716 23268 72772 23278
rect 72268 22092 72436 22148
rect 72492 23156 72548 23166
rect 72492 23042 72548 23100
rect 72492 22990 72494 23042
rect 72546 22990 72548 23042
rect 71708 21698 71764 21710
rect 71708 21646 71710 21698
rect 71762 21646 71764 21698
rect 71708 21588 71764 21646
rect 72268 21588 72324 22092
rect 72492 21812 72548 22990
rect 71708 21522 71764 21532
rect 71932 21586 72324 21588
rect 71932 21534 72270 21586
rect 72322 21534 72324 21586
rect 71932 21532 72324 21534
rect 71932 21140 71988 21532
rect 72268 21522 72324 21532
rect 72380 21756 72548 21812
rect 72604 21812 72660 21822
rect 72380 21364 72436 21756
rect 72604 21718 72660 21756
rect 72716 21810 72772 23212
rect 72828 23156 72884 23194
rect 72828 23090 72884 23100
rect 73052 22372 73108 23492
rect 73164 23266 73220 23278
rect 73164 23214 73166 23266
rect 73218 23214 73220 23266
rect 73164 22596 73220 23214
rect 73276 23044 73332 25228
rect 73388 24722 73444 27916
rect 73500 27748 73556 30268
rect 73500 27682 73556 27692
rect 73612 26402 73668 34300
rect 73724 30212 73780 30222
rect 73724 30118 73780 30156
rect 73836 29540 73892 34412
rect 73948 34018 74004 38332
rect 74060 36932 74116 36942
rect 74060 36482 74116 36876
rect 75068 36708 75124 36718
rect 75068 36614 75124 36652
rect 74060 36430 74062 36482
rect 74114 36430 74116 36482
rect 74060 36418 74116 36430
rect 75516 35924 75572 39200
rect 75516 35858 75572 35868
rect 76636 35924 76692 35934
rect 76636 35830 76692 35868
rect 75068 35812 75124 35822
rect 75068 35586 75124 35756
rect 75068 35534 75070 35586
rect 75122 35534 75124 35586
rect 75068 35522 75124 35534
rect 76076 35698 76132 35710
rect 76076 35646 76078 35698
rect 76130 35646 76132 35698
rect 76076 35308 76132 35646
rect 76076 35252 76356 35308
rect 75404 34690 75460 34702
rect 75404 34638 75406 34690
rect 75458 34638 75460 34690
rect 73948 33966 73950 34018
rect 74002 33966 74004 34018
rect 73948 33954 74004 33966
rect 75068 34132 75124 34142
rect 75404 34132 75460 34638
rect 76300 34690 76356 35252
rect 76300 34638 76302 34690
rect 76354 34638 76356 34690
rect 76300 34580 76356 34638
rect 76300 34514 76356 34524
rect 75628 34132 75684 34142
rect 75068 32450 75124 34076
rect 75068 32398 75070 32450
rect 75122 32398 75124 32450
rect 75068 32386 75124 32398
rect 75180 34130 75684 34132
rect 75180 34078 75630 34130
rect 75682 34078 75684 34130
rect 75180 34076 75684 34078
rect 73724 29484 73892 29540
rect 73948 31220 74004 31230
rect 73724 28420 73780 29484
rect 73836 29316 73892 29326
rect 73836 28644 73892 29260
rect 73948 29092 74004 31164
rect 74172 31108 74228 31118
rect 74172 31014 74228 31052
rect 74508 31106 74564 31118
rect 74508 31054 74510 31106
rect 74562 31054 74564 31106
rect 74508 30996 74564 31054
rect 74844 30996 74900 31006
rect 74508 30994 74900 30996
rect 74508 30942 74846 30994
rect 74898 30942 74900 30994
rect 74508 30940 74900 30942
rect 74732 30322 74788 30334
rect 74732 30270 74734 30322
rect 74786 30270 74788 30322
rect 74508 30212 74564 30222
rect 74396 29988 74452 29998
rect 74284 29986 74452 29988
rect 74284 29934 74398 29986
rect 74450 29934 74452 29986
rect 74284 29932 74452 29934
rect 74284 29426 74340 29932
rect 74396 29922 74452 29932
rect 74508 29650 74564 30156
rect 74508 29598 74510 29650
rect 74562 29598 74564 29650
rect 74508 29586 74564 29598
rect 74284 29374 74286 29426
rect 74338 29374 74340 29426
rect 74284 29362 74340 29374
rect 74732 29316 74788 30270
rect 74844 29426 74900 30940
rect 74844 29374 74846 29426
rect 74898 29374 74900 29426
rect 74844 29362 74900 29374
rect 74732 29250 74788 29260
rect 73948 29026 74004 29036
rect 73892 28588 74228 28644
rect 73836 28578 73892 28588
rect 73724 28364 73892 28420
rect 73724 28196 73780 28206
rect 73724 27298 73780 28140
rect 73724 27246 73726 27298
rect 73778 27246 73780 27298
rect 73724 27234 73780 27246
rect 73612 26350 73614 26402
rect 73666 26350 73668 26402
rect 73500 25508 73556 25518
rect 73500 25414 73556 25452
rect 73612 24948 73668 26350
rect 73724 27074 73780 27086
rect 73724 27022 73726 27074
rect 73778 27022 73780 27074
rect 73724 25618 73780 27022
rect 73724 25566 73726 25618
rect 73778 25566 73780 25618
rect 73724 25554 73780 25566
rect 73724 24948 73780 24958
rect 73612 24892 73724 24948
rect 73724 24882 73780 24892
rect 73836 24836 73892 28364
rect 74172 28082 74228 28588
rect 75180 28196 75236 34076
rect 75628 34066 75684 34076
rect 77980 34132 78036 39200
rect 78492 36092 78756 36102
rect 78548 36036 78596 36092
rect 78652 36036 78700 36092
rect 78492 36026 78756 36036
rect 78492 34524 78756 34534
rect 78548 34468 78596 34524
rect 78652 34468 78700 34524
rect 78492 34458 78756 34468
rect 77980 34066 78036 34076
rect 77980 33906 78036 33918
rect 77980 33854 77982 33906
rect 78034 33854 78036 33906
rect 77980 33460 78036 33854
rect 77980 33394 78036 33404
rect 76300 33236 76356 33246
rect 76300 33142 76356 33180
rect 75404 33124 75460 33134
rect 75460 33068 75684 33124
rect 75404 33030 75460 33068
rect 75628 32562 75684 33068
rect 78492 32956 78756 32966
rect 78548 32900 78596 32956
rect 78652 32900 78700 32956
rect 78492 32890 78756 32900
rect 75628 32510 75630 32562
rect 75682 32510 75684 32562
rect 75628 32498 75684 32510
rect 77980 32338 78036 32350
rect 77980 32286 77982 32338
rect 78034 32286 78036 32338
rect 75404 31778 75460 31790
rect 75404 31726 75406 31778
rect 75458 31726 75460 31778
rect 75180 28130 75236 28140
rect 75292 30884 75348 30894
rect 75292 30098 75348 30828
rect 75292 30046 75294 30098
rect 75346 30046 75348 30098
rect 74172 28030 74174 28082
rect 74226 28030 74228 28082
rect 74172 27076 74228 28030
rect 75068 27970 75124 27982
rect 75068 27918 75070 27970
rect 75122 27918 75124 27970
rect 74732 27860 74788 27870
rect 74396 27858 74788 27860
rect 74396 27806 74734 27858
rect 74786 27806 74788 27858
rect 74396 27804 74788 27806
rect 74396 27298 74452 27804
rect 74732 27794 74788 27804
rect 74396 27246 74398 27298
rect 74450 27246 74452 27298
rect 74396 27234 74452 27246
rect 74732 27076 74788 27086
rect 74172 27074 74788 27076
rect 74172 27022 74734 27074
rect 74786 27022 74788 27074
rect 74172 27020 74788 27022
rect 74732 27010 74788 27020
rect 73948 26404 74004 26414
rect 73948 25396 74004 26348
rect 74956 26404 75012 26414
rect 75068 26404 75124 27918
rect 75292 27860 75348 30046
rect 75404 30100 75460 31726
rect 75628 31556 75684 31566
rect 75628 31554 75796 31556
rect 75628 31502 75630 31554
rect 75682 31502 75796 31554
rect 75628 31500 75796 31502
rect 75628 31490 75684 31500
rect 75628 30882 75684 30894
rect 75628 30830 75630 30882
rect 75682 30830 75684 30882
rect 75404 30034 75460 30044
rect 75516 30210 75572 30222
rect 75516 30158 75518 30210
rect 75570 30158 75572 30210
rect 75516 29988 75572 30158
rect 75628 30212 75684 30830
rect 75628 30146 75684 30156
rect 75516 29922 75572 29932
rect 75628 29540 75684 29550
rect 75740 29540 75796 31500
rect 77980 30996 78036 32286
rect 78492 31388 78756 31398
rect 78548 31332 78596 31388
rect 78652 31332 78700 31388
rect 78492 31322 78756 31332
rect 77980 30930 78036 30940
rect 77756 30884 77812 30894
rect 77756 30790 77812 30828
rect 76636 30324 76692 30334
rect 76636 30230 76692 30268
rect 77308 30324 77364 30334
rect 76300 30100 76356 30110
rect 76300 30006 76356 30044
rect 76972 30098 77028 30110
rect 76972 30046 76974 30098
rect 77026 30046 77028 30098
rect 75628 29538 75796 29540
rect 75628 29486 75630 29538
rect 75682 29486 75796 29538
rect 75628 29484 75796 29486
rect 76972 29988 77028 30046
rect 75628 29474 75684 29484
rect 76524 29092 76580 29102
rect 75404 28754 75460 28766
rect 75404 28702 75406 28754
rect 75458 28702 75460 28754
rect 75404 28532 75460 28702
rect 75404 28466 75460 28476
rect 76300 28418 76356 28430
rect 76300 28366 76302 28418
rect 76354 28366 76356 28418
rect 75292 27794 75348 27804
rect 75628 27860 75684 27870
rect 76300 27860 76356 28366
rect 75628 27858 76356 27860
rect 75628 27806 75630 27858
rect 75682 27806 76356 27858
rect 75628 27804 76356 27806
rect 74956 26402 75124 26404
rect 74956 26350 74958 26402
rect 75010 26350 75124 26402
rect 74956 26348 75124 26350
rect 75180 27748 75236 27758
rect 74956 26338 75012 26348
rect 74284 26292 74340 26302
rect 74284 26290 74900 26292
rect 74284 26238 74286 26290
rect 74338 26238 74900 26290
rect 74284 26236 74900 26238
rect 74284 26226 74340 26236
rect 73948 25394 74228 25396
rect 73948 25342 73950 25394
rect 74002 25342 74228 25394
rect 73948 25340 74228 25342
rect 73948 25330 74004 25340
rect 73388 24670 73390 24722
rect 73442 24670 73444 24722
rect 73388 24658 73444 24670
rect 73724 24722 73780 24734
rect 73724 24670 73726 24722
rect 73778 24670 73780 24722
rect 73612 23492 73668 23502
rect 73612 23154 73668 23436
rect 73724 23268 73780 24670
rect 73836 23548 73892 24780
rect 73836 23492 74004 23548
rect 73724 23202 73780 23212
rect 73612 23102 73614 23154
rect 73666 23102 73668 23154
rect 73612 23090 73668 23102
rect 73276 22988 73444 23044
rect 73164 22530 73220 22540
rect 72716 21758 72718 21810
rect 72770 21758 72772 21810
rect 72492 21586 72548 21598
rect 72492 21534 72494 21586
rect 72546 21534 72548 21586
rect 72492 21476 72548 21534
rect 72492 21410 72548 21420
rect 71484 20188 71652 20244
rect 71820 21084 71988 21140
rect 72156 21308 72436 21364
rect 71260 20020 71316 20030
rect 71148 20018 71316 20020
rect 71148 19966 71262 20018
rect 71314 19966 71316 20018
rect 71148 19964 71316 19966
rect 71148 19346 71204 19964
rect 71260 19954 71316 19964
rect 71148 19294 71150 19346
rect 71202 19294 71204 19346
rect 71148 19282 71204 19294
rect 71372 18676 71428 18686
rect 71372 18562 71428 18620
rect 71372 18510 71374 18562
rect 71426 18510 71428 18562
rect 71372 18498 71428 18510
rect 71148 18450 71204 18462
rect 71148 18398 71150 18450
rect 71202 18398 71204 18450
rect 71148 18340 71204 18398
rect 71484 18340 71540 20188
rect 71596 20020 71652 20030
rect 71652 19964 71764 20020
rect 71596 19954 71652 19964
rect 71036 18284 71204 18340
rect 71372 18284 71540 18340
rect 71596 19794 71652 19806
rect 71596 19742 71598 19794
rect 71650 19742 71652 19794
rect 71036 17892 71092 18284
rect 71036 17826 71092 17836
rect 71148 17666 71204 17678
rect 71148 17614 71150 17666
rect 71202 17614 71204 17666
rect 71148 17444 71204 17614
rect 71148 17378 71204 17388
rect 71372 17444 71428 18284
rect 71484 17666 71540 17678
rect 71484 17614 71486 17666
rect 71538 17614 71540 17666
rect 71484 17556 71540 17614
rect 71484 17490 71540 17500
rect 71372 17378 71428 17388
rect 71372 17108 71428 17118
rect 71372 17014 71428 17052
rect 70700 16882 70756 16940
rect 70700 16830 70702 16882
rect 70754 16830 70756 16882
rect 70700 16818 70756 16830
rect 71484 16994 71540 17006
rect 71484 16942 71486 16994
rect 71538 16942 71540 16994
rect 71484 16772 71540 16942
rect 71596 16996 71652 19742
rect 71596 16930 71652 16940
rect 71484 16706 71540 16716
rect 71708 16882 71764 19964
rect 71820 19236 71876 21084
rect 71820 19170 71876 19180
rect 71932 20916 71988 20926
rect 71708 16830 71710 16882
rect 71762 16830 71764 16882
rect 71260 16548 71316 16558
rect 71036 14644 71092 14654
rect 71036 14550 71092 14588
rect 70588 13858 70644 13870
rect 70588 13806 70590 13858
rect 70642 13806 70644 13858
rect 70588 13748 70644 13806
rect 71148 13860 71204 13870
rect 71148 13766 71204 13804
rect 70588 13682 70644 13692
rect 70252 13468 70532 13524
rect 69692 12962 69860 12964
rect 69692 12910 69694 12962
rect 69746 12910 69860 12962
rect 69692 12908 69860 12910
rect 69692 12898 69748 12908
rect 69804 12402 69860 12908
rect 69804 12350 69806 12402
rect 69858 12350 69860 12402
rect 69804 12338 69860 12350
rect 70140 12178 70196 12190
rect 70140 12126 70142 12178
rect 70194 12126 70196 12178
rect 69468 9986 69524 9996
rect 69580 10722 69636 10734
rect 69580 10670 69582 10722
rect 69634 10670 69636 10722
rect 69244 9886 69246 9938
rect 69298 9886 69300 9938
rect 69244 9874 69300 9886
rect 68572 9266 68852 9268
rect 68572 9214 68574 9266
rect 68626 9214 68798 9266
rect 68850 9214 68852 9266
rect 68572 9212 68852 9214
rect 68572 9202 68628 9212
rect 68796 9202 68852 9212
rect 69580 9266 69636 10670
rect 70140 10724 70196 12126
rect 70252 11284 70308 13468
rect 70364 12850 70420 12862
rect 70364 12798 70366 12850
rect 70418 12798 70420 12850
rect 70364 12404 70420 12798
rect 70476 12404 70532 12414
rect 70364 12402 70532 12404
rect 70364 12350 70478 12402
rect 70530 12350 70532 12402
rect 70364 12348 70532 12350
rect 70476 12338 70532 12348
rect 70812 12292 70868 12302
rect 70812 12198 70868 12236
rect 70252 11218 70308 11228
rect 71260 10948 71316 16492
rect 71708 15148 71764 16830
rect 71820 18676 71876 18686
rect 71820 16548 71876 18620
rect 71820 16482 71876 16492
rect 71932 16100 71988 20860
rect 71932 16034 71988 16044
rect 71260 10882 71316 10892
rect 71372 15092 71764 15148
rect 71820 15092 71876 15102
rect 70140 10658 70196 10668
rect 70476 10724 70532 10734
rect 69916 10500 69972 10510
rect 69580 9214 69582 9266
rect 69634 9214 69636 9266
rect 69580 9202 69636 9214
rect 69804 9940 69860 9950
rect 69804 9266 69860 9884
rect 69804 9214 69806 9266
rect 69858 9214 69860 9266
rect 69804 9202 69860 9214
rect 69244 9044 69300 9054
rect 69244 8930 69300 8988
rect 69916 9044 69972 10444
rect 69916 8950 69972 8988
rect 70364 9044 70420 9054
rect 70364 8950 70420 8988
rect 69244 8878 69246 8930
rect 69298 8878 69300 8930
rect 68832 8652 69096 8662
rect 68888 8596 68936 8652
rect 68992 8596 69040 8652
rect 68832 8586 69096 8596
rect 68460 8530 68516 8540
rect 69244 8484 69300 8878
rect 69244 8418 69300 8428
rect 67116 8372 67172 8382
rect 67116 8278 67172 8316
rect 69804 8034 69860 8046
rect 69804 7982 69806 8034
rect 69858 7982 69860 8034
rect 69804 7812 69860 7982
rect 69580 7756 69860 7812
rect 68908 7362 68964 7374
rect 68908 7310 68910 7362
rect 68962 7310 68964 7362
rect 68908 7252 68964 7310
rect 68908 7186 68964 7196
rect 69244 7362 69300 7374
rect 69244 7310 69246 7362
rect 69298 7310 69300 7362
rect 68832 7084 69096 7094
rect 68888 7028 68936 7084
rect 68992 7028 69040 7084
rect 68832 7018 69096 7028
rect 68684 6578 68740 6590
rect 68684 6526 68686 6578
rect 68738 6526 68740 6578
rect 67340 6468 67396 6478
rect 68684 6468 68740 6526
rect 69020 6580 69076 6590
rect 69020 6486 69076 6524
rect 67340 6466 67620 6468
rect 67340 6414 67342 6466
rect 67394 6414 67620 6466
rect 67340 6412 67620 6414
rect 67340 6402 67396 6412
rect 67116 6132 67172 6142
rect 65884 6076 66052 6132
rect 67004 6130 67172 6132
rect 67004 6078 67118 6130
rect 67170 6078 67172 6130
rect 67004 6076 67172 6078
rect 65884 5908 65940 5918
rect 65884 5814 65940 5852
rect 65772 5030 65828 5068
rect 65548 5012 65604 5022
rect 64764 5010 65044 5012
rect 64764 4958 64766 5010
rect 64818 4958 65044 5010
rect 64764 4956 65044 4958
rect 64764 4946 64820 4956
rect 62860 4732 63588 4788
rect 63532 4226 63588 4732
rect 64988 4340 65044 4956
rect 65548 4918 65604 4956
rect 65996 5012 66052 6076
rect 66332 6020 66388 6030
rect 65996 4946 66052 4956
rect 66108 6018 66388 6020
rect 66108 5966 66334 6018
rect 66386 5966 66388 6018
rect 66108 5964 66388 5966
rect 65996 4452 66052 4462
rect 66108 4452 66164 5964
rect 66332 5954 66388 5964
rect 66668 5906 66724 5918
rect 66668 5854 66670 5906
rect 66722 5854 66724 5906
rect 66668 5346 66724 5854
rect 66668 5294 66670 5346
rect 66722 5294 66724 5346
rect 66668 5282 66724 5294
rect 65996 4450 66164 4452
rect 65996 4398 65998 4450
rect 66050 4398 66164 4450
rect 65996 4396 66164 4398
rect 66332 5122 66388 5134
rect 66332 5070 66334 5122
rect 66386 5070 66388 5122
rect 66332 5012 66388 5070
rect 65996 4386 66052 4396
rect 65212 4340 65268 4350
rect 64988 4338 65268 4340
rect 64988 4286 65214 4338
rect 65266 4286 65268 4338
rect 64988 4284 65268 4286
rect 65212 4274 65268 4284
rect 63532 4174 63534 4226
rect 63586 4174 63588 4226
rect 63532 4162 63588 4174
rect 66332 4228 66388 4956
rect 66332 4162 66388 4172
rect 67116 5012 67172 6076
rect 67564 5348 67620 6412
rect 69244 6468 69300 7310
rect 69580 6692 69636 7756
rect 69804 7700 69860 7756
rect 70364 8034 70420 8046
rect 70364 7982 70366 8034
rect 70418 7982 70420 8034
rect 69916 7700 69972 7710
rect 69804 7644 69916 7700
rect 69916 7634 69972 7644
rect 69692 7588 69748 7598
rect 69692 7586 69860 7588
rect 69692 7534 69694 7586
rect 69746 7534 69860 7586
rect 69692 7532 69860 7534
rect 69692 7522 69748 7532
rect 69580 6626 69636 6636
rect 69692 7252 69748 7262
rect 69692 6804 69748 7196
rect 69692 6690 69748 6748
rect 69692 6638 69694 6690
rect 69746 6638 69748 6690
rect 69692 6626 69748 6638
rect 69356 6468 69412 6478
rect 69244 6412 69356 6468
rect 68684 5908 68740 6412
rect 69356 6374 69412 6412
rect 69804 6468 69860 7532
rect 70364 7586 70420 7982
rect 70364 7534 70366 7586
rect 70418 7534 70420 7586
rect 69916 7476 69972 7486
rect 70364 7476 70420 7534
rect 69916 7474 70420 7476
rect 69916 7422 69918 7474
rect 69970 7422 70420 7474
rect 69916 7420 70420 7422
rect 69916 7364 69972 7420
rect 69916 7298 69972 7308
rect 70476 6580 70532 10668
rect 71372 9940 71428 15092
rect 71820 14532 71876 15036
rect 71820 14438 71876 14476
rect 71708 13748 71764 13758
rect 71708 13654 71764 13692
rect 71372 9846 71428 9884
rect 71708 10612 71764 10622
rect 70700 9828 70756 9838
rect 71708 9828 71764 10556
rect 70700 8260 70756 9772
rect 71484 9826 71764 9828
rect 71484 9774 71710 9826
rect 71762 9774 71764 9826
rect 71484 9772 71764 9774
rect 70476 6514 70532 6524
rect 70588 8258 70756 8260
rect 70588 8206 70702 8258
rect 70754 8206 70756 8258
rect 70588 8204 70756 8206
rect 70028 6468 70084 6478
rect 68684 5842 68740 5852
rect 69580 6244 69636 6254
rect 68460 5796 68516 5806
rect 67564 5292 68404 5348
rect 67228 5124 67284 5134
rect 67228 5030 67284 5068
rect 67564 5122 67620 5292
rect 67564 5070 67566 5122
rect 67618 5070 67620 5122
rect 67564 5058 67620 5070
rect 67900 5124 67956 5134
rect 67900 5030 67956 5068
rect 62412 3602 62468 3612
rect 64764 3668 64820 3678
rect 64764 3574 64820 3612
rect 67116 3666 67172 4956
rect 67676 5012 67732 5022
rect 67676 4918 67732 4956
rect 67116 3614 67118 3666
rect 67170 3614 67172 3666
rect 67116 3602 67172 3614
rect 67900 3556 67956 3566
rect 68012 3556 68068 5292
rect 68348 5122 68404 5292
rect 68460 5234 68516 5740
rect 69356 5796 69412 5806
rect 69356 5702 69412 5740
rect 68832 5516 69096 5526
rect 68888 5460 68936 5516
rect 68992 5460 69040 5516
rect 68832 5450 69096 5460
rect 68460 5182 68462 5234
rect 68514 5182 68516 5234
rect 68460 5170 68516 5182
rect 68348 5070 68350 5122
rect 68402 5070 68404 5122
rect 68348 5058 68404 5070
rect 69020 5124 69076 5134
rect 69020 5030 69076 5068
rect 69580 5122 69636 6188
rect 69580 5070 69582 5122
rect 69634 5070 69636 5122
rect 69580 5058 69636 5070
rect 68572 5012 68628 5022
rect 68460 4956 68572 5012
rect 68124 4228 68180 4238
rect 68124 4134 68180 4172
rect 67900 3554 68068 3556
rect 67900 3502 67902 3554
rect 67954 3502 68068 3554
rect 67900 3500 68068 3502
rect 68236 4116 68292 4126
rect 60620 3442 61012 3444
rect 60620 3390 60622 3442
rect 60674 3390 61012 3442
rect 60620 3388 61012 3390
rect 64092 3444 64148 3482
rect 64316 3444 64372 3454
rect 64092 3442 64372 3444
rect 64092 3390 64094 3442
rect 64146 3390 64318 3442
rect 64370 3390 64372 3442
rect 64092 3388 64372 3390
rect 60620 3378 60676 3388
rect 64092 800 64148 3388
rect 64316 3378 64372 3388
rect 67900 2884 67956 3500
rect 67900 2818 67956 2828
rect 68236 2100 68292 4060
rect 68348 3668 68404 3678
rect 68460 3668 68516 4956
rect 68572 4918 68628 4956
rect 69692 4452 69748 4462
rect 69804 4452 69860 6412
rect 69748 4396 69860 4452
rect 69916 6466 70084 6468
rect 69916 6414 70030 6466
rect 70082 6414 70084 6466
rect 69916 6412 70084 6414
rect 69916 5796 69972 6412
rect 70028 6402 70084 6412
rect 70140 6466 70196 6478
rect 70140 6414 70142 6466
rect 70194 6414 70196 6466
rect 70028 6244 70084 6254
rect 70028 5906 70084 6188
rect 70028 5854 70030 5906
rect 70082 5854 70084 5906
rect 70028 5842 70084 5854
rect 69692 4386 69748 4396
rect 68348 3666 68516 3668
rect 68348 3614 68350 3666
rect 68402 3614 68516 3666
rect 68348 3612 68516 3614
rect 68684 4338 68740 4350
rect 68684 4286 68686 4338
rect 68738 4286 68740 4338
rect 68684 3780 68740 4286
rect 69468 4116 69524 4126
rect 69468 4022 69524 4060
rect 68832 3948 69096 3958
rect 68888 3892 68936 3948
rect 68992 3892 69040 3948
rect 68832 3882 69096 3892
rect 68684 3666 68740 3724
rect 68684 3614 68686 3666
rect 68738 3614 68740 3666
rect 68348 3602 68404 3612
rect 68684 3602 68740 3614
rect 69916 2660 69972 5740
rect 70140 5236 70196 6414
rect 70252 6466 70308 6478
rect 70252 6414 70254 6466
rect 70306 6414 70308 6466
rect 70252 6356 70308 6414
rect 70308 6300 70420 6356
rect 70252 6290 70308 6300
rect 70252 5236 70308 5246
rect 70140 5234 70308 5236
rect 70140 5182 70254 5234
rect 70306 5182 70308 5234
rect 70140 5180 70308 5182
rect 70252 5170 70308 5180
rect 70364 5012 70420 6300
rect 70588 6244 70644 8204
rect 70700 8194 70756 8204
rect 71036 9380 71092 9390
rect 70700 7476 70756 7486
rect 70700 7474 70868 7476
rect 70700 7422 70702 7474
rect 70754 7422 70868 7474
rect 70700 7420 70868 7422
rect 70700 7410 70756 7420
rect 70700 6692 70756 6702
rect 70700 6598 70756 6636
rect 70588 6178 70644 6188
rect 70700 6132 70756 6142
rect 70588 5908 70644 5918
rect 70700 5908 70756 6076
rect 70588 5906 70756 5908
rect 70588 5854 70590 5906
rect 70642 5854 70756 5906
rect 70588 5852 70756 5854
rect 70588 5684 70644 5852
rect 70588 5618 70644 5628
rect 70812 5460 70868 7420
rect 70924 6578 70980 6590
rect 70924 6526 70926 6578
rect 70978 6526 70980 6578
rect 70924 6468 70980 6526
rect 70924 6402 70980 6412
rect 70924 5796 70980 5806
rect 70924 5702 70980 5740
rect 70812 5394 70868 5404
rect 70364 4946 70420 4956
rect 71036 4564 71092 9324
rect 71372 9268 71428 9278
rect 71484 9268 71540 9772
rect 71372 9266 71540 9268
rect 71372 9214 71374 9266
rect 71426 9214 71540 9266
rect 71372 9212 71540 9214
rect 71372 9202 71428 9212
rect 71260 8372 71316 8382
rect 71148 7700 71204 7710
rect 71148 7474 71204 7644
rect 71148 7422 71150 7474
rect 71202 7422 71204 7474
rect 71148 7410 71204 7422
rect 71260 6804 71316 8316
rect 71484 8148 71540 8158
rect 71484 8054 71540 8092
rect 71260 6578 71316 6748
rect 71260 6526 71262 6578
rect 71314 6526 71316 6578
rect 71260 6514 71316 6526
rect 71484 7364 71540 7374
rect 71372 6244 71428 6254
rect 71372 6130 71428 6188
rect 71372 6078 71374 6130
rect 71426 6078 71428 6130
rect 71372 6066 71428 6078
rect 71036 4498 71092 4508
rect 69916 2594 69972 2604
rect 71484 2548 71540 7308
rect 71708 6690 71764 9772
rect 72044 9828 72100 9838
rect 72044 9714 72100 9772
rect 72044 9662 72046 9714
rect 72098 9662 72100 9714
rect 72044 9650 72100 9662
rect 72156 8372 72212 21308
rect 72716 21140 72772 21758
rect 72716 21074 72772 21084
rect 72828 22036 72884 22046
rect 72828 20916 72884 21980
rect 72940 21588 72996 21598
rect 72940 21494 72996 21532
rect 72380 20860 72884 20916
rect 72268 18452 72324 18462
rect 72380 18452 72436 20860
rect 72828 20692 72884 20702
rect 72828 20598 72884 20636
rect 72716 20018 72772 20030
rect 72716 19966 72718 20018
rect 72770 19966 72772 20018
rect 72492 19908 72548 19918
rect 72716 19908 72772 19966
rect 72492 19906 72772 19908
rect 72492 19854 72494 19906
rect 72546 19854 72772 19906
rect 72492 19852 72772 19854
rect 72492 18788 72548 19852
rect 73052 19796 73108 22316
rect 73388 22260 73444 22988
rect 73276 22258 73444 22260
rect 73276 22206 73390 22258
rect 73442 22206 73444 22258
rect 73276 22204 73444 22206
rect 73276 21476 73332 22204
rect 73388 22194 73444 22204
rect 73500 22596 73556 22606
rect 73500 21812 73556 22540
rect 73948 22372 74004 23492
rect 73500 21718 73556 21756
rect 73612 22316 74004 22372
rect 74060 23492 74116 23502
rect 73276 21420 73444 21476
rect 72716 19740 73108 19796
rect 72492 18722 72548 18732
rect 72604 19124 72660 19134
rect 72380 18396 72548 18452
rect 72268 17668 72324 18396
rect 72268 17574 72324 17612
rect 72268 16996 72324 17006
rect 72268 16902 72324 16940
rect 72492 15148 72548 18396
rect 72604 17106 72660 19068
rect 72716 18338 72772 19740
rect 73276 19124 73332 19134
rect 73276 19030 73332 19068
rect 73388 18900 73444 21420
rect 73612 21026 73668 22316
rect 73836 22148 73892 22158
rect 73724 21700 73780 21710
rect 73724 21606 73780 21644
rect 73612 20974 73614 21026
rect 73666 20974 73668 21026
rect 73612 20962 73668 20974
rect 73724 20804 73780 20814
rect 73724 20710 73780 20748
rect 73836 19012 73892 22092
rect 74060 21924 74116 23436
rect 74172 22258 74228 25340
rect 74620 24948 74676 24958
rect 74620 24854 74676 24892
rect 74284 24834 74340 24846
rect 74284 24782 74286 24834
rect 74338 24782 74340 24834
rect 74284 23604 74340 24782
rect 74284 23538 74340 23548
rect 74844 24724 74900 26236
rect 75180 25506 75236 27692
rect 75516 27074 75572 27086
rect 75516 27022 75518 27074
rect 75570 27022 75572 27074
rect 75180 25454 75182 25506
rect 75234 25454 75236 25506
rect 75180 25442 75236 25454
rect 75292 26962 75348 26974
rect 75292 26910 75294 26962
rect 75346 26910 75348 26962
rect 75292 26180 75348 26910
rect 75292 25508 75348 26124
rect 75292 25442 75348 25452
rect 75516 25508 75572 27022
rect 75628 26516 75684 27804
rect 76412 27074 76468 27086
rect 76412 27022 76414 27074
rect 76466 27022 76468 27074
rect 75628 26450 75684 26460
rect 76188 26850 76244 26862
rect 76188 26798 76190 26850
rect 76242 26798 76244 26850
rect 75516 25442 75572 25452
rect 76076 24836 76132 24846
rect 76188 24836 76244 26798
rect 76300 25732 76356 25742
rect 76412 25732 76468 27022
rect 76300 25730 76468 25732
rect 76300 25678 76302 25730
rect 76354 25678 76468 25730
rect 76300 25676 76468 25678
rect 76300 25666 76356 25676
rect 76524 25620 76580 29036
rect 76636 25732 76692 25742
rect 76636 25638 76692 25676
rect 76076 24834 76244 24836
rect 76076 24782 76078 24834
rect 76130 24782 76244 24834
rect 76076 24780 76244 24782
rect 76412 25564 76580 25620
rect 76972 25620 77028 29932
rect 77084 26180 77140 26190
rect 77084 26086 77140 26124
rect 77308 25732 77364 30268
rect 77980 30324 78036 30334
rect 77980 30210 78036 30268
rect 77980 30158 77982 30210
rect 78034 30158 78036 30210
rect 77980 30146 78036 30158
rect 77420 30098 77476 30110
rect 77420 30046 77422 30098
rect 77474 30046 77476 30098
rect 77420 29316 77476 30046
rect 78492 29820 78756 29830
rect 78548 29764 78596 29820
rect 78652 29764 78700 29820
rect 78492 29754 78756 29764
rect 77756 29316 77812 29326
rect 77420 29314 77812 29316
rect 77420 29262 77758 29314
rect 77810 29262 77812 29314
rect 77420 29260 77812 29262
rect 77756 26964 77812 29260
rect 78492 28252 78756 28262
rect 78548 28196 78596 28252
rect 78652 28196 78700 28252
rect 78492 28186 78756 28196
rect 77756 26898 77812 26908
rect 77980 27634 78036 27646
rect 77980 27582 77982 27634
rect 78034 27582 78036 27634
rect 77980 26068 78036 27582
rect 78492 26684 78756 26694
rect 78548 26628 78596 26684
rect 78652 26628 78700 26684
rect 78492 26618 78756 26628
rect 77980 26002 78036 26012
rect 77308 25666 77364 25676
rect 77980 25732 78036 25742
rect 76972 25564 77140 25620
rect 76076 24770 76132 24780
rect 75292 24724 75348 24734
rect 74844 24722 75348 24724
rect 74844 24670 75294 24722
rect 75346 24670 75348 24722
rect 74844 24668 75348 24670
rect 74844 23492 74900 24668
rect 75292 24658 75348 24668
rect 75404 24050 75460 24062
rect 75404 23998 75406 24050
rect 75458 23998 75460 24050
rect 75404 23716 75460 23998
rect 75404 23650 75460 23660
rect 76412 23492 76468 25564
rect 76860 25508 76916 25518
rect 76860 25394 76916 25452
rect 76860 25342 76862 25394
rect 76914 25342 76916 25394
rect 76524 23716 76580 23726
rect 76524 23714 76692 23716
rect 76524 23662 76526 23714
rect 76578 23662 76692 23714
rect 76524 23660 76692 23662
rect 76524 23650 76580 23660
rect 76412 23436 76580 23492
rect 74844 23426 74900 23436
rect 74284 23044 74340 23054
rect 76412 23044 76468 23054
rect 74284 23042 74452 23044
rect 74284 22990 74286 23042
rect 74338 22990 74452 23042
rect 74284 22988 74452 22990
rect 74284 22978 74340 22988
rect 74172 22206 74174 22258
rect 74226 22206 74228 22258
rect 74172 22148 74228 22206
rect 74172 22082 74228 22092
rect 74060 21810 74116 21868
rect 74060 21758 74062 21810
rect 74114 21758 74116 21810
rect 74060 21746 74116 21758
rect 74396 21810 74452 22988
rect 76412 22950 76468 22988
rect 75628 22820 75684 22830
rect 75628 22482 75684 22764
rect 75628 22430 75630 22482
rect 75682 22430 75684 22482
rect 75628 22418 75684 22430
rect 74844 22370 74900 22382
rect 74844 22318 74846 22370
rect 74898 22318 74900 22370
rect 74844 22036 74900 22318
rect 74844 21970 74900 21980
rect 75068 22146 75124 22158
rect 75068 22094 75070 22146
rect 75122 22094 75124 22146
rect 74396 21758 74398 21810
rect 74450 21758 74452 21810
rect 74396 21746 74452 21758
rect 74732 21812 74788 21822
rect 74732 21698 74788 21756
rect 74732 21646 74734 21698
rect 74786 21646 74788 21698
rect 74732 21634 74788 21646
rect 74844 21588 74900 21598
rect 73948 21476 74004 21486
rect 74004 21420 74116 21476
rect 73948 21410 74004 21420
rect 73164 18844 73444 18900
rect 73724 18956 73892 19012
rect 73948 19234 74004 19246
rect 73948 19182 73950 19234
rect 74002 19182 74004 19234
rect 72716 18286 72718 18338
rect 72770 18286 72772 18338
rect 72716 18274 72772 18286
rect 72828 18562 72884 18574
rect 72828 18510 72830 18562
rect 72882 18510 72884 18562
rect 72604 17054 72606 17106
rect 72658 17054 72660 17106
rect 72604 17042 72660 17054
rect 72828 17108 72884 18510
rect 73052 18450 73108 18462
rect 73052 18398 73054 18450
rect 73106 18398 73108 18450
rect 73052 17778 73108 18398
rect 73052 17726 73054 17778
rect 73106 17726 73108 17778
rect 73052 17714 73108 17726
rect 73164 17556 73220 18844
rect 73164 17490 73220 17500
rect 73388 17892 73444 17902
rect 72828 17042 72884 17052
rect 73164 15204 73220 15214
rect 72492 15092 72772 15148
rect 72268 14306 72324 14318
rect 72268 14254 72270 14306
rect 72322 14254 72324 14306
rect 72268 13748 72324 14254
rect 72492 13748 72548 13758
rect 72716 13748 72772 15092
rect 72268 13692 72492 13748
rect 72492 13682 72548 13692
rect 72604 13746 72772 13748
rect 72604 13694 72718 13746
rect 72770 13694 72772 13746
rect 72604 13692 72772 13694
rect 72380 13522 72436 13534
rect 72380 13470 72382 13522
rect 72434 13470 72436 13522
rect 72380 12292 72436 13470
rect 72604 13074 72660 13692
rect 72716 13682 72772 13692
rect 72604 13022 72606 13074
rect 72658 13022 72660 13074
rect 72604 13010 72660 13022
rect 73164 12962 73220 15148
rect 73388 13972 73444 17836
rect 73724 17554 73780 18956
rect 73948 18900 74004 19182
rect 73836 18844 74004 18900
rect 73836 18228 73892 18844
rect 73948 18676 74004 18686
rect 73948 18450 74004 18620
rect 73948 18398 73950 18450
rect 74002 18398 74004 18450
rect 73948 18386 74004 18398
rect 73836 18172 74004 18228
rect 73724 17502 73726 17554
rect 73778 17502 73780 17554
rect 73724 16324 73780 17502
rect 73724 16258 73780 16268
rect 73836 16100 73892 16110
rect 73836 16006 73892 16044
rect 73948 15540 74004 18172
rect 73500 15484 74004 15540
rect 73500 15092 73556 15484
rect 73948 15316 74004 15326
rect 74060 15316 74116 21420
rect 74172 20578 74228 20590
rect 74172 20526 74174 20578
rect 74226 20526 74228 20578
rect 74172 20188 74228 20526
rect 74172 20132 74452 20188
rect 74396 19010 74452 20132
rect 74396 18958 74398 19010
rect 74450 18958 74452 19010
rect 74396 18228 74452 18958
rect 74396 18162 74452 18172
rect 74620 17666 74676 17678
rect 74620 17614 74622 17666
rect 74674 17614 74676 17666
rect 74620 17444 74676 17614
rect 74620 16884 74676 17388
rect 74396 16100 74452 16110
rect 74396 16006 74452 16044
rect 74172 15874 74228 15886
rect 74172 15822 74174 15874
rect 74226 15822 74228 15874
rect 74172 15540 74228 15822
rect 74172 15484 74564 15540
rect 74508 15426 74564 15484
rect 74508 15374 74510 15426
rect 74562 15374 74564 15426
rect 73948 15314 74060 15316
rect 73948 15262 73950 15314
rect 74002 15262 74060 15314
rect 73948 15260 74060 15262
rect 73948 15250 74004 15260
rect 74060 15222 74116 15260
rect 74396 15314 74452 15326
rect 74396 15262 74398 15314
rect 74450 15262 74452 15314
rect 74396 15204 74452 15262
rect 74396 15138 74452 15148
rect 73500 15026 73556 15036
rect 73612 15090 73668 15102
rect 73612 15038 73614 15090
rect 73666 15038 73668 15090
rect 73612 14420 73668 15038
rect 74172 14980 74228 14990
rect 73612 14364 74116 14420
rect 73388 13916 73668 13972
rect 73276 13860 73332 13870
rect 73276 13766 73332 13804
rect 73164 12910 73166 12962
rect 73218 12910 73220 12962
rect 73164 12898 73220 12910
rect 73388 13748 73444 13758
rect 72380 12226 72436 12236
rect 72940 12850 72996 12862
rect 72940 12798 72942 12850
rect 72994 12798 72996 12850
rect 72492 11282 72548 11294
rect 72492 11230 72494 11282
rect 72546 11230 72548 11282
rect 72268 11172 72324 11182
rect 72492 11172 72548 11230
rect 72604 11284 72660 11294
rect 72660 11228 72772 11284
rect 72604 11190 72660 11228
rect 72268 11170 72548 11172
rect 72268 11118 72270 11170
rect 72322 11118 72548 11170
rect 72268 11116 72548 11118
rect 72268 9380 72324 11116
rect 72268 9314 72324 9324
rect 72380 10948 72436 10958
rect 72380 10164 72436 10892
rect 72604 10724 72660 10734
rect 72604 10610 72660 10668
rect 72604 10558 72606 10610
rect 72658 10558 72660 10610
rect 72604 10546 72660 10558
rect 72716 10500 72772 11228
rect 72716 10434 72772 10444
rect 72828 11170 72884 11182
rect 72828 11118 72830 11170
rect 72882 11118 72884 11170
rect 72380 9266 72436 10108
rect 72380 9214 72382 9266
rect 72434 9214 72436 9266
rect 72380 9202 72436 9214
rect 72492 9828 72548 9838
rect 72156 8306 72212 8316
rect 72268 9042 72324 9054
rect 72268 8990 72270 9042
rect 72322 8990 72324 9042
rect 72268 7474 72324 8990
rect 72380 8148 72436 8158
rect 72380 7698 72436 8092
rect 72380 7646 72382 7698
rect 72434 7646 72436 7698
rect 72380 7634 72436 7646
rect 72492 7698 72548 9772
rect 72828 9826 72884 11118
rect 72828 9774 72830 9826
rect 72882 9774 72884 9826
rect 72828 9762 72884 9774
rect 72940 10052 72996 12798
rect 73276 12740 73332 12750
rect 73164 12684 73276 12740
rect 72940 9716 72996 9996
rect 72940 9650 72996 9660
rect 73052 12628 73108 12638
rect 72604 9044 72660 9054
rect 72604 9042 72772 9044
rect 72604 8990 72606 9042
rect 72658 8990 72772 9042
rect 72604 8988 72772 8990
rect 72604 8978 72660 8988
rect 72492 7646 72494 7698
rect 72546 7646 72548 7698
rect 72492 7634 72548 7646
rect 72716 7698 72772 8988
rect 72716 7646 72718 7698
rect 72770 7646 72772 7698
rect 72716 7634 72772 7646
rect 72940 8930 72996 8942
rect 72940 8878 72942 8930
rect 72994 8878 72996 8930
rect 72268 7422 72270 7474
rect 72322 7422 72324 7474
rect 72268 7364 72324 7422
rect 72268 7298 72324 7308
rect 72940 7364 72996 8878
rect 72940 7298 72996 7308
rect 73052 7140 73108 12572
rect 73164 7700 73220 12684
rect 73276 12646 73332 12684
rect 73388 10724 73444 13692
rect 73388 10658 73444 10668
rect 73388 10498 73444 10510
rect 73612 10500 73668 13916
rect 73724 13860 73780 13870
rect 73724 12850 73780 13804
rect 74060 13858 74116 14364
rect 74060 13806 74062 13858
rect 74114 13806 74116 13858
rect 74060 13794 74116 13806
rect 73948 12964 74004 12974
rect 73948 12870 74004 12908
rect 73724 12798 73726 12850
rect 73778 12798 73780 12850
rect 73724 12786 73780 12798
rect 74172 12628 74228 14924
rect 74508 14084 74564 15374
rect 74620 14980 74676 16828
rect 74620 14914 74676 14924
rect 74732 15316 74788 15326
rect 74508 14018 74564 14028
rect 74620 14306 74676 14318
rect 74620 14254 74622 14306
rect 74674 14254 74676 14306
rect 74620 13972 74676 14254
rect 74620 13906 74676 13916
rect 74396 13860 74452 13870
rect 74396 13766 74452 13804
rect 74732 13634 74788 15260
rect 74732 13582 74734 13634
rect 74786 13582 74788 13634
rect 74732 13570 74788 13582
rect 74844 13412 74900 21532
rect 75068 20804 75124 22094
rect 76300 22146 76356 22158
rect 76300 22094 76302 22146
rect 76354 22094 76356 22146
rect 75180 21924 75236 21934
rect 75180 21586 75236 21868
rect 76300 21812 76356 22094
rect 76300 21746 76356 21756
rect 75852 21700 75908 21710
rect 75852 21606 75908 21644
rect 75180 21534 75182 21586
rect 75234 21534 75236 21586
rect 75180 21522 75236 21534
rect 75068 20738 75124 20748
rect 75292 20578 75348 20590
rect 75292 20526 75294 20578
rect 75346 20526 75348 20578
rect 75292 20244 75348 20526
rect 76300 20578 76356 20590
rect 76300 20526 76302 20578
rect 76354 20526 76356 20578
rect 75292 20178 75348 20188
rect 75740 20244 75796 20254
rect 76300 20188 76356 20526
rect 75740 20018 75796 20188
rect 75740 19966 75742 20018
rect 75794 19966 75796 20018
rect 75740 19954 75796 19966
rect 76188 20132 76356 20188
rect 75068 19794 75124 19806
rect 75068 19742 75070 19794
rect 75122 19742 75124 19794
rect 74956 19348 75012 19358
rect 74956 19254 75012 19292
rect 75068 18676 75124 19742
rect 76188 19460 76244 20132
rect 76188 19234 76244 19404
rect 76188 19182 76190 19234
rect 76242 19182 76244 19234
rect 76188 19170 76244 19182
rect 75628 19124 75684 19134
rect 75628 19030 75684 19068
rect 75292 19012 75348 19022
rect 75292 18918 75348 18956
rect 75516 19010 75572 19022
rect 75516 18958 75518 19010
rect 75570 18958 75572 19010
rect 75068 18610 75124 18620
rect 75292 18452 75348 18462
rect 75516 18452 75572 18958
rect 75348 18396 75572 18452
rect 75292 18338 75348 18396
rect 75292 18286 75294 18338
rect 75346 18286 75348 18338
rect 75292 18274 75348 18286
rect 76412 17892 76468 17902
rect 75516 17780 75572 17790
rect 75516 17686 75572 17724
rect 74956 17668 75012 17678
rect 74956 16770 75012 17612
rect 76412 17666 76468 17836
rect 76412 17614 76414 17666
rect 76466 17614 76468 17666
rect 76412 17602 76468 17614
rect 75180 17444 75236 17454
rect 75180 17350 75236 17388
rect 75628 17444 75684 17454
rect 76188 17444 76244 17454
rect 75628 17442 76188 17444
rect 75628 17390 75630 17442
rect 75682 17390 76188 17442
rect 75628 17388 76188 17390
rect 75628 17378 75684 17388
rect 76188 17350 76244 17388
rect 76300 17442 76356 17454
rect 76300 17390 76302 17442
rect 76354 17390 76356 17442
rect 76300 17108 76356 17390
rect 76524 17220 76580 23436
rect 76636 22820 76692 23660
rect 76860 23156 76916 25342
rect 76636 22594 76692 22764
rect 76636 22542 76638 22594
rect 76690 22542 76692 22594
rect 76636 22530 76692 22542
rect 76748 23154 76916 23156
rect 76748 23102 76862 23154
rect 76914 23102 76916 23154
rect 76748 23100 76916 23102
rect 76748 20188 76804 23100
rect 76860 23090 76916 23100
rect 76972 23266 77028 23278
rect 76972 23214 76974 23266
rect 77026 23214 77028 23266
rect 76972 22708 77028 23214
rect 76972 22642 77028 22652
rect 76636 20132 76804 20188
rect 76860 22260 76916 22270
rect 77084 22260 77140 25564
rect 77980 25618 78036 25676
rect 77980 25566 77982 25618
rect 78034 25566 78036 25618
rect 77980 25554 78036 25566
rect 77420 25396 77476 25406
rect 77420 25302 77476 25340
rect 78204 25396 78260 25406
rect 78204 24610 78260 25340
rect 78492 25116 78756 25126
rect 78548 25060 78596 25116
rect 78652 25060 78700 25116
rect 78492 25050 78756 25060
rect 78204 24558 78206 24610
rect 78258 24558 78260 24610
rect 78204 24546 78260 24558
rect 78492 23548 78756 23558
rect 78548 23492 78596 23548
rect 78652 23492 78700 23548
rect 78492 23482 78756 23492
rect 76860 22258 77140 22260
rect 76860 22206 76862 22258
rect 76914 22206 77140 22258
rect 76860 22204 77140 22206
rect 77196 23044 77252 23054
rect 77196 22258 77252 22988
rect 77644 22930 77700 22942
rect 77644 22878 77646 22930
rect 77698 22878 77700 22930
rect 77644 22820 77700 22878
rect 77980 22932 78036 22942
rect 77980 22930 78148 22932
rect 77980 22878 77982 22930
rect 78034 22878 78148 22930
rect 77980 22876 78148 22878
rect 77980 22866 78036 22876
rect 77644 22754 77700 22764
rect 77196 22206 77198 22258
rect 77250 22206 77252 22258
rect 76636 19346 76692 20132
rect 76636 19294 76638 19346
rect 76690 19294 76692 19346
rect 76636 17780 76692 19294
rect 76860 19348 76916 22204
rect 77196 22194 77252 22206
rect 77980 22708 78036 22718
rect 77868 22146 77924 22158
rect 77868 22094 77870 22146
rect 77922 22094 77924 22146
rect 77868 21700 77924 22094
rect 77868 21634 77924 21644
rect 77980 21474 78036 22652
rect 78092 22370 78148 22876
rect 78092 22318 78094 22370
rect 78146 22318 78148 22370
rect 78092 22306 78148 22318
rect 78492 21980 78756 21990
rect 78548 21924 78596 21980
rect 78652 21924 78700 21980
rect 78492 21914 78756 21924
rect 77980 21422 77982 21474
rect 78034 21422 78036 21474
rect 77980 21410 78036 21422
rect 77980 21140 78036 21150
rect 77980 19906 78036 21084
rect 78492 20412 78756 20422
rect 78548 20356 78596 20412
rect 78652 20356 78700 20412
rect 78492 20346 78756 20356
rect 77980 19854 77982 19906
rect 78034 19854 78036 19906
rect 77980 19842 78036 19854
rect 76860 19282 76916 19292
rect 78092 19348 78148 19358
rect 78092 19254 78148 19292
rect 77644 19124 77700 19134
rect 77980 19124 78036 19134
rect 77700 19122 78036 19124
rect 77700 19070 77982 19122
rect 78034 19070 78036 19122
rect 77700 19068 78036 19070
rect 77644 19030 77700 19068
rect 77980 19058 78036 19068
rect 77196 19012 77252 19022
rect 77420 19012 77476 19022
rect 77196 18918 77252 18956
rect 77308 19010 77476 19012
rect 77308 18958 77422 19010
rect 77474 18958 77476 19010
rect 77308 18956 77476 18958
rect 77308 17892 77364 18956
rect 77420 18946 77476 18956
rect 77532 19010 77588 19022
rect 77532 18958 77534 19010
rect 77586 18958 77588 19010
rect 77420 18564 77476 18574
rect 77532 18564 77588 18958
rect 78492 18844 78756 18854
rect 78548 18788 78596 18844
rect 78652 18788 78700 18844
rect 78492 18778 78756 18788
rect 77420 18562 77588 18564
rect 77420 18510 77422 18562
rect 77474 18510 77588 18562
rect 77420 18508 77588 18510
rect 77420 18498 77476 18508
rect 78092 18452 78148 18462
rect 77308 17826 77364 17836
rect 77868 18450 78148 18452
rect 77868 18398 78094 18450
rect 78146 18398 78148 18450
rect 77868 18396 78148 18398
rect 76636 17714 76692 17724
rect 76748 17668 76804 17678
rect 76972 17668 77028 17678
rect 76748 17666 77028 17668
rect 76748 17614 76750 17666
rect 76802 17614 76974 17666
rect 77026 17614 77028 17666
rect 76748 17612 77028 17614
rect 76748 17602 76804 17612
rect 76972 17602 77028 17612
rect 77196 17668 77252 17678
rect 77196 17554 77252 17612
rect 77196 17502 77198 17554
rect 77250 17502 77252 17554
rect 77196 17490 77252 17502
rect 77308 17554 77364 17566
rect 77308 17502 77310 17554
rect 77362 17502 77364 17554
rect 77308 17444 77364 17502
rect 77308 17378 77364 17388
rect 76524 17164 77252 17220
rect 76300 17052 77140 17108
rect 77084 16994 77140 17052
rect 77084 16942 77086 16994
rect 77138 16942 77140 16994
rect 77084 16930 77140 16942
rect 77196 16772 77252 17164
rect 77868 16884 77924 18396
rect 78092 18386 78148 18396
rect 78492 17276 78756 17286
rect 78548 17220 78596 17276
rect 78652 17220 78700 17276
rect 78492 17210 78756 17220
rect 74956 16718 74958 16770
rect 75010 16718 75012 16770
rect 74956 16706 75012 16718
rect 77084 16716 77252 16772
rect 77756 16882 77924 16884
rect 77756 16830 77870 16882
rect 77922 16830 77924 16882
rect 77756 16828 77924 16830
rect 76412 16212 76468 16222
rect 76412 16118 76468 16156
rect 76972 16212 77028 16222
rect 76972 16098 77028 16156
rect 76972 16046 76974 16098
rect 77026 16046 77028 16098
rect 76972 16034 77028 16046
rect 76748 15876 76804 15886
rect 76524 15874 76804 15876
rect 76524 15822 76750 15874
rect 76802 15822 76804 15874
rect 76524 15820 76804 15822
rect 76524 15540 76580 15820
rect 76748 15810 76804 15820
rect 76076 15484 76580 15540
rect 76076 15314 76132 15484
rect 76076 15262 76078 15314
rect 76130 15262 76132 15314
rect 76076 15250 76132 15262
rect 76188 15092 76244 15102
rect 75628 14532 75684 14542
rect 75628 14438 75684 14476
rect 76188 14530 76244 15036
rect 76188 14478 76190 14530
rect 76242 14478 76244 14530
rect 76188 14466 76244 14478
rect 76860 14532 76916 14542
rect 74508 13356 74900 13412
rect 76300 14420 76356 14430
rect 74508 13186 74564 13356
rect 74508 13134 74510 13186
rect 74562 13134 74564 13186
rect 74508 13122 74564 13134
rect 74172 12562 74228 12572
rect 74732 12068 74788 13356
rect 74844 12852 74900 12862
rect 75292 12852 75348 12862
rect 74844 12850 75348 12852
rect 74844 12798 74846 12850
rect 74898 12798 75294 12850
rect 75346 12798 75348 12850
rect 74844 12796 75348 12798
rect 74844 12786 74900 12796
rect 75292 12786 75348 12796
rect 75628 12740 75684 12750
rect 75628 12646 75684 12684
rect 74956 12068 75012 12078
rect 74732 12066 75012 12068
rect 74732 12014 74958 12066
rect 75010 12014 75012 12066
rect 74732 12012 75012 12014
rect 74956 12002 75012 12012
rect 75628 11396 75684 11406
rect 75628 11302 75684 11340
rect 74620 11172 74676 11182
rect 74620 11078 74676 11116
rect 73388 10446 73390 10498
rect 73442 10446 73444 10498
rect 73388 10276 73444 10446
rect 73388 10210 73444 10220
rect 73500 10444 73668 10500
rect 74172 10724 74228 10734
rect 73500 9828 73556 10444
rect 74060 10276 74116 10286
rect 73612 10164 73668 10174
rect 73668 10108 73780 10164
rect 73612 10098 73668 10108
rect 73500 9734 73556 9772
rect 73612 9940 73668 9950
rect 73276 9602 73332 9614
rect 73276 9550 73278 9602
rect 73330 9550 73332 9602
rect 73276 9380 73332 9550
rect 73388 9604 73444 9614
rect 73388 9602 73556 9604
rect 73388 9550 73390 9602
rect 73442 9550 73556 9602
rect 73388 9548 73556 9550
rect 73388 9538 73444 9548
rect 73500 9492 73556 9548
rect 73500 9426 73556 9436
rect 73276 9314 73332 9324
rect 73612 9266 73668 9884
rect 73612 9214 73614 9266
rect 73666 9214 73668 9266
rect 73612 9202 73668 9214
rect 73612 8372 73668 8382
rect 73724 8372 73780 10108
rect 73836 9716 73892 9726
rect 73836 9714 74004 9716
rect 73836 9662 73838 9714
rect 73890 9662 74004 9714
rect 73836 9660 74004 9662
rect 73836 9380 73892 9660
rect 73836 9314 73892 9324
rect 73948 9266 74004 9660
rect 74060 9492 74116 10220
rect 74060 9426 74116 9436
rect 73948 9214 73950 9266
rect 74002 9214 74004 9266
rect 73948 9202 74004 9214
rect 73612 8370 73780 8372
rect 73612 8318 73614 8370
rect 73666 8318 73780 8370
rect 73612 8316 73780 8318
rect 73612 8306 73668 8316
rect 73164 7634 73220 7644
rect 73276 7364 73332 7374
rect 73276 7270 73332 7308
rect 72380 7084 73444 7140
rect 71708 6638 71710 6690
rect 71762 6638 71764 6690
rect 71596 6580 71652 6590
rect 71596 5906 71652 6524
rect 71708 6356 71764 6638
rect 71708 6290 71764 6300
rect 72156 6692 72212 6702
rect 72156 6130 72212 6636
rect 72156 6078 72158 6130
rect 72210 6078 72212 6130
rect 72156 6066 72212 6078
rect 72268 6466 72324 6478
rect 72268 6414 72270 6466
rect 72322 6414 72324 6466
rect 71596 5854 71598 5906
rect 71650 5854 71652 5906
rect 71596 5842 71652 5854
rect 72268 5796 72324 6414
rect 72380 6130 72436 7084
rect 72380 6078 72382 6130
rect 72434 6078 72436 6130
rect 72380 6066 72436 6078
rect 72604 6466 72660 6478
rect 72604 6414 72606 6466
rect 72658 6414 72660 6466
rect 72492 5908 72548 5918
rect 72604 5908 72660 6414
rect 72492 5906 72660 5908
rect 72492 5854 72494 5906
rect 72546 5854 72660 5906
rect 72492 5852 72660 5854
rect 72492 5796 72548 5852
rect 72324 5740 72548 5796
rect 72268 5730 72324 5740
rect 72716 5684 72772 7084
rect 72940 6132 72996 6142
rect 72940 6038 72996 6076
rect 73388 6130 73444 7084
rect 73388 6078 73390 6130
rect 73442 6078 73444 6130
rect 73388 6066 73444 6078
rect 74172 6132 74228 10668
rect 75516 10500 75572 10510
rect 75516 10406 75572 10444
rect 76076 10498 76132 10510
rect 76076 10446 76078 10498
rect 76130 10446 76132 10498
rect 75740 10388 75796 10398
rect 75628 10386 75796 10388
rect 75628 10334 75742 10386
rect 75794 10334 75796 10386
rect 75628 10332 75796 10334
rect 74284 10052 74340 10062
rect 74284 9826 74340 9996
rect 74284 9774 74286 9826
rect 74338 9774 74340 9826
rect 74284 9762 74340 9774
rect 74172 6066 74228 6076
rect 72492 5628 72772 5684
rect 72380 5460 72436 5470
rect 71484 2482 71540 2492
rect 72156 3556 72212 3566
rect 72156 3442 72212 3500
rect 72156 3390 72158 3442
rect 72210 3390 72212 3442
rect 68124 2044 68292 2100
rect 68124 800 68180 2044
rect 72156 800 72212 3390
rect 72380 3330 72436 5404
rect 72492 5234 72548 5628
rect 72492 5182 72494 5234
rect 72546 5182 72548 5234
rect 72492 5170 72548 5182
rect 75628 4338 75684 10332
rect 75740 10322 75796 10332
rect 76076 10388 76132 10446
rect 76076 10322 76132 10332
rect 76300 9604 76356 14364
rect 76860 14418 76916 14476
rect 76860 14366 76862 14418
rect 76914 14366 76916 14418
rect 76860 14354 76916 14366
rect 76524 14308 76580 14318
rect 76524 14214 76580 14252
rect 76860 13860 76916 13870
rect 76860 13766 76916 13804
rect 77084 12852 77140 16716
rect 77196 14420 77252 14430
rect 77196 14326 77252 14364
rect 77644 14420 77700 14430
rect 77644 14326 77700 14364
rect 77756 14308 77812 16828
rect 77868 16818 77924 16828
rect 77980 16212 78036 16222
rect 77980 15202 78036 16156
rect 78492 15708 78756 15718
rect 78548 15652 78596 15708
rect 78652 15652 78700 15708
rect 78492 15642 78756 15652
rect 77980 15150 77982 15202
rect 78034 15150 78036 15202
rect 77980 15138 78036 15150
rect 77644 13748 77700 13758
rect 77756 13748 77812 14252
rect 78492 14140 78756 14150
rect 78548 14084 78596 14140
rect 78652 14084 78700 14140
rect 78492 14074 78756 14084
rect 77644 13746 77812 13748
rect 77644 13694 77646 13746
rect 77698 13694 77812 13746
rect 77644 13692 77812 13694
rect 77644 13682 77700 13692
rect 77084 12796 77252 12852
rect 76860 12740 76916 12750
rect 76916 12684 77140 12740
rect 76860 12674 76916 12684
rect 77084 12290 77140 12684
rect 77084 12238 77086 12290
rect 77138 12238 77140 12290
rect 77084 12226 77140 12238
rect 76524 11620 76580 11630
rect 76412 11170 76468 11182
rect 76412 11118 76414 11170
rect 76466 11118 76468 11170
rect 76412 10836 76468 11118
rect 76412 10770 76468 10780
rect 76524 10948 76580 11564
rect 76748 11396 76804 11406
rect 76748 11282 76804 11340
rect 76748 11230 76750 11282
rect 76802 11230 76804 11282
rect 76748 11218 76804 11230
rect 77084 11282 77140 11294
rect 77084 11230 77086 11282
rect 77138 11230 77140 11282
rect 76524 10892 76916 10948
rect 76524 10834 76580 10892
rect 76524 10782 76526 10834
rect 76578 10782 76580 10834
rect 76524 10770 76580 10782
rect 76748 10724 76804 10734
rect 76636 10722 76804 10724
rect 76636 10670 76750 10722
rect 76802 10670 76804 10722
rect 76636 10668 76804 10670
rect 76524 10388 76580 10398
rect 76636 10388 76692 10668
rect 76748 10658 76804 10668
rect 76860 10612 76916 10892
rect 76972 10836 77028 10846
rect 77084 10836 77140 11230
rect 77028 10780 77140 10836
rect 76972 10770 77028 10780
rect 76972 10612 77028 10622
rect 76860 10610 77028 10612
rect 76860 10558 76974 10610
rect 77026 10558 77028 10610
rect 76860 10556 77028 10558
rect 76972 10546 77028 10556
rect 76524 10386 76692 10388
rect 76524 10334 76526 10386
rect 76578 10334 76692 10386
rect 76524 10332 76692 10334
rect 76524 10322 76580 10332
rect 76412 9828 76468 9838
rect 76412 9826 76916 9828
rect 76412 9774 76414 9826
rect 76466 9774 76916 9826
rect 76412 9772 76916 9774
rect 76412 9762 76468 9772
rect 76860 9716 76916 9772
rect 77084 9716 77140 9726
rect 76860 9714 77140 9716
rect 76860 9662 77086 9714
rect 77138 9662 77140 9714
rect 76860 9660 77140 9662
rect 76748 9604 76804 9614
rect 76300 9538 76356 9548
rect 76524 9602 76804 9604
rect 76524 9550 76750 9602
rect 76802 9550 76804 9602
rect 76524 9548 76804 9550
rect 76524 9268 76580 9548
rect 76748 9538 76804 9548
rect 76076 9212 76580 9268
rect 76076 9042 76132 9212
rect 76076 8990 76078 9042
rect 76130 8990 76132 9042
rect 76076 8978 76132 8990
rect 76972 7924 77028 7934
rect 76748 7588 76804 7598
rect 76076 7586 76804 7588
rect 76076 7534 76750 7586
rect 76802 7534 76804 7586
rect 76076 7532 76804 7534
rect 76076 5906 76132 7532
rect 76748 7522 76804 7532
rect 76972 7476 77028 7868
rect 76860 7474 77028 7476
rect 76860 7422 76974 7474
rect 77026 7422 77028 7474
rect 76860 7420 77028 7422
rect 76524 7364 76580 7374
rect 76860 7364 76916 7420
rect 76972 7410 77028 7420
rect 76524 7362 76916 7364
rect 76524 7310 76526 7362
rect 76578 7310 76916 7362
rect 76524 7308 76916 7310
rect 76524 7298 76580 7308
rect 76076 5854 76078 5906
rect 76130 5854 76132 5906
rect 76076 5842 76132 5854
rect 76972 7252 77028 7262
rect 76972 5234 77028 7196
rect 76972 5182 76974 5234
rect 77026 5182 77028 5234
rect 76972 5170 77028 5182
rect 75740 5124 75796 5134
rect 76412 5124 76468 5134
rect 75740 5122 76468 5124
rect 75740 5070 75742 5122
rect 75794 5070 76414 5122
rect 76466 5070 76468 5122
rect 75740 5068 76468 5070
rect 75740 5058 75796 5068
rect 75628 4286 75630 4338
rect 75682 4286 75684 4338
rect 75628 4274 75684 4286
rect 72604 3556 72660 3566
rect 72604 3462 72660 3500
rect 72380 3278 72382 3330
rect 72434 3278 72436 3330
rect 72380 3266 72436 3278
rect 75516 3442 75572 3454
rect 75516 3390 75518 3442
rect 75570 3390 75572 3442
rect 75516 1428 75572 3390
rect 76412 3388 76468 5068
rect 75516 1362 75572 1372
rect 76188 3332 76468 3388
rect 77084 3332 77140 9660
rect 77196 7364 77252 12796
rect 77756 12178 77812 13692
rect 78492 12572 78756 12582
rect 78548 12516 78596 12572
rect 78652 12516 78700 12572
rect 78492 12506 78756 12516
rect 77756 12126 77758 12178
rect 77810 12126 77812 12178
rect 77756 12114 77812 12126
rect 78492 11004 78756 11014
rect 78548 10948 78596 11004
rect 78652 10948 78700 11004
rect 78492 10938 78756 10948
rect 77420 10724 77476 10734
rect 77196 7298 77252 7308
rect 77308 10722 77476 10724
rect 77308 10670 77422 10722
rect 77474 10670 77476 10722
rect 77308 10668 77476 10670
rect 77308 7140 77364 10668
rect 77420 10658 77476 10668
rect 77644 10610 77700 10622
rect 77644 10558 77646 10610
rect 77698 10558 77700 10610
rect 77644 10388 77700 10558
rect 77644 10322 77700 10332
rect 78492 9436 78756 9446
rect 78548 9380 78596 9436
rect 78652 9380 78700 9436
rect 78492 9370 78756 9380
rect 77980 8820 78036 8830
rect 77980 8726 78036 8764
rect 78492 7868 78756 7878
rect 78548 7812 78596 7868
rect 78652 7812 78700 7868
rect 78492 7802 78756 7812
rect 77196 7084 77364 7140
rect 77196 3554 77252 7084
rect 78492 6300 78756 6310
rect 78548 6244 78596 6300
rect 78652 6244 78700 6300
rect 78492 6234 78756 6244
rect 77980 6132 78036 6142
rect 77980 5794 78036 6076
rect 77980 5742 77982 5794
rect 78034 5742 78036 5794
rect 77980 5730 78036 5742
rect 78492 4732 78756 4742
rect 78548 4676 78596 4732
rect 78652 4676 78700 4732
rect 78492 4666 78756 4676
rect 77980 4114 78036 4126
rect 77980 4062 77982 4114
rect 78034 4062 78036 4114
rect 77980 3892 78036 4062
rect 77980 3826 78036 3836
rect 77196 3502 77198 3554
rect 77250 3502 77252 3554
rect 77196 3490 77252 3502
rect 76188 800 76244 3332
rect 77084 3266 77140 3276
rect 78492 3164 78756 3174
rect 78548 3108 78596 3164
rect 78652 3108 78700 3164
rect 78492 3098 78756 3108
rect 3948 700 4676 756
rect 7616 0 7728 800
rect 11648 0 11760 800
rect 15680 0 15792 800
rect 19712 0 19824 800
rect 23744 0 23856 800
rect 27776 0 27888 800
rect 31808 0 31920 800
rect 35840 0 35952 800
rect 39872 0 39984 800
rect 43904 0 44016 800
rect 47936 0 48048 800
rect 51968 0 52080 800
rect 56000 0 56112 800
rect 60032 0 60144 800
rect 64064 0 64176 800
rect 68096 0 68208 800
rect 72128 0 72240 800
rect 76160 0 76272 800
<< via2 >>
rect 3388 38332 3444 38388
rect 1932 35868 1988 35924
rect 2940 35138 2996 35140
rect 2940 35086 2942 35138
rect 2942 35086 2994 35138
rect 2994 35086 2996 35138
rect 2940 35084 2996 35086
rect 10872 36874 10928 36876
rect 10872 36822 10874 36874
rect 10874 36822 10926 36874
rect 10926 36822 10928 36874
rect 10872 36820 10928 36822
rect 10976 36874 11032 36876
rect 10976 36822 10978 36874
rect 10978 36822 11030 36874
rect 11030 36822 11032 36874
rect 10976 36820 11032 36822
rect 11080 36874 11136 36876
rect 11080 36822 11082 36874
rect 11082 36822 11134 36874
rect 11134 36822 11136 36874
rect 11080 36820 11136 36822
rect 14476 37548 14532 37604
rect 7308 36370 7364 36372
rect 7308 36318 7310 36370
rect 7310 36318 7362 36370
rect 7362 36318 7364 36370
rect 7308 36316 7364 36318
rect 3948 35084 4004 35140
rect 1820 34972 1876 35028
rect 3500 35026 3556 35028
rect 3500 34974 3502 35026
rect 3502 34974 3554 35026
rect 3554 34974 3556 35026
rect 3500 34972 3556 34974
rect 1932 33404 1988 33460
rect 1932 30940 1988 30996
rect 2268 28700 2324 28756
rect 1932 28476 1988 28532
rect 1820 26684 1876 26740
rect 1932 26012 1988 26068
rect 1820 23884 1876 23940
rect 1932 23548 1988 23604
rect 3052 34300 3108 34356
rect 4284 33964 4340 34020
rect 4844 34018 4900 34020
rect 4844 33966 4846 34018
rect 4846 33966 4898 34018
rect 4898 33966 4900 34018
rect 4844 33964 4900 33966
rect 4732 33292 4788 33348
rect 4284 31778 4340 31780
rect 4284 31726 4286 31778
rect 4286 31726 4338 31778
rect 4338 31726 4340 31778
rect 4284 31724 4340 31726
rect 4060 31164 4116 31220
rect 3724 30098 3780 30100
rect 3724 30046 3726 30098
rect 3726 30046 3778 30098
rect 3778 30046 3780 30098
rect 3724 30044 3780 30046
rect 2492 29426 2548 29428
rect 2492 29374 2494 29426
rect 2494 29374 2546 29426
rect 2546 29374 2548 29426
rect 2492 29372 2548 29374
rect 2940 28642 2996 28644
rect 2940 28590 2942 28642
rect 2942 28590 2994 28642
rect 2994 28590 2996 28642
rect 2940 28588 2996 28590
rect 2380 23324 2436 23380
rect 3164 22258 3220 22260
rect 3164 22206 3166 22258
rect 3166 22206 3218 22258
rect 3218 22206 3220 22258
rect 3164 22204 3220 22206
rect 3836 22258 3892 22260
rect 3836 22206 3838 22258
rect 3838 22206 3890 22258
rect 3890 22206 3892 22258
rect 3836 22204 3892 22206
rect 9884 34972 9940 35028
rect 10872 35306 10928 35308
rect 10872 35254 10874 35306
rect 10874 35254 10926 35306
rect 10926 35254 10928 35306
rect 10872 35252 10928 35254
rect 10976 35306 11032 35308
rect 10976 35254 10978 35306
rect 10978 35254 11030 35306
rect 11030 35254 11032 35306
rect 10976 35252 11032 35254
rect 11080 35306 11136 35308
rect 11080 35254 11082 35306
rect 11082 35254 11134 35306
rect 11134 35254 11136 35306
rect 11080 35252 11136 35254
rect 10332 34076 10388 34132
rect 11004 34130 11060 34132
rect 11004 34078 11006 34130
rect 11006 34078 11058 34130
rect 11058 34078 11060 34130
rect 11004 34076 11060 34078
rect 10872 33738 10928 33740
rect 10872 33686 10874 33738
rect 10874 33686 10926 33738
rect 10926 33686 10928 33738
rect 10872 33684 10928 33686
rect 10976 33738 11032 33740
rect 10976 33686 10978 33738
rect 10978 33686 11030 33738
rect 11030 33686 11032 33738
rect 10976 33684 11032 33686
rect 11080 33738 11136 33740
rect 11080 33686 11082 33738
rect 11082 33686 11134 33738
rect 11134 33686 11136 33738
rect 11080 33684 11136 33686
rect 20860 37324 20916 37380
rect 19628 36652 19684 36708
rect 16380 36428 16436 36484
rect 17052 36482 17108 36484
rect 17052 36430 17054 36482
rect 17054 36430 17106 36482
rect 17106 36430 17108 36482
rect 17052 36428 17108 36430
rect 13804 36204 13860 36260
rect 17724 36258 17780 36260
rect 17724 36206 17726 36258
rect 17726 36206 17778 36258
rect 17778 36206 17780 36258
rect 17724 36204 17780 36206
rect 20532 36090 20588 36092
rect 20532 36038 20534 36090
rect 20534 36038 20586 36090
rect 20586 36038 20588 36090
rect 20532 36036 20588 36038
rect 20636 36090 20692 36092
rect 20636 36038 20638 36090
rect 20638 36038 20690 36090
rect 20690 36038 20692 36090
rect 20636 36036 20692 36038
rect 20740 36090 20796 36092
rect 20740 36038 20742 36090
rect 20742 36038 20794 36090
rect 20794 36038 20796 36090
rect 20740 36036 20796 36038
rect 17276 35868 17332 35924
rect 14700 35756 14756 35812
rect 13244 35586 13300 35588
rect 13244 35534 13246 35586
rect 13246 35534 13298 35586
rect 13298 35534 13300 35586
rect 13244 35532 13300 35534
rect 12236 35308 12292 35364
rect 15372 35532 15428 35588
rect 14476 34412 14532 34468
rect 16604 35420 16660 35476
rect 17052 35420 17108 35476
rect 15372 34914 15428 34916
rect 15372 34862 15374 34914
rect 15374 34862 15426 34914
rect 15426 34862 15428 34914
rect 15372 34860 15428 34862
rect 13804 34076 13860 34132
rect 11676 33516 11732 33572
rect 12572 33570 12628 33572
rect 12572 33518 12574 33570
rect 12574 33518 12626 33570
rect 12626 33518 12628 33570
rect 12572 33516 12628 33518
rect 11228 33404 11284 33460
rect 13468 33458 13524 33460
rect 13468 33406 13470 33458
rect 13470 33406 13522 33458
rect 13522 33406 13524 33458
rect 13468 33404 13524 33406
rect 13580 33234 13636 33236
rect 13580 33182 13582 33234
rect 13582 33182 13634 33234
rect 13634 33182 13636 33234
rect 13580 33180 13636 33182
rect 15932 34690 15988 34692
rect 15932 34638 15934 34690
rect 15934 34638 15986 34690
rect 15986 34638 15988 34690
rect 15932 34636 15988 34638
rect 16268 34914 16324 34916
rect 16268 34862 16270 34914
rect 16270 34862 16322 34914
rect 16322 34862 16324 34914
rect 16268 34860 16324 34862
rect 16940 34860 16996 34916
rect 15820 34412 15876 34468
rect 14476 33346 14532 33348
rect 14476 33294 14478 33346
rect 14478 33294 14530 33346
rect 14530 33294 14532 33346
rect 14476 33292 14532 33294
rect 12684 32732 12740 32788
rect 13916 32674 13972 32676
rect 13916 32622 13918 32674
rect 13918 32622 13970 32674
rect 13970 32622 13972 32674
rect 13916 32620 13972 32622
rect 10872 32170 10928 32172
rect 10872 32118 10874 32170
rect 10874 32118 10926 32170
rect 10926 32118 10928 32170
rect 10872 32116 10928 32118
rect 10976 32170 11032 32172
rect 10976 32118 10978 32170
rect 10978 32118 11030 32170
rect 11030 32118 11032 32170
rect 10976 32116 11032 32118
rect 11080 32170 11136 32172
rect 11080 32118 11082 32170
rect 11082 32118 11134 32170
rect 11134 32118 11136 32170
rect 11080 32116 11136 32118
rect 5180 31052 5236 31108
rect 9548 31388 9604 31444
rect 9996 31388 10052 31444
rect 5740 30044 5796 30100
rect 4956 29484 5012 29540
rect 4284 27916 4340 27972
rect 5292 29148 5348 29204
rect 6748 29538 6804 29540
rect 6748 29486 6750 29538
rect 6750 29486 6802 29538
rect 6802 29486 6804 29538
rect 6748 29484 6804 29486
rect 6524 29260 6580 29316
rect 6076 29202 6132 29204
rect 6076 29150 6078 29202
rect 6078 29150 6130 29202
rect 6130 29150 6132 29202
rect 6076 29148 6132 29150
rect 5628 28588 5684 28644
rect 5292 27804 5348 27860
rect 4284 25228 4340 25284
rect 6076 25340 6132 25396
rect 4844 25282 4900 25284
rect 4844 25230 4846 25282
rect 4846 25230 4898 25282
rect 4898 25230 4900 25282
rect 4844 25228 4900 25230
rect 4732 24834 4788 24836
rect 4732 24782 4734 24834
rect 4734 24782 4786 24834
rect 4786 24782 4788 24834
rect 4732 24780 4788 24782
rect 4284 24108 4340 24164
rect 4060 21756 4116 21812
rect 5516 24834 5572 24836
rect 5516 24782 5518 24834
rect 5518 24782 5570 24834
rect 5570 24782 5572 24834
rect 5516 24780 5572 24782
rect 4844 24556 4900 24612
rect 4844 24108 4900 24164
rect 5740 23938 5796 23940
rect 5740 23886 5742 23938
rect 5742 23886 5794 23938
rect 5794 23886 5796 23938
rect 5740 23884 5796 23886
rect 5740 23324 5796 23380
rect 4956 22370 5012 22372
rect 4956 22318 4958 22370
rect 4958 22318 5010 22370
rect 5010 22318 5012 22370
rect 4956 22316 5012 22318
rect 5740 22316 5796 22372
rect 4172 21644 4228 21700
rect 2716 21026 2772 21028
rect 2716 20974 2718 21026
rect 2718 20974 2770 21026
rect 2770 20974 2772 21026
rect 2716 20972 2772 20974
rect 1932 18620 1988 18676
rect 4956 21756 5012 21812
rect 4956 20860 5012 20916
rect 5740 20748 5796 20804
rect 4956 20690 5012 20692
rect 4956 20638 4958 20690
rect 4958 20638 5010 20690
rect 5010 20638 5012 20690
rect 4956 20636 5012 20638
rect 5852 20690 5908 20692
rect 5852 20638 5854 20690
rect 5854 20638 5906 20690
rect 5906 20638 5908 20690
rect 5852 20636 5908 20638
rect 4396 19740 4452 19796
rect 1932 16156 1988 16212
rect 3836 17052 3892 17108
rect 5404 19292 5460 19348
rect 5068 17778 5124 17780
rect 5068 17726 5070 17778
rect 5070 17726 5122 17778
rect 5122 17726 5124 17778
rect 5068 17724 5124 17726
rect 5292 17612 5348 17668
rect 4732 17052 4788 17108
rect 3724 16098 3780 16100
rect 3724 16046 3726 16098
rect 3726 16046 3778 16098
rect 3778 16046 3780 16098
rect 3724 16044 3780 16046
rect 4396 15986 4452 15988
rect 4396 15934 4398 15986
rect 4398 15934 4450 15986
rect 4450 15934 4452 15986
rect 4396 15932 4452 15934
rect 5292 15932 5348 15988
rect 2716 15820 2772 15876
rect 4060 15874 4116 15876
rect 4060 15822 4062 15874
rect 4062 15822 4114 15874
rect 4114 15822 4116 15874
rect 4060 15820 4116 15822
rect 1932 13692 1988 13748
rect 4844 15260 4900 15316
rect 5740 18450 5796 18452
rect 5740 18398 5742 18450
rect 5742 18398 5794 18450
rect 5794 18398 5796 18450
rect 5740 18396 5796 18398
rect 5852 17500 5908 17556
rect 5628 16156 5684 16212
rect 5740 16044 5796 16100
rect 6188 24556 6244 24612
rect 7420 29314 7476 29316
rect 7420 29262 7422 29314
rect 7422 29262 7474 29314
rect 7474 29262 7476 29314
rect 7420 29260 7476 29262
rect 6748 29148 6804 29204
rect 7084 28700 7140 28756
rect 8540 29372 8596 29428
rect 8316 28028 8372 28084
rect 9660 28082 9716 28084
rect 9660 28030 9662 28082
rect 9662 28030 9714 28082
rect 9714 28030 9716 28082
rect 9660 28028 9716 28030
rect 6748 27804 6804 27860
rect 6860 27746 6916 27748
rect 6860 27694 6862 27746
rect 6862 27694 6914 27746
rect 6914 27694 6916 27746
rect 6860 27692 6916 27694
rect 6748 27074 6804 27076
rect 6748 27022 6750 27074
rect 6750 27022 6802 27074
rect 6802 27022 6804 27074
rect 6748 27020 6804 27022
rect 6300 22204 6356 22260
rect 6188 21756 6244 21812
rect 8092 26290 8148 26292
rect 8092 26238 8094 26290
rect 8094 26238 8146 26290
rect 8146 26238 8148 26290
rect 8092 26236 8148 26238
rect 8876 26402 8932 26404
rect 8876 26350 8878 26402
rect 8878 26350 8930 26402
rect 8930 26350 8932 26402
rect 8876 26348 8932 26350
rect 10872 30602 10928 30604
rect 10872 30550 10874 30602
rect 10874 30550 10926 30602
rect 10926 30550 10928 30602
rect 10872 30548 10928 30550
rect 10976 30602 11032 30604
rect 10976 30550 10978 30602
rect 10978 30550 11030 30602
rect 11030 30550 11032 30602
rect 10976 30548 11032 30550
rect 11080 30602 11136 30604
rect 11080 30550 11082 30602
rect 11082 30550 11134 30602
rect 11134 30550 11136 30602
rect 11080 30548 11136 30550
rect 9996 29426 10052 29428
rect 9996 29374 9998 29426
rect 9998 29374 10050 29426
rect 10050 29374 10052 29426
rect 9996 29372 10052 29374
rect 10220 29260 10276 29316
rect 10220 27692 10276 27748
rect 13132 30156 13188 30212
rect 11340 29372 11396 29428
rect 10872 29034 10928 29036
rect 10872 28982 10874 29034
rect 10874 28982 10926 29034
rect 10926 28982 10928 29034
rect 10872 28980 10928 28982
rect 10976 29034 11032 29036
rect 10976 28982 10978 29034
rect 10978 28982 11030 29034
rect 11030 28982 11032 29034
rect 10976 28980 11032 28982
rect 11080 29034 11136 29036
rect 11080 28982 11082 29034
rect 11082 28982 11134 29034
rect 11134 28982 11136 29034
rect 11080 28980 11136 28982
rect 9996 27634 10052 27636
rect 9996 27582 9998 27634
rect 9998 27582 10050 27634
rect 10050 27582 10052 27634
rect 9996 27580 10052 27582
rect 9884 26684 9940 26740
rect 10108 27074 10164 27076
rect 10108 27022 10110 27074
rect 10110 27022 10162 27074
rect 10162 27022 10164 27074
rect 10108 27020 10164 27022
rect 9548 26236 9604 26292
rect 9884 26348 9940 26404
rect 8428 25116 8484 25172
rect 9660 25116 9716 25172
rect 8428 24556 8484 24612
rect 9548 24892 9604 24948
rect 8652 23378 8708 23380
rect 8652 23326 8654 23378
rect 8654 23326 8706 23378
rect 8706 23326 8708 23378
rect 8652 23324 8708 23326
rect 7196 23266 7252 23268
rect 7196 23214 7198 23266
rect 7198 23214 7250 23266
rect 7250 23214 7252 23266
rect 7196 23212 7252 23214
rect 9100 23212 9156 23268
rect 8652 22988 8708 23044
rect 6860 20690 6916 20692
rect 6860 20638 6862 20690
rect 6862 20638 6914 20690
rect 6914 20638 6916 20690
rect 6860 20636 6916 20638
rect 7308 20130 7364 20132
rect 7308 20078 7310 20130
rect 7310 20078 7362 20130
rect 7362 20078 7364 20130
rect 7308 20076 7364 20078
rect 6412 18450 6468 18452
rect 6412 18398 6414 18450
rect 6414 18398 6466 18450
rect 6466 18398 6468 18450
rect 6412 18396 6468 18398
rect 6076 17778 6132 17780
rect 6076 17726 6078 17778
rect 6078 17726 6130 17778
rect 6130 17726 6132 17778
rect 6076 17724 6132 17726
rect 6636 17554 6692 17556
rect 6636 17502 6638 17554
rect 6638 17502 6690 17554
rect 6690 17502 6692 17554
rect 6636 17500 6692 17502
rect 6188 15932 6244 15988
rect 5964 15484 6020 15540
rect 6748 17388 6804 17444
rect 5628 15314 5684 15316
rect 5628 15262 5630 15314
rect 5630 15262 5682 15314
rect 5682 15262 5684 15314
rect 5628 15260 5684 15262
rect 2716 13020 2772 13076
rect 1820 12124 1876 12180
rect 1932 11228 1988 11284
rect 1932 8818 1988 8820
rect 1932 8766 1934 8818
rect 1934 8766 1986 8818
rect 1986 8766 1988 8818
rect 1932 8764 1988 8766
rect 3612 12962 3668 12964
rect 3612 12910 3614 12962
rect 3614 12910 3666 12962
rect 3666 12910 3668 12962
rect 3612 12908 3668 12910
rect 3164 10780 3220 10836
rect 4284 11452 4340 11508
rect 4172 9826 4228 9828
rect 4172 9774 4174 9826
rect 4174 9774 4226 9826
rect 4226 9774 4228 9826
rect 4172 9772 4228 9774
rect 3164 9714 3220 9716
rect 3164 9662 3166 9714
rect 3166 9662 3218 9714
rect 3218 9662 3220 9714
rect 3164 9660 3220 9662
rect 3836 9714 3892 9716
rect 3836 9662 3838 9714
rect 3838 9662 3890 9714
rect 3890 9662 3892 9714
rect 3836 9660 3892 9662
rect 4284 9212 4340 9268
rect 2716 7644 2772 7700
rect 3836 7980 3892 8036
rect 4284 6690 4340 6692
rect 4284 6638 4286 6690
rect 4286 6638 4338 6690
rect 4338 6638 4340 6690
rect 4284 6636 4340 6638
rect 2492 6578 2548 6580
rect 2492 6526 2494 6578
rect 2494 6526 2546 6578
rect 2546 6526 2548 6578
rect 2492 6524 2548 6526
rect 5068 14252 5124 14308
rect 4844 13916 4900 13972
rect 4732 10834 4788 10836
rect 4732 10782 4734 10834
rect 4734 10782 4786 10834
rect 4786 10782 4788 10834
rect 4732 10780 4788 10782
rect 4620 10332 4676 10388
rect 4732 9884 4788 9940
rect 4620 9772 4676 9828
rect 7196 15036 7252 15092
rect 8540 20076 8596 20132
rect 8092 20018 8148 20020
rect 8092 19966 8094 20018
rect 8094 19966 8146 20018
rect 8146 19966 8148 20018
rect 8092 19964 8148 19966
rect 7532 18396 7588 18452
rect 7980 17388 8036 17444
rect 7532 15932 7588 15988
rect 6076 14252 6132 14308
rect 5740 12908 5796 12964
rect 5516 12178 5572 12180
rect 5516 12126 5518 12178
rect 5518 12126 5570 12178
rect 5570 12126 5572 12178
rect 5516 12124 5572 12126
rect 5068 11506 5124 11508
rect 5068 11454 5070 11506
rect 5070 11454 5122 11506
rect 5122 11454 5124 11506
rect 5068 11452 5124 11454
rect 6972 11506 7028 11508
rect 6972 11454 6974 11506
rect 6974 11454 7026 11506
rect 7026 11454 7028 11506
rect 6972 11452 7028 11454
rect 6188 10780 6244 10836
rect 5180 10668 5236 10724
rect 5068 10386 5124 10388
rect 5068 10334 5070 10386
rect 5070 10334 5122 10386
rect 5122 10334 5124 10386
rect 5068 10332 5124 10334
rect 5068 9996 5124 10052
rect 5852 10722 5908 10724
rect 5852 10670 5854 10722
rect 5854 10670 5906 10722
rect 5906 10670 5908 10722
rect 5852 10668 5908 10670
rect 5628 10610 5684 10612
rect 5628 10558 5630 10610
rect 5630 10558 5682 10610
rect 5682 10558 5684 10610
rect 5628 10556 5684 10558
rect 7644 15538 7700 15540
rect 7644 15486 7646 15538
rect 7646 15486 7698 15538
rect 7698 15486 7700 15538
rect 7644 15484 7700 15486
rect 6972 10556 7028 10612
rect 6412 9996 6468 10052
rect 6636 10444 6692 10500
rect 6188 9938 6244 9940
rect 6188 9886 6190 9938
rect 6190 9886 6242 9938
rect 6242 9886 6244 9938
rect 6188 9884 6244 9886
rect 5740 9826 5796 9828
rect 5740 9774 5742 9826
rect 5742 9774 5794 9826
rect 5794 9774 5796 9826
rect 5740 9772 5796 9774
rect 4844 6690 4900 6692
rect 4844 6638 4846 6690
rect 4846 6638 4898 6690
rect 4898 6638 4900 6690
rect 4844 6636 4900 6638
rect 4396 4956 4452 5012
rect 1932 4114 1988 4116
rect 1932 4062 1934 4114
rect 1934 4062 1986 4114
rect 1986 4062 1988 4114
rect 1932 4060 1988 4062
rect 4284 3724 4340 3780
rect 4284 3554 4340 3556
rect 4284 3502 4286 3554
rect 4286 3502 4338 3554
rect 4338 3502 4340 3554
rect 4284 3500 4340 3502
rect 1932 1484 1988 1540
rect 5292 9212 5348 9268
rect 5516 9154 5572 9156
rect 5516 9102 5518 9154
rect 5518 9102 5570 9154
rect 5570 9102 5572 9154
rect 5516 9100 5572 9102
rect 5628 8034 5684 8036
rect 5628 7982 5630 8034
rect 5630 7982 5682 8034
rect 5682 7982 5684 8034
rect 5628 7980 5684 7982
rect 7868 13020 7924 13076
rect 6076 7308 6132 7364
rect 5180 3724 5236 3780
rect 5740 4060 5796 4116
rect 5740 3500 5796 3556
rect 7756 11116 7812 11172
rect 7532 10668 7588 10724
rect 7084 9100 7140 9156
rect 8540 16098 8596 16100
rect 8540 16046 8542 16098
rect 8542 16046 8594 16098
rect 8594 16046 8596 16098
rect 8540 16044 8596 16046
rect 8092 15036 8148 15092
rect 9436 21532 9492 21588
rect 8988 21474 9044 21476
rect 8988 21422 8990 21474
rect 8990 21422 9042 21474
rect 9042 21422 9044 21474
rect 8988 21420 9044 21422
rect 10668 28700 10724 28756
rect 11788 29314 11844 29316
rect 11788 29262 11790 29314
rect 11790 29262 11842 29314
rect 11842 29262 11844 29314
rect 11788 29260 11844 29262
rect 13244 29202 13300 29204
rect 13244 29150 13246 29202
rect 13246 29150 13298 29202
rect 13298 29150 13300 29202
rect 13244 29148 13300 29150
rect 13804 30044 13860 30100
rect 11340 28588 11396 28644
rect 11004 27692 11060 27748
rect 10872 27466 10928 27468
rect 10872 27414 10874 27466
rect 10874 27414 10926 27466
rect 10926 27414 10928 27466
rect 10872 27412 10928 27414
rect 10976 27466 11032 27468
rect 10976 27414 10978 27466
rect 10978 27414 11030 27466
rect 11030 27414 11032 27466
rect 10976 27412 11032 27414
rect 11080 27466 11136 27468
rect 11080 27414 11082 27466
rect 11082 27414 11134 27466
rect 11134 27414 11136 27466
rect 11080 27412 11136 27414
rect 11228 26684 11284 26740
rect 10556 26348 10612 26404
rect 10872 25898 10928 25900
rect 10872 25846 10874 25898
rect 10874 25846 10926 25898
rect 10926 25846 10928 25898
rect 10872 25844 10928 25846
rect 10976 25898 11032 25900
rect 10976 25846 10978 25898
rect 10978 25846 11030 25898
rect 11030 25846 11032 25898
rect 10976 25844 11032 25846
rect 11080 25898 11136 25900
rect 11080 25846 11082 25898
rect 11082 25846 11134 25898
rect 11134 25846 11136 25898
rect 11080 25844 11136 25846
rect 11564 26236 11620 26292
rect 10220 24892 10276 24948
rect 9660 23324 9716 23380
rect 10220 22876 10276 22932
rect 9996 21644 10052 21700
rect 9884 21532 9940 21588
rect 9996 20802 10052 20804
rect 9996 20750 9998 20802
rect 9998 20750 10050 20802
rect 10050 20750 10052 20802
rect 9996 20748 10052 20750
rect 10108 20578 10164 20580
rect 10108 20526 10110 20578
rect 10110 20526 10162 20578
rect 10162 20526 10164 20578
rect 10108 20524 10164 20526
rect 9660 20018 9716 20020
rect 9660 19966 9662 20018
rect 9662 19966 9714 20018
rect 9714 19966 9716 20018
rect 9660 19964 9716 19966
rect 10108 20018 10164 20020
rect 10108 19966 10110 20018
rect 10110 19966 10162 20018
rect 10162 19966 10164 20018
rect 10108 19964 10164 19966
rect 10108 19068 10164 19124
rect 8988 16770 9044 16772
rect 8988 16718 8990 16770
rect 8990 16718 9042 16770
rect 9042 16718 9044 16770
rect 8988 16716 9044 16718
rect 9324 16044 9380 16100
rect 8652 13916 8708 13972
rect 8652 13692 8708 13748
rect 8316 11506 8372 11508
rect 8316 11454 8318 11506
rect 8318 11454 8370 11506
rect 8370 11454 8372 11506
rect 8316 11452 8372 11454
rect 8764 11170 8820 11172
rect 8764 11118 8766 11170
rect 8766 11118 8818 11170
rect 8818 11118 8820 11170
rect 8764 11116 8820 11118
rect 7980 10668 8036 10724
rect 9548 10722 9604 10724
rect 9548 10670 9550 10722
rect 9550 10670 9602 10722
rect 9602 10670 9604 10722
rect 9548 10668 9604 10670
rect 7868 9436 7924 9492
rect 7420 8764 7476 8820
rect 8428 9154 8484 9156
rect 8428 9102 8430 9154
rect 8430 9102 8482 9154
rect 8482 9102 8484 9154
rect 8428 9100 8484 9102
rect 7420 7362 7476 7364
rect 7420 7310 7422 7362
rect 7422 7310 7474 7362
rect 7474 7310 7476 7362
rect 7420 7308 7476 7310
rect 8876 7532 8932 7588
rect 8652 7308 8708 7364
rect 10108 15932 10164 15988
rect 9996 14700 10052 14756
rect 10872 24330 10928 24332
rect 10872 24278 10874 24330
rect 10874 24278 10926 24330
rect 10926 24278 10928 24330
rect 10872 24276 10928 24278
rect 10976 24330 11032 24332
rect 10976 24278 10978 24330
rect 10978 24278 11030 24330
rect 11030 24278 11032 24330
rect 10976 24276 11032 24278
rect 11080 24330 11136 24332
rect 11080 24278 11082 24330
rect 11082 24278 11134 24330
rect 11134 24278 11136 24330
rect 11080 24276 11136 24278
rect 10872 22762 10928 22764
rect 10872 22710 10874 22762
rect 10874 22710 10926 22762
rect 10926 22710 10928 22762
rect 10872 22708 10928 22710
rect 10976 22762 11032 22764
rect 10976 22710 10978 22762
rect 10978 22710 11030 22762
rect 11030 22710 11032 22762
rect 10976 22708 11032 22710
rect 11080 22762 11136 22764
rect 11080 22710 11082 22762
rect 11082 22710 11134 22762
rect 11134 22710 11136 22762
rect 11080 22708 11136 22710
rect 10556 21756 10612 21812
rect 11340 22092 11396 22148
rect 10444 21644 10500 21700
rect 10332 21586 10388 21588
rect 10332 21534 10334 21586
rect 10334 21534 10386 21586
rect 10386 21534 10388 21586
rect 10332 21532 10388 21534
rect 10556 21308 10612 21364
rect 10444 20802 10500 20804
rect 10444 20750 10446 20802
rect 10446 20750 10498 20802
rect 10498 20750 10500 20802
rect 10444 20748 10500 20750
rect 11116 21586 11172 21588
rect 11116 21534 11118 21586
rect 11118 21534 11170 21586
rect 11170 21534 11172 21586
rect 11116 21532 11172 21534
rect 13804 27804 13860 27860
rect 12124 27580 12180 27636
rect 11788 26684 11844 26740
rect 11676 24444 11732 24500
rect 12012 25730 12068 25732
rect 12012 25678 12014 25730
rect 12014 25678 12066 25730
rect 12066 25678 12068 25730
rect 12012 25676 12068 25678
rect 11788 21756 11844 21812
rect 11564 21644 11620 21700
rect 10872 21194 10928 21196
rect 10872 21142 10874 21194
rect 10874 21142 10926 21194
rect 10926 21142 10928 21194
rect 10872 21140 10928 21142
rect 10976 21194 11032 21196
rect 10976 21142 10978 21194
rect 10978 21142 11030 21194
rect 11030 21142 11032 21194
rect 10976 21140 11032 21142
rect 11080 21194 11136 21196
rect 11080 21142 11082 21194
rect 11082 21142 11134 21194
rect 11134 21142 11136 21194
rect 11080 21140 11136 21142
rect 10332 20188 10388 20244
rect 10668 20188 10724 20244
rect 10780 20412 10836 20468
rect 11004 20748 11060 20804
rect 11452 21474 11508 21476
rect 11452 21422 11454 21474
rect 11454 21422 11506 21474
rect 11506 21422 11508 21474
rect 11452 21420 11508 21422
rect 11900 21308 11956 21364
rect 12012 21532 12068 21588
rect 11676 20914 11732 20916
rect 11676 20862 11678 20914
rect 11678 20862 11730 20914
rect 11730 20862 11732 20914
rect 11676 20860 11732 20862
rect 11228 20636 11284 20692
rect 10556 19404 10612 19460
rect 10872 19626 10928 19628
rect 10872 19574 10874 19626
rect 10874 19574 10926 19626
rect 10926 19574 10928 19626
rect 10872 19572 10928 19574
rect 10976 19626 11032 19628
rect 10976 19574 10978 19626
rect 10978 19574 11030 19626
rect 11030 19574 11032 19626
rect 10976 19572 11032 19574
rect 11080 19626 11136 19628
rect 11080 19574 11082 19626
rect 11082 19574 11134 19626
rect 11134 19574 11136 19626
rect 11080 19572 11136 19574
rect 10892 19122 10948 19124
rect 10892 19070 10894 19122
rect 10894 19070 10946 19122
rect 10946 19070 10948 19122
rect 10892 19068 10948 19070
rect 11340 19122 11396 19124
rect 11340 19070 11342 19122
rect 11342 19070 11394 19122
rect 11394 19070 11396 19122
rect 11340 19068 11396 19070
rect 11228 18844 11284 18900
rect 10872 18058 10928 18060
rect 10872 18006 10874 18058
rect 10874 18006 10926 18058
rect 10926 18006 10928 18058
rect 10872 18004 10928 18006
rect 10976 18058 11032 18060
rect 10976 18006 10978 18058
rect 10978 18006 11030 18058
rect 11030 18006 11032 18058
rect 10976 18004 11032 18006
rect 11080 18058 11136 18060
rect 11080 18006 11082 18058
rect 11082 18006 11134 18058
rect 11134 18006 11136 18058
rect 11080 18004 11136 18006
rect 11788 20636 11844 20692
rect 11676 20578 11732 20580
rect 11676 20526 11678 20578
rect 11678 20526 11730 20578
rect 11730 20526 11732 20578
rect 11676 20524 11732 20526
rect 11676 20018 11732 20020
rect 11676 19966 11678 20018
rect 11678 19966 11730 20018
rect 11730 19966 11732 20018
rect 11676 19964 11732 19966
rect 11900 20076 11956 20132
rect 11788 17724 11844 17780
rect 11676 17554 11732 17556
rect 11676 17502 11678 17554
rect 11678 17502 11730 17554
rect 11730 17502 11732 17554
rect 11676 17500 11732 17502
rect 11676 17106 11732 17108
rect 11676 17054 11678 17106
rect 11678 17054 11730 17106
rect 11730 17054 11732 17106
rect 11676 17052 11732 17054
rect 10892 16604 10948 16660
rect 11340 16882 11396 16884
rect 11340 16830 11342 16882
rect 11342 16830 11394 16882
rect 11394 16830 11396 16882
rect 11340 16828 11396 16830
rect 12908 25676 12964 25732
rect 12796 25506 12852 25508
rect 12796 25454 12798 25506
rect 12798 25454 12850 25506
rect 12850 25454 12852 25506
rect 12796 25452 12852 25454
rect 13580 25452 13636 25508
rect 12572 25394 12628 25396
rect 12572 25342 12574 25394
rect 12574 25342 12626 25394
rect 12626 25342 12628 25394
rect 12572 25340 12628 25342
rect 13468 24610 13524 24612
rect 13468 24558 13470 24610
rect 13470 24558 13522 24610
rect 13522 24558 13524 24610
rect 13468 24556 13524 24558
rect 13580 22876 13636 22932
rect 14252 32786 14308 32788
rect 14252 32734 14254 32786
rect 14254 32734 14306 32786
rect 14306 32734 14308 32786
rect 14252 32732 14308 32734
rect 14588 32732 14644 32788
rect 14588 32562 14644 32564
rect 14588 32510 14590 32562
rect 14590 32510 14642 32562
rect 14642 32510 14644 32562
rect 14588 32508 14644 32510
rect 14140 31724 14196 31780
rect 14924 32844 14980 32900
rect 15708 33068 15764 33124
rect 18284 35420 18340 35476
rect 18956 35420 19012 35476
rect 18060 34914 18116 34916
rect 18060 34862 18062 34914
rect 18062 34862 18114 34914
rect 18114 34862 18116 34914
rect 18060 34860 18116 34862
rect 17500 34636 17556 34692
rect 17612 34188 17668 34244
rect 18284 34188 18340 34244
rect 16044 34076 16100 34132
rect 15148 32562 15204 32564
rect 15148 32510 15150 32562
rect 15150 32510 15202 32562
rect 15202 32510 15204 32562
rect 15148 32508 15204 32510
rect 17836 34130 17892 34132
rect 17836 34078 17838 34130
rect 17838 34078 17890 34130
rect 17890 34078 17892 34130
rect 17836 34076 17892 34078
rect 18172 33964 18228 34020
rect 15372 32396 15428 32452
rect 15036 31724 15092 31780
rect 14812 31500 14868 31556
rect 14924 30882 14980 30884
rect 14924 30830 14926 30882
rect 14926 30830 14978 30882
rect 14978 30830 14980 30882
rect 14924 30828 14980 30830
rect 14476 30604 14532 30660
rect 14700 30210 14756 30212
rect 14700 30158 14702 30210
rect 14702 30158 14754 30210
rect 14754 30158 14756 30210
rect 14700 30156 14756 30158
rect 14364 30044 14420 30100
rect 14700 28754 14756 28756
rect 14700 28702 14702 28754
rect 14702 28702 14754 28754
rect 14754 28702 14756 28754
rect 14700 28700 14756 28702
rect 14252 28028 14308 28084
rect 14252 24556 14308 24612
rect 13916 24498 13972 24500
rect 13916 24446 13918 24498
rect 13918 24446 13970 24498
rect 13970 24446 13972 24498
rect 13916 24444 13972 24446
rect 12684 21810 12740 21812
rect 12684 21758 12686 21810
rect 12686 21758 12738 21810
rect 12738 21758 12740 21810
rect 12684 21756 12740 21758
rect 12124 21084 12180 21140
rect 13468 22146 13524 22148
rect 13468 22094 13470 22146
rect 13470 22094 13522 22146
rect 13522 22094 13524 22146
rect 13468 22092 13524 22094
rect 13804 22146 13860 22148
rect 13804 22094 13806 22146
rect 13806 22094 13858 22146
rect 13858 22094 13860 22146
rect 13804 22092 13860 22094
rect 13468 21810 13524 21812
rect 13468 21758 13470 21810
rect 13470 21758 13522 21810
rect 13522 21758 13524 21810
rect 13468 21756 13524 21758
rect 12236 20412 12292 20468
rect 12572 20188 12628 20244
rect 12124 19234 12180 19236
rect 12124 19182 12126 19234
rect 12126 19182 12178 19234
rect 12178 19182 12180 19234
rect 12124 19180 12180 19182
rect 12684 19180 12740 19236
rect 12348 18396 12404 18452
rect 13020 18620 13076 18676
rect 13132 18450 13188 18452
rect 13132 18398 13134 18450
rect 13134 18398 13186 18450
rect 13186 18398 13188 18450
rect 13132 18396 13188 18398
rect 12908 17836 12964 17892
rect 12572 17778 12628 17780
rect 12572 17726 12574 17778
rect 12574 17726 12626 17778
rect 12626 17726 12628 17778
rect 12572 17724 12628 17726
rect 11228 16716 11284 16772
rect 12348 16770 12404 16772
rect 12348 16718 12350 16770
rect 12350 16718 12402 16770
rect 12402 16718 12404 16770
rect 12348 16716 12404 16718
rect 10872 16490 10928 16492
rect 10872 16438 10874 16490
rect 10874 16438 10926 16490
rect 10926 16438 10928 16490
rect 10872 16436 10928 16438
rect 10976 16490 11032 16492
rect 10976 16438 10978 16490
rect 10978 16438 11030 16490
rect 11030 16438 11032 16490
rect 10976 16436 11032 16438
rect 11080 16490 11136 16492
rect 11080 16438 11082 16490
rect 11082 16438 11134 16490
rect 11134 16438 11136 16490
rect 11228 16492 11284 16548
rect 11080 16436 11136 16438
rect 10556 16268 10612 16324
rect 11564 16380 11620 16436
rect 10332 16210 10388 16212
rect 10332 16158 10334 16210
rect 10334 16158 10386 16210
rect 10386 16158 10388 16210
rect 10332 16156 10388 16158
rect 11116 16156 11172 16212
rect 11340 15986 11396 15988
rect 11340 15934 11342 15986
rect 11342 15934 11394 15986
rect 11394 15934 11396 15986
rect 11340 15932 11396 15934
rect 11900 16268 11956 16324
rect 10444 15260 10500 15316
rect 11564 15314 11620 15316
rect 11564 15262 11566 15314
rect 11566 15262 11618 15314
rect 11618 15262 11620 15314
rect 11564 15260 11620 15262
rect 10556 15036 10612 15092
rect 10872 14922 10928 14924
rect 10872 14870 10874 14922
rect 10874 14870 10926 14922
rect 10926 14870 10928 14922
rect 10872 14868 10928 14870
rect 10976 14922 11032 14924
rect 10976 14870 10978 14922
rect 10978 14870 11030 14922
rect 11030 14870 11032 14922
rect 10976 14868 11032 14870
rect 11080 14922 11136 14924
rect 11080 14870 11082 14922
rect 11082 14870 11134 14922
rect 11134 14870 11136 14922
rect 11080 14868 11136 14870
rect 10556 13916 10612 13972
rect 11452 13916 11508 13972
rect 10108 10444 10164 10500
rect 10444 11116 10500 11172
rect 10220 9324 10276 9380
rect 9996 8818 10052 8820
rect 9996 8766 9998 8818
rect 9998 8766 10050 8818
rect 10050 8766 10052 8818
rect 9996 8764 10052 8766
rect 9660 7532 9716 7588
rect 9212 6860 9268 6916
rect 9772 6748 9828 6804
rect 8988 6076 9044 6132
rect 10556 10498 10612 10500
rect 10556 10446 10558 10498
rect 10558 10446 10610 10498
rect 10610 10446 10612 10498
rect 10556 10444 10612 10446
rect 12012 15148 12068 15204
rect 12124 16604 12180 16660
rect 11452 13468 11508 13524
rect 10872 13354 10928 13356
rect 10872 13302 10874 13354
rect 10874 13302 10926 13354
rect 10926 13302 10928 13354
rect 10872 13300 10928 13302
rect 10976 13354 11032 13356
rect 10976 13302 10978 13354
rect 10978 13302 11030 13354
rect 11030 13302 11032 13354
rect 10976 13300 11032 13302
rect 11080 13354 11136 13356
rect 11080 13302 11082 13354
rect 11082 13302 11134 13354
rect 11134 13302 11136 13354
rect 11080 13300 11136 13302
rect 12460 16156 12516 16212
rect 12684 17500 12740 17556
rect 12684 16940 12740 16996
rect 12236 15260 12292 15316
rect 12348 15932 12404 15988
rect 12908 16156 12964 16212
rect 13020 16828 13076 16884
rect 12348 14028 12404 14084
rect 10872 11786 10928 11788
rect 10872 11734 10874 11786
rect 10874 11734 10926 11786
rect 10926 11734 10928 11786
rect 10872 11732 10928 11734
rect 10976 11786 11032 11788
rect 10976 11734 10978 11786
rect 10978 11734 11030 11786
rect 11030 11734 11032 11786
rect 10976 11732 11032 11734
rect 11080 11786 11136 11788
rect 11080 11734 11082 11786
rect 11082 11734 11134 11786
rect 11134 11734 11136 11786
rect 11080 11732 11136 11734
rect 12348 12796 12404 12852
rect 12012 12124 12068 12180
rect 13132 15314 13188 15316
rect 13132 15262 13134 15314
rect 13134 15262 13186 15314
rect 13186 15262 13188 15314
rect 13132 15260 13188 15262
rect 13580 21196 13636 21252
rect 13468 17724 13524 17780
rect 13580 17836 13636 17892
rect 13580 16268 13636 16324
rect 14252 22146 14308 22148
rect 14252 22094 14254 22146
rect 14254 22094 14306 22146
rect 14306 22094 14308 22146
rect 14252 22092 14308 22094
rect 13916 19740 13972 19796
rect 14028 21868 14084 21924
rect 13356 14812 13412 14868
rect 13804 17948 13860 18004
rect 13020 13970 13076 13972
rect 13020 13918 13022 13970
rect 13022 13918 13074 13970
rect 13074 13918 13076 13970
rect 13020 13916 13076 13918
rect 13244 13804 13300 13860
rect 12684 12178 12740 12180
rect 12684 12126 12686 12178
rect 12686 12126 12738 12178
rect 12738 12126 12740 12178
rect 12684 12124 12740 12126
rect 11788 11170 11844 11172
rect 11788 11118 11790 11170
rect 11790 11118 11842 11170
rect 11842 11118 11844 11170
rect 11788 11116 11844 11118
rect 11228 10668 11284 10724
rect 11340 10444 11396 10500
rect 10872 10218 10928 10220
rect 10872 10166 10874 10218
rect 10874 10166 10926 10218
rect 10926 10166 10928 10218
rect 10872 10164 10928 10166
rect 10976 10218 11032 10220
rect 10976 10166 10978 10218
rect 10978 10166 11030 10218
rect 11030 10166 11032 10218
rect 10976 10164 11032 10166
rect 11080 10218 11136 10220
rect 11080 10166 11082 10218
rect 11082 10166 11134 10218
rect 11134 10166 11136 10218
rect 11080 10164 11136 10166
rect 10668 9100 10724 9156
rect 10780 9436 10836 9492
rect 11676 10108 11732 10164
rect 11788 10556 11844 10612
rect 11788 9772 11844 9828
rect 11452 9154 11508 9156
rect 11452 9102 11454 9154
rect 11454 9102 11506 9154
rect 11506 9102 11508 9154
rect 11452 9100 11508 9102
rect 10872 8650 10928 8652
rect 10872 8598 10874 8650
rect 10874 8598 10926 8650
rect 10926 8598 10928 8650
rect 10872 8596 10928 8598
rect 10976 8650 11032 8652
rect 10976 8598 10978 8650
rect 10978 8598 11030 8650
rect 11030 8598 11032 8650
rect 10976 8596 11032 8598
rect 11080 8650 11136 8652
rect 11080 8598 11082 8650
rect 11082 8598 11134 8650
rect 11134 8598 11136 8650
rect 11080 8596 11136 8598
rect 10444 8204 10500 8260
rect 11340 7644 11396 7700
rect 11116 7586 11172 7588
rect 11116 7534 11118 7586
rect 11118 7534 11170 7586
rect 11170 7534 11172 7586
rect 11116 7532 11172 7534
rect 10872 7082 10928 7084
rect 10872 7030 10874 7082
rect 10874 7030 10926 7082
rect 10926 7030 10928 7082
rect 10872 7028 10928 7030
rect 10976 7082 11032 7084
rect 10976 7030 10978 7082
rect 10978 7030 11030 7082
rect 11030 7030 11032 7082
rect 10976 7028 11032 7030
rect 11080 7082 11136 7084
rect 11080 7030 11082 7082
rect 11082 7030 11134 7082
rect 11134 7030 11136 7082
rect 11080 7028 11136 7030
rect 9996 6076 10052 6132
rect 8988 5628 9044 5684
rect 11116 6018 11172 6020
rect 11116 5966 11118 6018
rect 11118 5966 11170 6018
rect 11170 5966 11172 6018
rect 11116 5964 11172 5966
rect 10872 5514 10928 5516
rect 10872 5462 10874 5514
rect 10874 5462 10926 5514
rect 10926 5462 10928 5514
rect 10872 5460 10928 5462
rect 10976 5514 11032 5516
rect 10976 5462 10978 5514
rect 10978 5462 11030 5514
rect 11030 5462 11032 5514
rect 10976 5460 11032 5462
rect 11080 5514 11136 5516
rect 11080 5462 11082 5514
rect 11082 5462 11134 5514
rect 11134 5462 11136 5514
rect 11080 5460 11136 5462
rect 9212 4898 9268 4900
rect 9212 4846 9214 4898
rect 9214 4846 9266 4898
rect 9266 4846 9268 4898
rect 9212 4844 9268 4846
rect 10780 5010 10836 5012
rect 10780 4958 10782 5010
rect 10782 4958 10834 5010
rect 10834 4958 10836 5010
rect 10780 4956 10836 4958
rect 10332 4844 10388 4900
rect 10872 3946 10928 3948
rect 10872 3894 10874 3946
rect 10874 3894 10926 3946
rect 10926 3894 10928 3946
rect 10872 3892 10928 3894
rect 10976 3946 11032 3948
rect 10976 3894 10978 3946
rect 10978 3894 11030 3946
rect 11030 3894 11032 3946
rect 10976 3892 11032 3894
rect 11080 3946 11136 3948
rect 11080 3894 11082 3946
rect 11082 3894 11134 3946
rect 11134 3894 11136 3946
rect 11080 3892 11136 3894
rect 6972 2380 7028 2436
rect 8204 3442 8260 3444
rect 8204 3390 8206 3442
rect 8206 3390 8258 3442
rect 8258 3390 8260 3442
rect 8204 3388 8260 3390
rect 11788 7532 11844 7588
rect 11564 5682 11620 5684
rect 11564 5630 11566 5682
rect 11566 5630 11618 5682
rect 11618 5630 11620 5682
rect 11564 5628 11620 5630
rect 12124 11340 12180 11396
rect 12012 10668 12068 10724
rect 12684 11788 12740 11844
rect 12012 10108 12068 10164
rect 12348 9324 12404 9380
rect 12460 8540 12516 8596
rect 13020 12796 13076 12852
rect 12908 12012 12964 12068
rect 13020 11788 13076 11844
rect 12796 11340 12852 11396
rect 12796 10556 12852 10612
rect 12908 10444 12964 10500
rect 12124 7644 12180 7700
rect 12572 8428 12628 8484
rect 12012 7308 12068 7364
rect 12460 4732 12516 4788
rect 12796 9100 12852 9156
rect 12684 5906 12740 5908
rect 12684 5854 12686 5906
rect 12686 5854 12738 5906
rect 12738 5854 12740 5906
rect 12684 5852 12740 5854
rect 13692 14028 13748 14084
rect 14140 21810 14196 21812
rect 14140 21758 14142 21810
rect 14142 21758 14194 21810
rect 14194 21758 14196 21810
rect 14140 21756 14196 21758
rect 14364 21308 14420 21364
rect 14588 25452 14644 25508
rect 15036 30044 15092 30100
rect 14924 28700 14980 28756
rect 14924 28028 14980 28084
rect 15932 32450 15988 32452
rect 15932 32398 15934 32450
rect 15934 32398 15986 32450
rect 15986 32398 15988 32450
rect 15932 32396 15988 32398
rect 16716 33122 16772 33124
rect 16716 33070 16718 33122
rect 16718 33070 16770 33122
rect 16770 33070 16772 33122
rect 16716 33068 16772 33070
rect 16268 32732 16324 32788
rect 16380 32956 16436 33012
rect 16380 32396 16436 32452
rect 16716 32284 16772 32340
rect 15260 30716 15316 30772
rect 15596 30210 15652 30212
rect 15596 30158 15598 30210
rect 15598 30158 15650 30210
rect 15650 30158 15652 30210
rect 15596 30156 15652 30158
rect 15484 30044 15540 30100
rect 15484 29596 15540 29652
rect 20532 34522 20588 34524
rect 20532 34470 20534 34522
rect 20534 34470 20586 34522
rect 20586 34470 20588 34522
rect 20532 34468 20588 34470
rect 20636 34522 20692 34524
rect 20636 34470 20638 34522
rect 20638 34470 20690 34522
rect 20690 34470 20692 34522
rect 20636 34468 20692 34470
rect 20740 34522 20796 34524
rect 20740 34470 20742 34522
rect 20742 34470 20794 34522
rect 20794 34470 20796 34522
rect 20740 34468 20796 34470
rect 18508 33292 18564 33348
rect 18732 33964 18788 34020
rect 18620 33234 18676 33236
rect 18620 33182 18622 33234
rect 18622 33182 18674 33234
rect 18674 33182 18676 33234
rect 18620 33180 18676 33182
rect 20524 34130 20580 34132
rect 20524 34078 20526 34130
rect 20526 34078 20578 34130
rect 20578 34078 20580 34130
rect 20524 34076 20580 34078
rect 19516 34018 19572 34020
rect 19516 33966 19518 34018
rect 19518 33966 19570 34018
rect 19570 33966 19572 34018
rect 19516 33964 19572 33966
rect 21644 37436 21700 37492
rect 21532 35084 21588 35140
rect 21420 34076 21476 34132
rect 19740 33516 19796 33572
rect 16044 31554 16100 31556
rect 16044 31502 16046 31554
rect 16046 31502 16098 31554
rect 16098 31502 16100 31554
rect 16044 31500 16100 31502
rect 17836 31666 17892 31668
rect 17836 31614 17838 31666
rect 17838 31614 17890 31666
rect 17890 31614 17892 31666
rect 17836 31612 17892 31614
rect 18508 31836 18564 31892
rect 18396 31276 18452 31332
rect 18956 31836 19012 31892
rect 16492 30434 16548 30436
rect 16492 30382 16494 30434
rect 16494 30382 16546 30434
rect 16546 30382 16548 30434
rect 16492 30380 16548 30382
rect 16156 30268 16212 30324
rect 17948 30940 18004 30996
rect 16380 30098 16436 30100
rect 16380 30046 16382 30098
rect 16382 30046 16434 30098
rect 16434 30046 16436 30098
rect 16380 30044 16436 30046
rect 15932 29932 15988 29988
rect 16268 29650 16324 29652
rect 16268 29598 16270 29650
rect 16270 29598 16322 29650
rect 16322 29598 16324 29650
rect 16268 29596 16324 29598
rect 15708 29148 15764 29204
rect 15596 28364 15652 28420
rect 14812 25116 14868 25172
rect 14812 24892 14868 24948
rect 14812 24220 14868 24276
rect 15596 27746 15652 27748
rect 15596 27694 15598 27746
rect 15598 27694 15650 27746
rect 15650 27694 15652 27746
rect 15596 27692 15652 27694
rect 16156 29036 16212 29092
rect 16268 27746 16324 27748
rect 16268 27694 16270 27746
rect 16270 27694 16322 27746
rect 16322 27694 16324 27746
rect 16268 27692 16324 27694
rect 15484 25618 15540 25620
rect 15484 25566 15486 25618
rect 15486 25566 15538 25618
rect 15538 25566 15540 25618
rect 15484 25564 15540 25566
rect 15820 25564 15876 25620
rect 15708 25452 15764 25508
rect 15484 25116 15540 25172
rect 15820 24892 15876 24948
rect 15484 24556 15540 24612
rect 15484 24220 15540 24276
rect 15036 23042 15092 23044
rect 15036 22990 15038 23042
rect 15038 22990 15090 23042
rect 15090 22990 15092 23042
rect 15036 22988 15092 22990
rect 14476 21810 14532 21812
rect 14476 21758 14478 21810
rect 14478 21758 14530 21810
rect 14530 21758 14532 21810
rect 14476 21756 14532 21758
rect 14476 21196 14532 21252
rect 14924 21980 14980 22036
rect 14364 19010 14420 19012
rect 14364 18958 14366 19010
rect 14366 18958 14418 19010
rect 14418 18958 14420 19010
rect 14364 18956 14420 18958
rect 14252 18620 14308 18676
rect 14812 19404 14868 19460
rect 14812 19122 14868 19124
rect 14812 19070 14814 19122
rect 14814 19070 14866 19122
rect 14866 19070 14868 19122
rect 14812 19068 14868 19070
rect 14700 18508 14756 18564
rect 14588 18284 14644 18340
rect 14252 17724 14308 17780
rect 14700 17778 14756 17780
rect 14700 17726 14702 17778
rect 14702 17726 14754 17778
rect 14754 17726 14756 17778
rect 14700 17724 14756 17726
rect 14028 17164 14084 17220
rect 13916 15260 13972 15316
rect 13916 13858 13972 13860
rect 13916 13806 13918 13858
rect 13918 13806 13970 13858
rect 13970 13806 13972 13858
rect 13916 13804 13972 13806
rect 14364 16044 14420 16100
rect 15372 23548 15428 23604
rect 15820 23548 15876 23604
rect 16156 23884 16212 23940
rect 16268 23378 16324 23380
rect 16268 23326 16270 23378
rect 16270 23326 16322 23378
rect 16322 23326 16324 23378
rect 16268 23324 16324 23326
rect 15372 23154 15428 23156
rect 15372 23102 15374 23154
rect 15374 23102 15426 23154
rect 15426 23102 15428 23154
rect 15372 23100 15428 23102
rect 15484 22988 15540 23044
rect 15484 21868 15540 21924
rect 15596 21698 15652 21700
rect 15596 21646 15598 21698
rect 15598 21646 15650 21698
rect 15650 21646 15652 21698
rect 15596 21644 15652 21646
rect 15036 19404 15092 19460
rect 15708 20524 15764 20580
rect 16044 23266 16100 23268
rect 16044 23214 16046 23266
rect 16046 23214 16098 23266
rect 16098 23214 16100 23266
rect 16044 23212 16100 23214
rect 15932 23154 15988 23156
rect 15932 23102 15934 23154
rect 15934 23102 15986 23154
rect 15986 23102 15988 23154
rect 15932 23100 15988 23102
rect 15932 22316 15988 22372
rect 16268 22258 16324 22260
rect 16268 22206 16270 22258
rect 16270 22206 16322 22258
rect 16322 22206 16324 22258
rect 16268 22204 16324 22206
rect 15932 21586 15988 21588
rect 15932 21534 15934 21586
rect 15934 21534 15986 21586
rect 15986 21534 15988 21586
rect 15932 21532 15988 21534
rect 16716 29932 16772 29988
rect 16716 29426 16772 29428
rect 16716 29374 16718 29426
rect 16718 29374 16770 29426
rect 16770 29374 16772 29426
rect 16716 29372 16772 29374
rect 16604 29314 16660 29316
rect 16604 29262 16606 29314
rect 16606 29262 16658 29314
rect 16658 29262 16660 29314
rect 16604 29260 16660 29262
rect 16828 28924 16884 28980
rect 17052 30828 17108 30884
rect 17388 30380 17444 30436
rect 17276 30210 17332 30212
rect 17276 30158 17278 30210
rect 17278 30158 17330 30210
rect 17330 30158 17332 30210
rect 17276 30156 17332 30158
rect 17612 30044 17668 30100
rect 17500 29650 17556 29652
rect 17500 29598 17502 29650
rect 17502 29598 17554 29650
rect 17554 29598 17556 29650
rect 17500 29596 17556 29598
rect 17500 29036 17556 29092
rect 17164 28418 17220 28420
rect 17164 28366 17166 28418
rect 17166 28366 17218 28418
rect 17218 28366 17220 28418
rect 17164 28364 17220 28366
rect 16828 27804 16884 27860
rect 16492 27634 16548 27636
rect 16492 27582 16494 27634
rect 16494 27582 16546 27634
rect 16546 27582 16548 27634
rect 16492 27580 16548 27582
rect 16828 26962 16884 26964
rect 16828 26910 16830 26962
rect 16830 26910 16882 26962
rect 16882 26910 16884 26962
rect 16828 26908 16884 26910
rect 17388 26908 17444 26964
rect 16380 21196 16436 21252
rect 16492 25676 16548 25732
rect 16716 25506 16772 25508
rect 16716 25454 16718 25506
rect 16718 25454 16770 25506
rect 16770 25454 16772 25506
rect 16716 25452 16772 25454
rect 16716 24892 16772 24948
rect 17836 29260 17892 29316
rect 18284 29260 18340 29316
rect 18396 28364 18452 28420
rect 17836 27858 17892 27860
rect 17836 27806 17838 27858
rect 17838 27806 17890 27858
rect 17890 27806 17892 27858
rect 17836 27804 17892 27806
rect 16604 24556 16660 24612
rect 16716 24444 16772 24500
rect 17500 24332 17556 24388
rect 17612 27580 17668 27636
rect 16716 23938 16772 23940
rect 16716 23886 16718 23938
rect 16718 23886 16770 23938
rect 16770 23886 16772 23938
rect 16716 23884 16772 23886
rect 17500 23324 17556 23380
rect 16604 23042 16660 23044
rect 16604 22990 16606 23042
rect 16606 22990 16658 23042
rect 16658 22990 16660 23042
rect 16604 22988 16660 22990
rect 16380 20636 16436 20692
rect 16380 20018 16436 20020
rect 16380 19966 16382 20018
rect 16382 19966 16434 20018
rect 16434 19966 16436 20018
rect 16380 19964 16436 19966
rect 16268 19852 16324 19908
rect 16156 19740 16212 19796
rect 15820 19628 15876 19684
rect 15372 18284 15428 18340
rect 15036 18226 15092 18228
rect 15036 18174 15038 18226
rect 15038 18174 15090 18226
rect 15090 18174 15092 18226
rect 15036 18172 15092 18174
rect 14924 17164 14980 17220
rect 14700 15874 14756 15876
rect 14700 15822 14702 15874
rect 14702 15822 14754 15874
rect 14754 15822 14756 15874
rect 14700 15820 14756 15822
rect 14588 15314 14644 15316
rect 14588 15262 14590 15314
rect 14590 15262 14642 15314
rect 14642 15262 14644 15314
rect 14588 15260 14644 15262
rect 14700 15202 14756 15204
rect 14700 15150 14702 15202
rect 14702 15150 14754 15202
rect 14754 15150 14756 15202
rect 14700 15148 14756 15150
rect 13916 13522 13972 13524
rect 13916 13470 13918 13522
rect 13918 13470 13970 13522
rect 13970 13470 13972 13522
rect 13916 13468 13972 13470
rect 14028 12850 14084 12852
rect 14028 12798 14030 12850
rect 14030 12798 14082 12850
rect 14082 12798 14084 12850
rect 14028 12796 14084 12798
rect 13804 11788 13860 11844
rect 14028 11116 14084 11172
rect 13580 9826 13636 9828
rect 13580 9774 13582 9826
rect 13582 9774 13634 9826
rect 13634 9774 13636 9826
rect 13580 9772 13636 9774
rect 13580 9154 13636 9156
rect 13580 9102 13582 9154
rect 13582 9102 13634 9154
rect 13634 9102 13636 9154
rect 13580 9100 13636 9102
rect 13468 8428 13524 8484
rect 13580 7644 13636 7700
rect 13132 6860 13188 6916
rect 14252 9938 14308 9940
rect 14252 9886 14254 9938
rect 14254 9886 14306 9938
rect 14306 9886 14308 9938
rect 14252 9884 14308 9886
rect 13916 9324 13972 9380
rect 14028 9154 14084 9156
rect 14028 9102 14030 9154
rect 14030 9102 14082 9154
rect 14082 9102 14084 9154
rect 14028 9100 14084 9102
rect 13804 7420 13860 7476
rect 14028 7084 14084 7140
rect 14252 7644 14308 7700
rect 15036 15148 15092 15204
rect 15260 15372 15316 15428
rect 14924 14364 14980 14420
rect 15260 14364 15316 14420
rect 14924 13468 14980 13524
rect 15036 13356 15092 13412
rect 15708 17666 15764 17668
rect 15708 17614 15710 17666
rect 15710 17614 15762 17666
rect 15762 17614 15764 17666
rect 15708 17612 15764 17614
rect 15708 17276 15764 17332
rect 15708 16940 15764 16996
rect 15596 16044 15652 16100
rect 15708 16770 15764 16772
rect 15708 16718 15710 16770
rect 15710 16718 15762 16770
rect 15762 16718 15764 16770
rect 15708 16716 15764 16718
rect 16044 19010 16100 19012
rect 16044 18958 16046 19010
rect 16046 18958 16098 19010
rect 16098 18958 16100 19010
rect 16044 18956 16100 18958
rect 15932 18732 15988 18788
rect 17052 22204 17108 22260
rect 16828 21868 16884 21924
rect 16604 21810 16660 21812
rect 16604 21758 16606 21810
rect 16606 21758 16658 21810
rect 16658 21758 16660 21810
rect 16604 21756 16660 21758
rect 16940 21644 16996 21700
rect 16716 21196 16772 21252
rect 16716 20690 16772 20692
rect 16716 20638 16718 20690
rect 16718 20638 16770 20690
rect 16770 20638 16772 20690
rect 16716 20636 16772 20638
rect 16604 20300 16660 20356
rect 16940 20860 16996 20916
rect 16604 19628 16660 19684
rect 16380 18844 16436 18900
rect 16156 18338 16212 18340
rect 16156 18286 16158 18338
rect 16158 18286 16210 18338
rect 16210 18286 16212 18338
rect 16156 18284 16212 18286
rect 16156 17836 16212 17892
rect 15932 17554 15988 17556
rect 15932 17502 15934 17554
rect 15934 17502 15986 17554
rect 15986 17502 15988 17554
rect 15932 17500 15988 17502
rect 15820 16156 15876 16212
rect 16268 17442 16324 17444
rect 16268 17390 16270 17442
rect 16270 17390 16322 17442
rect 16322 17390 16324 17442
rect 16268 17388 16324 17390
rect 16492 18060 16548 18116
rect 16828 19068 16884 19124
rect 16716 18620 16772 18676
rect 17388 21644 17444 21700
rect 17276 21532 17332 21588
rect 17276 20636 17332 20692
rect 17164 20578 17220 20580
rect 17164 20526 17166 20578
rect 17166 20526 17218 20578
rect 17218 20526 17220 20578
rect 17164 20524 17220 20526
rect 17164 19852 17220 19908
rect 17276 19740 17332 19796
rect 17500 19906 17556 19908
rect 17500 19854 17502 19906
rect 17502 19854 17554 19906
rect 17554 19854 17556 19906
rect 17500 19852 17556 19854
rect 18172 27356 18228 27412
rect 18284 27580 18340 27636
rect 18620 29596 18676 29652
rect 18732 27970 18788 27972
rect 18732 27918 18734 27970
rect 18734 27918 18786 27970
rect 18786 27918 18788 27970
rect 18732 27916 18788 27918
rect 18620 27468 18676 27524
rect 17724 24610 17780 24612
rect 17724 24558 17726 24610
rect 17726 24558 17778 24610
rect 17778 24558 17780 24610
rect 17724 24556 17780 24558
rect 17948 24556 18004 24612
rect 17948 23996 18004 24052
rect 18172 26012 18228 26068
rect 20524 33180 20580 33236
rect 20300 33122 20356 33124
rect 20300 33070 20302 33122
rect 20302 33070 20354 33122
rect 20354 33070 20356 33122
rect 20300 33068 20356 33070
rect 20860 33404 20916 33460
rect 22092 36876 22148 36932
rect 24780 36428 24836 36484
rect 22092 36316 22148 36372
rect 21868 35644 21924 35700
rect 21868 34860 21924 34916
rect 24108 36370 24164 36372
rect 24108 36318 24110 36370
rect 24110 36318 24162 36370
rect 24162 36318 24164 36370
rect 24108 36316 24164 36318
rect 22204 34802 22260 34804
rect 22204 34750 22206 34802
rect 22206 34750 22258 34802
rect 22258 34750 22260 34802
rect 22204 34748 22260 34750
rect 20636 33068 20692 33124
rect 19292 32844 19348 32900
rect 20532 32954 20588 32956
rect 20532 32902 20534 32954
rect 20534 32902 20586 32954
rect 20586 32902 20588 32954
rect 20532 32900 20588 32902
rect 20636 32954 20692 32956
rect 20636 32902 20638 32954
rect 20638 32902 20690 32954
rect 20690 32902 20692 32954
rect 20636 32900 20692 32902
rect 20740 32954 20796 32956
rect 20740 32902 20742 32954
rect 20742 32902 20794 32954
rect 20794 32902 20796 32954
rect 20740 32900 20796 32902
rect 19292 32562 19348 32564
rect 19292 32510 19294 32562
rect 19294 32510 19346 32562
rect 19346 32510 19348 32562
rect 19292 32508 19348 32510
rect 19516 32396 19572 32452
rect 19964 32562 20020 32564
rect 19964 32510 19966 32562
rect 19966 32510 20018 32562
rect 20018 32510 20020 32562
rect 19964 32508 20020 32510
rect 19068 31388 19124 31444
rect 19404 31276 19460 31332
rect 19068 30322 19124 30324
rect 19068 30270 19070 30322
rect 19070 30270 19122 30322
rect 19122 30270 19124 30322
rect 19068 30268 19124 30270
rect 19292 30156 19348 30212
rect 19180 30044 19236 30100
rect 19068 29932 19124 29988
rect 19516 30210 19572 30212
rect 19516 30158 19518 30210
rect 19518 30158 19570 30210
rect 19570 30158 19572 30210
rect 19516 30156 19572 30158
rect 19628 29932 19684 29988
rect 19292 29036 19348 29092
rect 19068 27804 19124 27860
rect 19292 28082 19348 28084
rect 19292 28030 19294 28082
rect 19294 28030 19346 28082
rect 19346 28030 19348 28082
rect 19292 28028 19348 28030
rect 19292 27580 19348 27636
rect 18732 26178 18788 26180
rect 18732 26126 18734 26178
rect 18734 26126 18786 26178
rect 18786 26126 18788 26178
rect 18732 26124 18788 26126
rect 18732 25900 18788 25956
rect 18732 24722 18788 24724
rect 18732 24670 18734 24722
rect 18734 24670 18786 24722
rect 18786 24670 18788 24722
rect 18732 24668 18788 24670
rect 18732 24220 18788 24276
rect 18396 23996 18452 24052
rect 20412 32450 20468 32452
rect 20412 32398 20414 32450
rect 20414 32398 20466 32450
rect 20466 32398 20468 32450
rect 20412 32396 20468 32398
rect 19852 31106 19908 31108
rect 19852 31054 19854 31106
rect 19854 31054 19906 31106
rect 19906 31054 19908 31106
rect 19852 31052 19908 31054
rect 20076 31106 20132 31108
rect 20076 31054 20078 31106
rect 20078 31054 20130 31106
rect 20130 31054 20132 31106
rect 20076 31052 20132 31054
rect 20076 30716 20132 30772
rect 20188 30492 20244 30548
rect 20188 30156 20244 30212
rect 19740 29314 19796 29316
rect 19740 29262 19742 29314
rect 19742 29262 19794 29314
rect 19794 29262 19796 29314
rect 19740 29260 19796 29262
rect 19628 27468 19684 27524
rect 20532 31386 20588 31388
rect 20532 31334 20534 31386
rect 20534 31334 20586 31386
rect 20586 31334 20588 31386
rect 20532 31332 20588 31334
rect 20636 31386 20692 31388
rect 20636 31334 20638 31386
rect 20638 31334 20690 31386
rect 20690 31334 20692 31386
rect 20636 31332 20692 31334
rect 20740 31386 20796 31388
rect 20740 31334 20742 31386
rect 20742 31334 20794 31386
rect 20794 31334 20796 31386
rect 20740 31332 20796 31334
rect 20748 30492 20804 30548
rect 20300 30044 20356 30100
rect 20524 30098 20580 30100
rect 20524 30046 20526 30098
rect 20526 30046 20578 30098
rect 20578 30046 20580 30098
rect 20524 30044 20580 30046
rect 20532 29818 20588 29820
rect 20532 29766 20534 29818
rect 20534 29766 20586 29818
rect 20586 29766 20588 29818
rect 20532 29764 20588 29766
rect 20636 29818 20692 29820
rect 20636 29766 20638 29818
rect 20638 29766 20690 29818
rect 20690 29766 20692 29818
rect 20636 29764 20692 29766
rect 20740 29818 20796 29820
rect 20740 29766 20742 29818
rect 20742 29766 20794 29818
rect 20794 29766 20796 29818
rect 20740 29764 20796 29766
rect 20300 29596 20356 29652
rect 20748 29650 20804 29652
rect 20748 29598 20750 29650
rect 20750 29598 20802 29650
rect 20802 29598 20804 29650
rect 20748 29596 20804 29598
rect 20636 29538 20692 29540
rect 20636 29486 20638 29538
rect 20638 29486 20690 29538
rect 20690 29486 20692 29538
rect 20636 29484 20692 29486
rect 21868 33404 21924 33460
rect 20972 32956 21028 33012
rect 20972 32786 21028 32788
rect 20972 32734 20974 32786
rect 20974 32734 21026 32786
rect 21026 32734 21028 32786
rect 20972 32732 21028 32734
rect 21644 33234 21700 33236
rect 21644 33182 21646 33234
rect 21646 33182 21698 33234
rect 21698 33182 21700 33234
rect 21644 33180 21700 33182
rect 22092 33068 22148 33124
rect 21532 32956 21588 33012
rect 21308 32620 21364 32676
rect 21308 30828 21364 30884
rect 21420 30716 21476 30772
rect 21196 30044 21252 30100
rect 20524 29148 20580 29204
rect 20748 28924 20804 28980
rect 20076 27970 20132 27972
rect 20076 27918 20078 27970
rect 20078 27918 20130 27970
rect 20130 27918 20132 27970
rect 20076 27916 20132 27918
rect 20188 27356 20244 27412
rect 19964 27020 20020 27076
rect 19852 26460 19908 26516
rect 19404 26290 19460 26292
rect 19404 26238 19406 26290
rect 19406 26238 19458 26290
rect 19458 26238 19460 26290
rect 19404 26236 19460 26238
rect 19068 26066 19124 26068
rect 19068 26014 19070 26066
rect 19070 26014 19122 26066
rect 19122 26014 19124 26066
rect 19068 26012 19124 26014
rect 18956 25900 19012 25956
rect 19404 24722 19460 24724
rect 19404 24670 19406 24722
rect 19406 24670 19458 24722
rect 19458 24670 19460 24722
rect 19404 24668 19460 24670
rect 19068 24498 19124 24500
rect 19068 24446 19070 24498
rect 19070 24446 19122 24498
rect 19122 24446 19124 24498
rect 19068 24444 19124 24446
rect 18172 22876 18228 22932
rect 19068 23266 19124 23268
rect 19068 23214 19070 23266
rect 19070 23214 19122 23266
rect 19122 23214 19124 23266
rect 19068 23212 19124 23214
rect 18284 22428 18340 22484
rect 18732 22540 18788 22596
rect 18396 22146 18452 22148
rect 18396 22094 18398 22146
rect 18398 22094 18450 22146
rect 18450 22094 18452 22146
rect 18396 22092 18452 22094
rect 18396 21868 18452 21924
rect 17836 21084 17892 21140
rect 18284 21308 18340 21364
rect 17836 20914 17892 20916
rect 17836 20862 17838 20914
rect 17838 20862 17890 20914
rect 17890 20862 17892 20914
rect 17836 20860 17892 20862
rect 18284 20748 18340 20804
rect 18508 21810 18564 21812
rect 18508 21758 18510 21810
rect 18510 21758 18562 21810
rect 18562 21758 18564 21810
rect 18508 21756 18564 21758
rect 18732 21698 18788 21700
rect 18732 21646 18734 21698
rect 18734 21646 18786 21698
rect 18786 21646 18788 21698
rect 18732 21644 18788 21646
rect 18284 20578 18340 20580
rect 18284 20526 18286 20578
rect 18286 20526 18338 20578
rect 18338 20526 18340 20578
rect 18284 20524 18340 20526
rect 18620 21084 18676 21140
rect 18508 20524 18564 20580
rect 16828 18508 16884 18564
rect 16828 18338 16884 18340
rect 16828 18286 16830 18338
rect 16830 18286 16882 18338
rect 16882 18286 16884 18338
rect 16828 18284 16884 18286
rect 17836 19068 17892 19124
rect 17388 18844 17444 18900
rect 17164 18172 17220 18228
rect 16716 17554 16772 17556
rect 16716 17502 16718 17554
rect 16718 17502 16770 17554
rect 16770 17502 16772 17554
rect 16716 17500 16772 17502
rect 16268 16994 16324 16996
rect 16268 16942 16270 16994
rect 16270 16942 16322 16994
rect 16322 16942 16324 16994
rect 16268 16940 16324 16942
rect 16380 16882 16436 16884
rect 16380 16830 16382 16882
rect 16382 16830 16434 16882
rect 16434 16830 16436 16882
rect 16380 16828 16436 16830
rect 15708 15484 15764 15540
rect 15260 13132 15316 13188
rect 14364 6748 14420 6804
rect 14476 9772 14532 9828
rect 15148 11788 15204 11844
rect 13132 6130 13188 6132
rect 13132 6078 13134 6130
rect 13134 6078 13186 6130
rect 13186 6078 13188 6130
rect 13132 6076 13188 6078
rect 13580 5852 13636 5908
rect 12908 5234 12964 5236
rect 12908 5182 12910 5234
rect 12910 5182 12962 5234
rect 12962 5182 12964 5234
rect 12908 5180 12964 5182
rect 12796 4956 12852 5012
rect 14252 6130 14308 6132
rect 14252 6078 14254 6130
rect 14254 6078 14306 6130
rect 14306 6078 14308 6130
rect 14252 6076 14308 6078
rect 14252 5628 14308 5684
rect 16716 17164 16772 17220
rect 16156 15426 16212 15428
rect 16156 15374 16158 15426
rect 16158 15374 16210 15426
rect 16210 15374 16212 15426
rect 16156 15372 16212 15374
rect 15932 14140 15988 14196
rect 15708 13132 15764 13188
rect 16044 13746 16100 13748
rect 16044 13694 16046 13746
rect 16046 13694 16098 13746
rect 16098 13694 16100 13746
rect 16044 13692 16100 13694
rect 17164 17836 17220 17892
rect 17836 18844 17892 18900
rect 17500 17890 17556 17892
rect 17500 17838 17502 17890
rect 17502 17838 17554 17890
rect 17554 17838 17556 17890
rect 17500 17836 17556 17838
rect 18060 17948 18116 18004
rect 18396 19180 18452 19236
rect 18284 19122 18340 19124
rect 18284 19070 18286 19122
rect 18286 19070 18338 19122
rect 18338 19070 18340 19122
rect 18284 19068 18340 19070
rect 18396 18844 18452 18900
rect 18956 20578 19012 20580
rect 18956 20526 18958 20578
rect 18958 20526 19010 20578
rect 19010 20526 19012 20578
rect 18956 20524 19012 20526
rect 18732 20412 18788 20468
rect 18620 19234 18676 19236
rect 18620 19182 18622 19234
rect 18622 19182 18674 19234
rect 18674 19182 18676 19234
rect 18620 19180 18676 19182
rect 19068 20412 19124 20468
rect 19852 26290 19908 26292
rect 19852 26238 19854 26290
rect 19854 26238 19906 26290
rect 19906 26238 19908 26290
rect 19852 26236 19908 26238
rect 19740 24892 19796 24948
rect 19628 24332 19684 24388
rect 19852 24220 19908 24276
rect 20076 26236 20132 26292
rect 20076 26012 20132 26068
rect 20188 24780 20244 24836
rect 20972 28812 21028 28868
rect 21084 28700 21140 28756
rect 20860 28588 20916 28644
rect 20532 28250 20588 28252
rect 20532 28198 20534 28250
rect 20534 28198 20586 28250
rect 20586 28198 20588 28250
rect 20532 28196 20588 28198
rect 20636 28250 20692 28252
rect 20636 28198 20638 28250
rect 20638 28198 20690 28250
rect 20690 28198 20692 28250
rect 20636 28196 20692 28198
rect 20740 28250 20796 28252
rect 20740 28198 20742 28250
rect 20742 28198 20794 28250
rect 20794 28198 20796 28250
rect 20740 28196 20796 28198
rect 20748 28028 20804 28084
rect 20524 27746 20580 27748
rect 20524 27694 20526 27746
rect 20526 27694 20578 27746
rect 20578 27694 20580 27746
rect 20524 27692 20580 27694
rect 20524 27132 20580 27188
rect 20748 27020 20804 27076
rect 20532 26682 20588 26684
rect 20532 26630 20534 26682
rect 20534 26630 20586 26682
rect 20586 26630 20588 26682
rect 20532 26628 20588 26630
rect 20636 26682 20692 26684
rect 20636 26630 20638 26682
rect 20638 26630 20690 26682
rect 20690 26630 20692 26682
rect 20636 26628 20692 26630
rect 20740 26682 20796 26684
rect 20740 26630 20742 26682
rect 20742 26630 20794 26682
rect 20794 26630 20796 26682
rect 20740 26628 20796 26630
rect 20636 26012 20692 26068
rect 20748 25506 20804 25508
rect 20748 25454 20750 25506
rect 20750 25454 20802 25506
rect 20802 25454 20804 25506
rect 20748 25452 20804 25454
rect 20532 25114 20588 25116
rect 20532 25062 20534 25114
rect 20534 25062 20586 25114
rect 20586 25062 20588 25114
rect 20532 25060 20588 25062
rect 20636 25114 20692 25116
rect 20636 25062 20638 25114
rect 20638 25062 20690 25114
rect 20690 25062 20692 25114
rect 20636 25060 20692 25062
rect 20740 25114 20796 25116
rect 20740 25062 20742 25114
rect 20742 25062 20794 25114
rect 20794 25062 20796 25114
rect 20740 25060 20796 25062
rect 19740 23212 19796 23268
rect 19404 22482 19460 22484
rect 19404 22430 19406 22482
rect 19406 22430 19458 22482
rect 19458 22430 19460 22482
rect 19404 22428 19460 22430
rect 19852 23100 19908 23156
rect 19852 22540 19908 22596
rect 19292 21756 19348 21812
rect 19292 21586 19348 21588
rect 19292 21534 19294 21586
rect 19294 21534 19346 21586
rect 19346 21534 19348 21586
rect 19292 21532 19348 21534
rect 19404 21420 19460 21476
rect 19628 21084 19684 21140
rect 19404 20524 19460 20580
rect 18172 17724 18228 17780
rect 16828 16210 16884 16212
rect 16828 16158 16830 16210
rect 16830 16158 16882 16210
rect 16882 16158 16884 16210
rect 16828 16156 16884 16158
rect 17052 17388 17108 17444
rect 17164 16828 17220 16884
rect 16940 15932 16996 15988
rect 16604 15260 16660 15316
rect 16268 13020 16324 13076
rect 15820 12684 15876 12740
rect 15484 11788 15540 11844
rect 15708 12178 15764 12180
rect 15708 12126 15710 12178
rect 15710 12126 15762 12178
rect 15762 12126 15764 12178
rect 15708 12124 15764 12126
rect 15820 12066 15876 12068
rect 15820 12014 15822 12066
rect 15822 12014 15874 12066
rect 15874 12014 15876 12066
rect 15820 12012 15876 12014
rect 15484 11282 15540 11284
rect 15484 11230 15486 11282
rect 15486 11230 15538 11282
rect 15538 11230 15540 11282
rect 15484 11228 15540 11230
rect 15484 10220 15540 10276
rect 15372 9884 15428 9940
rect 15708 10498 15764 10500
rect 15708 10446 15710 10498
rect 15710 10446 15762 10498
rect 15762 10446 15764 10498
rect 15708 10444 15764 10446
rect 16156 12738 16212 12740
rect 16156 12686 16158 12738
rect 16158 12686 16210 12738
rect 16210 12686 16212 12738
rect 16156 12684 16212 12686
rect 16268 12012 16324 12068
rect 16716 14700 16772 14756
rect 16828 14476 16884 14532
rect 16492 12124 16548 12180
rect 16716 12572 16772 12628
rect 16492 11340 16548 11396
rect 15932 10780 15988 10836
rect 16044 10386 16100 10388
rect 16044 10334 16046 10386
rect 16046 10334 16098 10386
rect 16098 10334 16100 10386
rect 16044 10332 16100 10334
rect 15708 10220 15764 10276
rect 16940 13916 16996 13972
rect 18620 18396 18676 18452
rect 18508 18284 18564 18340
rect 18396 17164 18452 17220
rect 18956 18620 19012 18676
rect 19068 18562 19124 18564
rect 19068 18510 19070 18562
rect 19070 18510 19122 18562
rect 19122 18510 19124 18562
rect 19068 18508 19124 18510
rect 18956 18396 19012 18452
rect 18844 17442 18900 17444
rect 18844 17390 18846 17442
rect 18846 17390 18898 17442
rect 18898 17390 18900 17442
rect 18844 17388 18900 17390
rect 18844 16940 18900 16996
rect 17948 15932 18004 15988
rect 17388 14700 17444 14756
rect 17164 14306 17220 14308
rect 17164 14254 17166 14306
rect 17166 14254 17218 14306
rect 17218 14254 17220 14306
rect 17164 14252 17220 14254
rect 17612 14924 17668 14980
rect 17500 14476 17556 14532
rect 17724 14476 17780 14532
rect 18396 15202 18452 15204
rect 18396 15150 18398 15202
rect 18398 15150 18450 15202
rect 18450 15150 18452 15202
rect 18396 15148 18452 15150
rect 18060 14924 18116 14980
rect 17948 14306 18004 14308
rect 17948 14254 17950 14306
rect 17950 14254 18002 14306
rect 18002 14254 18004 14306
rect 17948 14252 18004 14254
rect 17836 13970 17892 13972
rect 17836 13918 17838 13970
rect 17838 13918 17890 13970
rect 17890 13918 17892 13970
rect 17836 13916 17892 13918
rect 16940 13074 16996 13076
rect 16940 13022 16942 13074
rect 16942 13022 16994 13074
rect 16994 13022 16996 13074
rect 16940 13020 16996 13022
rect 17724 13746 17780 13748
rect 17724 13694 17726 13746
rect 17726 13694 17778 13746
rect 17778 13694 17780 13746
rect 17724 13692 17780 13694
rect 17612 13468 17668 13524
rect 17836 13580 17892 13636
rect 18396 14924 18452 14980
rect 18284 14642 18340 14644
rect 18284 14590 18286 14642
rect 18286 14590 18338 14642
rect 18338 14590 18340 14642
rect 18284 14588 18340 14590
rect 18060 13580 18116 13636
rect 18284 13468 18340 13524
rect 17276 12684 17332 12740
rect 16828 12460 16884 12516
rect 17276 11564 17332 11620
rect 16828 11394 16884 11396
rect 16828 11342 16830 11394
rect 16830 11342 16882 11394
rect 16882 11342 16884 11394
rect 16828 11340 16884 11342
rect 16940 11228 16996 11284
rect 16380 11170 16436 11172
rect 16380 11118 16382 11170
rect 16382 11118 16434 11170
rect 16434 11118 16436 11170
rect 16380 11116 16436 11118
rect 17836 12850 17892 12852
rect 17836 12798 17838 12850
rect 17838 12798 17890 12850
rect 17890 12798 17892 12850
rect 17836 12796 17892 12798
rect 17948 12572 18004 12628
rect 17612 11564 17668 11620
rect 17500 11116 17556 11172
rect 18060 11116 18116 11172
rect 17276 10834 17332 10836
rect 17276 10782 17278 10834
rect 17278 10782 17330 10834
rect 17330 10782 17332 10834
rect 17276 10780 17332 10782
rect 17500 10444 17556 10500
rect 17388 10220 17444 10276
rect 17836 9714 17892 9716
rect 17836 9662 17838 9714
rect 17838 9662 17890 9714
rect 17890 9662 17892 9714
rect 17836 9660 17892 9662
rect 16156 8540 16212 8596
rect 17276 8540 17332 8596
rect 15148 7196 15204 7252
rect 18284 13020 18340 13076
rect 18732 16492 18788 16548
rect 19180 18060 19236 18116
rect 18956 16380 19012 16436
rect 18956 16098 19012 16100
rect 18956 16046 18958 16098
rect 18958 16046 19010 16098
rect 19010 16046 19012 16098
rect 18956 16044 19012 16046
rect 19292 16380 19348 16436
rect 19068 14924 19124 14980
rect 18844 14588 18900 14644
rect 18956 14530 19012 14532
rect 18956 14478 18958 14530
rect 18958 14478 19010 14530
rect 19010 14478 19012 14530
rect 18956 14476 19012 14478
rect 19180 13916 19236 13972
rect 18284 12460 18340 12516
rect 18284 11788 18340 11844
rect 18396 11676 18452 11732
rect 18620 12012 18676 12068
rect 18620 11282 18676 11284
rect 18620 11230 18622 11282
rect 18622 11230 18674 11282
rect 18674 11230 18676 11282
rect 18620 11228 18676 11230
rect 18844 12850 18900 12852
rect 18844 12798 18846 12850
rect 18846 12798 18898 12850
rect 18898 12798 18900 12850
rect 18844 12796 18900 12798
rect 19516 19852 19572 19908
rect 19740 20578 19796 20580
rect 19740 20526 19742 20578
rect 19742 20526 19794 20578
rect 19794 20526 19796 20578
rect 19740 20524 19796 20526
rect 20524 23884 20580 23940
rect 20188 23772 20244 23828
rect 20532 23546 20588 23548
rect 20188 23436 20244 23492
rect 20532 23494 20534 23546
rect 20534 23494 20586 23546
rect 20586 23494 20588 23546
rect 20532 23492 20588 23494
rect 20636 23546 20692 23548
rect 20636 23494 20638 23546
rect 20638 23494 20690 23546
rect 20690 23494 20692 23546
rect 20636 23492 20692 23494
rect 20740 23546 20796 23548
rect 20740 23494 20742 23546
rect 20742 23494 20794 23546
rect 20794 23494 20796 23546
rect 20740 23492 20796 23494
rect 20300 22876 20356 22932
rect 20532 21978 20588 21980
rect 20532 21926 20534 21978
rect 20534 21926 20586 21978
rect 20586 21926 20588 21978
rect 20532 21924 20588 21926
rect 20636 21978 20692 21980
rect 20636 21926 20638 21978
rect 20638 21926 20690 21978
rect 20690 21926 20692 21978
rect 20636 21924 20692 21926
rect 20740 21978 20796 21980
rect 20740 21926 20742 21978
rect 20742 21926 20794 21978
rect 20794 21926 20796 21978
rect 20740 21924 20796 21926
rect 20300 21698 20356 21700
rect 20300 21646 20302 21698
rect 20302 21646 20354 21698
rect 20354 21646 20356 21698
rect 20300 21644 20356 21646
rect 20188 21196 20244 21252
rect 20636 20972 20692 21028
rect 21308 28028 21364 28084
rect 21084 27804 21140 27860
rect 21644 29708 21700 29764
rect 21532 29148 21588 29204
rect 21756 29596 21812 29652
rect 21644 28924 21700 28980
rect 21868 27970 21924 27972
rect 21868 27918 21870 27970
rect 21870 27918 21922 27970
rect 21922 27918 21924 27970
rect 21868 27916 21924 27918
rect 21980 29932 22036 29988
rect 22092 29538 22148 29540
rect 22092 29486 22094 29538
rect 22094 29486 22146 29538
rect 22146 29486 22148 29538
rect 22092 29484 22148 29486
rect 23436 34412 23492 34468
rect 22316 34076 22372 34132
rect 22988 34130 23044 34132
rect 22988 34078 22990 34130
rect 22990 34078 23042 34130
rect 23042 34078 23044 34130
rect 22988 34076 23044 34078
rect 25004 35084 25060 35140
rect 23660 34300 23716 34356
rect 24220 34748 24276 34804
rect 24444 34690 24500 34692
rect 24444 34638 24446 34690
rect 24446 34638 24498 34690
rect 24498 34638 24500 34690
rect 24444 34636 24500 34638
rect 24444 34300 24500 34356
rect 23548 33404 23604 33460
rect 22876 33292 22932 33348
rect 24108 33964 24164 34020
rect 22876 32956 22932 33012
rect 22540 32620 22596 32676
rect 22428 30380 22484 30436
rect 23324 33122 23380 33124
rect 23324 33070 23326 33122
rect 23326 33070 23378 33122
rect 23378 33070 23380 33122
rect 23324 33068 23380 33070
rect 24332 33122 24388 33124
rect 24332 33070 24334 33122
rect 24334 33070 24386 33122
rect 24386 33070 24388 33122
rect 24332 33068 24388 33070
rect 23772 32956 23828 33012
rect 23324 31890 23380 31892
rect 23324 31838 23326 31890
rect 23326 31838 23378 31890
rect 23378 31838 23380 31890
rect 23324 31836 23380 31838
rect 22764 31778 22820 31780
rect 22764 31726 22766 31778
rect 22766 31726 22818 31778
rect 22818 31726 22820 31778
rect 22764 31724 22820 31726
rect 22540 29932 22596 29988
rect 22652 30268 22708 30324
rect 21532 27580 21588 27636
rect 21084 26908 21140 26964
rect 21084 26684 21140 26740
rect 21196 26012 21252 26068
rect 21308 24780 21364 24836
rect 21420 26908 21476 26964
rect 21644 27020 21700 27076
rect 21868 26684 21924 26740
rect 21644 25506 21700 25508
rect 21644 25454 21646 25506
rect 21646 25454 21698 25506
rect 21698 25454 21700 25506
rect 21644 25452 21700 25454
rect 21756 23996 21812 24052
rect 22428 29820 22484 29876
rect 22428 29036 22484 29092
rect 22092 28588 22148 28644
rect 22540 28588 22596 28644
rect 22316 28252 22372 28308
rect 22092 26514 22148 26516
rect 22092 26462 22094 26514
rect 22094 26462 22146 26514
rect 22146 26462 22148 26514
rect 22092 26460 22148 26462
rect 21980 25228 22036 25284
rect 22316 25394 22372 25396
rect 22316 25342 22318 25394
rect 22318 25342 22370 25394
rect 22370 25342 22372 25394
rect 22316 25340 22372 25342
rect 22428 26066 22484 26068
rect 22428 26014 22430 26066
rect 22430 26014 22482 26066
rect 22482 26014 22484 26066
rect 22428 26012 22484 26014
rect 22092 24332 22148 24388
rect 21308 23938 21364 23940
rect 21308 23886 21310 23938
rect 21310 23886 21362 23938
rect 21362 23886 21364 23938
rect 21308 23884 21364 23886
rect 21756 23772 21812 23828
rect 21420 23548 21476 23604
rect 21868 23660 21924 23716
rect 21980 23884 22036 23940
rect 21196 22988 21252 23044
rect 21084 20972 21140 21028
rect 19964 20748 20020 20804
rect 20860 20748 20916 20804
rect 20532 20410 20588 20412
rect 20532 20358 20534 20410
rect 20534 20358 20586 20410
rect 20586 20358 20588 20410
rect 20532 20356 20588 20358
rect 20636 20410 20692 20412
rect 20636 20358 20638 20410
rect 20638 20358 20690 20410
rect 20690 20358 20692 20410
rect 20636 20356 20692 20358
rect 20740 20410 20796 20412
rect 20740 20358 20742 20410
rect 20742 20358 20794 20410
rect 20794 20358 20796 20410
rect 20740 20356 20796 20358
rect 20188 19906 20244 19908
rect 20188 19854 20190 19906
rect 20190 19854 20242 19906
rect 20242 19854 20244 19906
rect 20188 19852 20244 19854
rect 20188 18956 20244 19012
rect 20076 18396 20132 18452
rect 20532 18842 20588 18844
rect 20532 18790 20534 18842
rect 20534 18790 20586 18842
rect 20586 18790 20588 18842
rect 20532 18788 20588 18790
rect 20636 18842 20692 18844
rect 20636 18790 20638 18842
rect 20638 18790 20690 18842
rect 20690 18790 20692 18842
rect 20636 18788 20692 18790
rect 20740 18842 20796 18844
rect 20740 18790 20742 18842
rect 20742 18790 20794 18842
rect 20794 18790 20796 18842
rect 20740 18788 20796 18790
rect 20300 18338 20356 18340
rect 20300 18286 20302 18338
rect 20302 18286 20354 18338
rect 20354 18286 20356 18338
rect 20300 18284 20356 18286
rect 20188 17948 20244 18004
rect 20300 17500 20356 17556
rect 19516 15372 19572 15428
rect 19964 17442 20020 17444
rect 19964 17390 19966 17442
rect 19966 17390 20018 17442
rect 20018 17390 20020 17442
rect 19964 17388 20020 17390
rect 19516 12962 19572 12964
rect 19516 12910 19518 12962
rect 19518 12910 19570 12962
rect 19570 12910 19572 12962
rect 19516 12908 19572 12910
rect 18844 11900 18900 11956
rect 19292 12012 19348 12068
rect 19180 11618 19236 11620
rect 19180 11566 19182 11618
rect 19182 11566 19234 11618
rect 19234 11566 19236 11618
rect 19180 11564 19236 11566
rect 19516 11900 19572 11956
rect 18508 10498 18564 10500
rect 18508 10446 18510 10498
rect 18510 10446 18562 10498
rect 18562 10446 18564 10498
rect 18508 10444 18564 10446
rect 18284 8652 18340 8708
rect 18844 9042 18900 9044
rect 18844 8990 18846 9042
rect 18846 8990 18898 9042
rect 18898 8990 18900 9042
rect 18844 8988 18900 8990
rect 18956 8652 19012 8708
rect 15932 7980 15988 8036
rect 17500 7698 17556 7700
rect 17500 7646 17502 7698
rect 17502 7646 17554 7698
rect 17554 7646 17556 7698
rect 17500 7644 17556 7646
rect 15820 6076 15876 6132
rect 16044 6748 16100 6804
rect 14588 5906 14644 5908
rect 14588 5854 14590 5906
rect 14590 5854 14642 5906
rect 14642 5854 14644 5906
rect 14588 5852 14644 5854
rect 13916 5234 13972 5236
rect 13916 5182 13918 5234
rect 13918 5182 13970 5234
rect 13970 5182 13972 5234
rect 13916 5180 13972 5182
rect 14476 5180 14532 5236
rect 13692 4732 13748 4788
rect 14700 5404 14756 5460
rect 15036 5404 15092 5460
rect 15148 5628 15204 5684
rect 14476 4732 14532 4788
rect 14700 4450 14756 4452
rect 14700 4398 14702 4450
rect 14702 4398 14754 4450
rect 14754 4398 14756 4450
rect 14700 4396 14756 4398
rect 11340 2940 11396 2996
rect 15708 5628 15764 5684
rect 15372 4396 15428 4452
rect 15148 2716 15204 2772
rect 16268 5122 16324 5124
rect 16268 5070 16270 5122
rect 16270 5070 16322 5122
rect 16322 5070 16324 5122
rect 16268 5068 16324 5070
rect 16604 4508 16660 4564
rect 16716 5740 16772 5796
rect 17948 8034 18004 8036
rect 17948 7982 17950 8034
rect 17950 7982 18002 8034
rect 18002 7982 18004 8034
rect 17948 7980 18004 7982
rect 18732 7644 18788 7700
rect 18396 5740 18452 5796
rect 17500 5682 17556 5684
rect 17500 5630 17502 5682
rect 17502 5630 17554 5682
rect 17554 5630 17556 5682
rect 17500 5628 17556 5630
rect 16716 4396 16772 4452
rect 17948 5180 18004 5236
rect 17612 4562 17668 4564
rect 17612 4510 17614 4562
rect 17614 4510 17666 4562
rect 17666 4510 17668 4562
rect 17612 4508 17668 4510
rect 19068 8540 19124 8596
rect 19068 8258 19124 8260
rect 19068 8206 19070 8258
rect 19070 8206 19122 8258
rect 19122 8206 19124 8258
rect 19068 8204 19124 8206
rect 19740 16828 19796 16884
rect 20860 18396 20916 18452
rect 20748 18284 20804 18340
rect 21084 18284 21140 18340
rect 20748 17948 20804 18004
rect 20748 17666 20804 17668
rect 20748 17614 20750 17666
rect 20750 17614 20802 17666
rect 20802 17614 20804 17666
rect 20748 17612 20804 17614
rect 20532 17274 20588 17276
rect 20532 17222 20534 17274
rect 20534 17222 20586 17274
rect 20586 17222 20588 17274
rect 20532 17220 20588 17222
rect 20636 17274 20692 17276
rect 20636 17222 20638 17274
rect 20638 17222 20690 17274
rect 20690 17222 20692 17274
rect 20636 17220 20692 17222
rect 20740 17274 20796 17276
rect 20740 17222 20742 17274
rect 20742 17222 20794 17274
rect 20794 17222 20796 17274
rect 20740 17220 20796 17222
rect 19852 15986 19908 15988
rect 19852 15934 19854 15986
rect 19854 15934 19906 15986
rect 19906 15934 19908 15986
rect 19852 15932 19908 15934
rect 20188 15874 20244 15876
rect 20188 15822 20190 15874
rect 20190 15822 20242 15874
rect 20242 15822 20244 15874
rect 20188 15820 20244 15822
rect 20636 15874 20692 15876
rect 20636 15822 20638 15874
rect 20638 15822 20690 15874
rect 20690 15822 20692 15874
rect 20636 15820 20692 15822
rect 20532 15706 20588 15708
rect 20532 15654 20534 15706
rect 20534 15654 20586 15706
rect 20586 15654 20588 15706
rect 20532 15652 20588 15654
rect 20636 15706 20692 15708
rect 20636 15654 20638 15706
rect 20638 15654 20690 15706
rect 20690 15654 20692 15706
rect 20636 15652 20692 15654
rect 20740 15706 20796 15708
rect 20740 15654 20742 15706
rect 20742 15654 20794 15706
rect 20794 15654 20796 15706
rect 20740 15652 20796 15654
rect 20412 15148 20468 15204
rect 21420 21532 21476 21588
rect 22204 23436 22260 23492
rect 22876 30156 22932 30212
rect 23660 31724 23716 31780
rect 23884 31724 23940 31780
rect 23548 31500 23604 31556
rect 23548 30940 23604 30996
rect 23884 30940 23940 30996
rect 23324 30380 23380 30436
rect 23436 29596 23492 29652
rect 22764 28588 22820 28644
rect 22876 28924 22932 28980
rect 22652 28476 22708 28532
rect 22876 28252 22932 28308
rect 22876 27970 22932 27972
rect 22876 27918 22878 27970
rect 22878 27918 22930 27970
rect 22930 27918 22932 27970
rect 22876 27916 22932 27918
rect 23100 28812 23156 28868
rect 23100 28364 23156 28420
rect 23212 28700 23268 28756
rect 24220 31500 24276 31556
rect 24108 30380 24164 30436
rect 23996 30210 24052 30212
rect 23996 30158 23998 30210
rect 23998 30158 24050 30210
rect 24050 30158 24052 30210
rect 23996 30156 24052 30158
rect 23660 29820 23716 29876
rect 22652 26962 22708 26964
rect 22652 26910 22654 26962
rect 22654 26910 22706 26962
rect 22706 26910 22708 26962
rect 22652 26908 22708 26910
rect 23548 27020 23604 27076
rect 22652 25452 22708 25508
rect 22540 24220 22596 24276
rect 22988 25452 23044 25508
rect 23884 28642 23940 28644
rect 23884 28590 23886 28642
rect 23886 28590 23938 28642
rect 23938 28590 23940 28642
rect 23884 28588 23940 28590
rect 23772 28364 23828 28420
rect 23548 24722 23604 24724
rect 23548 24670 23550 24722
rect 23550 24670 23602 24722
rect 23602 24670 23604 24722
rect 23548 24668 23604 24670
rect 23100 23996 23156 24052
rect 22988 23826 23044 23828
rect 22988 23774 22990 23826
rect 22990 23774 23042 23826
rect 23042 23774 23044 23826
rect 22988 23772 23044 23774
rect 23436 24444 23492 24500
rect 22988 23548 23044 23604
rect 23996 27746 24052 27748
rect 23996 27694 23998 27746
rect 23998 27694 24050 27746
rect 24050 27694 24052 27746
rect 23996 27692 24052 27694
rect 23436 23938 23492 23940
rect 23436 23886 23438 23938
rect 23438 23886 23490 23938
rect 23490 23886 23492 23938
rect 23436 23884 23492 23886
rect 23884 24332 23940 24388
rect 23324 23772 23380 23828
rect 22092 22370 22148 22372
rect 22092 22318 22094 22370
rect 22094 22318 22146 22370
rect 22146 22318 22148 22370
rect 22092 22316 22148 22318
rect 21980 22092 22036 22148
rect 21308 20636 21364 20692
rect 21532 20802 21588 20804
rect 21532 20750 21534 20802
rect 21534 20750 21586 20802
rect 21586 20750 21588 20802
rect 21532 20748 21588 20750
rect 21756 20690 21812 20692
rect 21756 20638 21758 20690
rect 21758 20638 21810 20690
rect 21810 20638 21812 20690
rect 21756 20636 21812 20638
rect 21868 19852 21924 19908
rect 22092 20636 22148 20692
rect 22428 21474 22484 21476
rect 22428 21422 22430 21474
rect 22430 21422 22482 21474
rect 22482 21422 22484 21474
rect 22428 21420 22484 21422
rect 21980 19628 22036 19684
rect 21868 19516 21924 19572
rect 22316 19516 22372 19572
rect 21644 19122 21700 19124
rect 21644 19070 21646 19122
rect 21646 19070 21698 19122
rect 21698 19070 21700 19122
rect 21644 19068 21700 19070
rect 21980 19068 22036 19124
rect 21868 19010 21924 19012
rect 21868 18958 21870 19010
rect 21870 18958 21922 19010
rect 21922 18958 21924 19010
rect 21868 18956 21924 18958
rect 21980 18844 22036 18900
rect 21756 18508 21812 18564
rect 21644 17612 21700 17668
rect 21420 17500 21476 17556
rect 21532 15484 21588 15540
rect 20860 14924 20916 14980
rect 20188 14252 20244 14308
rect 20076 14028 20132 14084
rect 20076 12796 20132 12852
rect 19964 12684 20020 12740
rect 19740 11676 19796 11732
rect 20076 12124 20132 12180
rect 20532 14138 20588 14140
rect 20532 14086 20534 14138
rect 20534 14086 20586 14138
rect 20586 14086 20588 14138
rect 20532 14084 20588 14086
rect 20636 14138 20692 14140
rect 20636 14086 20638 14138
rect 20638 14086 20690 14138
rect 20690 14086 20692 14138
rect 20636 14084 20692 14086
rect 20740 14138 20796 14140
rect 20740 14086 20742 14138
rect 20742 14086 20794 14138
rect 20794 14086 20796 14138
rect 20740 14084 20796 14086
rect 21308 14306 21364 14308
rect 21308 14254 21310 14306
rect 21310 14254 21362 14306
rect 21362 14254 21364 14306
rect 21308 14252 21364 14254
rect 20860 13804 20916 13860
rect 20188 13580 20244 13636
rect 20076 11954 20132 11956
rect 20076 11902 20078 11954
rect 20078 11902 20130 11954
rect 20130 11902 20132 11954
rect 20076 11900 20132 11902
rect 19628 10444 19684 10500
rect 19852 10668 19908 10724
rect 20524 13580 20580 13636
rect 20300 12850 20356 12852
rect 20300 12798 20302 12850
rect 20302 12798 20354 12850
rect 20354 12798 20356 12850
rect 20300 12796 20356 12798
rect 20532 12570 20588 12572
rect 20532 12518 20534 12570
rect 20534 12518 20586 12570
rect 20586 12518 20588 12570
rect 20532 12516 20588 12518
rect 20636 12570 20692 12572
rect 20636 12518 20638 12570
rect 20638 12518 20690 12570
rect 20690 12518 20692 12570
rect 20636 12516 20692 12518
rect 20740 12570 20796 12572
rect 20740 12518 20742 12570
rect 20742 12518 20794 12570
rect 20794 12518 20796 12570
rect 20740 12516 20796 12518
rect 19852 10444 19908 10500
rect 20860 11900 20916 11956
rect 20972 11676 21028 11732
rect 20860 11340 20916 11396
rect 20412 11228 20468 11284
rect 20532 11002 20588 11004
rect 20532 10950 20534 11002
rect 20534 10950 20586 11002
rect 20586 10950 20588 11002
rect 20532 10948 20588 10950
rect 20636 11002 20692 11004
rect 20636 10950 20638 11002
rect 20638 10950 20690 11002
rect 20690 10950 20692 11002
rect 20636 10948 20692 10950
rect 20740 11002 20796 11004
rect 20740 10950 20742 11002
rect 20742 10950 20794 11002
rect 20794 10950 20796 11002
rect 20740 10948 20796 10950
rect 21532 13692 21588 13748
rect 21980 18226 22036 18228
rect 21980 18174 21982 18226
rect 21982 18174 22034 18226
rect 22034 18174 22036 18226
rect 21980 18172 22036 18174
rect 22092 17612 22148 17668
rect 22316 17276 22372 17332
rect 22092 16492 22148 16548
rect 22092 16210 22148 16212
rect 22092 16158 22094 16210
rect 22094 16158 22146 16210
rect 22146 16158 22148 16210
rect 22092 16156 22148 16158
rect 22204 15538 22260 15540
rect 22204 15486 22206 15538
rect 22206 15486 22258 15538
rect 22258 15486 22260 15538
rect 22204 15484 22260 15486
rect 22540 20300 22596 20356
rect 22764 21868 22820 21924
rect 22540 18396 22596 18452
rect 22652 18284 22708 18340
rect 22540 18172 22596 18228
rect 22988 21810 23044 21812
rect 22988 21758 22990 21810
rect 22990 21758 23042 21810
rect 23042 21758 23044 21810
rect 22988 21756 23044 21758
rect 23100 20018 23156 20020
rect 23100 19966 23102 20018
rect 23102 19966 23154 20018
rect 23154 19966 23156 20018
rect 23100 19964 23156 19966
rect 23436 23660 23492 23716
rect 23548 21980 23604 22036
rect 23436 21586 23492 21588
rect 23436 21534 23438 21586
rect 23438 21534 23490 21586
rect 23490 21534 23492 21586
rect 23436 21532 23492 21534
rect 23548 20300 23604 20356
rect 23548 19906 23604 19908
rect 23548 19854 23550 19906
rect 23550 19854 23602 19906
rect 23602 19854 23604 19906
rect 23548 19852 23604 19854
rect 23324 19740 23380 19796
rect 23100 19458 23156 19460
rect 23100 19406 23102 19458
rect 23102 19406 23154 19458
rect 23154 19406 23156 19458
rect 23100 19404 23156 19406
rect 22876 18396 22932 18452
rect 21868 14140 21924 14196
rect 21756 13580 21812 13636
rect 22092 14028 22148 14084
rect 21980 13468 22036 13524
rect 21532 13020 21588 13076
rect 21756 13020 21812 13076
rect 21756 12684 21812 12740
rect 21756 12012 21812 12068
rect 21308 11506 21364 11508
rect 21308 11454 21310 11506
rect 21310 11454 21362 11506
rect 21362 11454 21364 11506
rect 21308 11452 21364 11454
rect 19740 9884 19796 9940
rect 20300 9996 20356 10052
rect 19628 9714 19684 9716
rect 19628 9662 19630 9714
rect 19630 9662 19682 9714
rect 19682 9662 19684 9714
rect 19628 9660 19684 9662
rect 21420 10780 21476 10836
rect 21532 10332 21588 10388
rect 21196 10108 21252 10164
rect 21308 10050 21364 10052
rect 21308 9998 21310 10050
rect 21310 9998 21362 10050
rect 21362 9998 21364 10050
rect 21308 9996 21364 9998
rect 21532 9996 21588 10052
rect 20748 9884 20804 9940
rect 20636 9602 20692 9604
rect 20636 9550 20638 9602
rect 20638 9550 20690 9602
rect 20690 9550 20692 9602
rect 20636 9548 20692 9550
rect 19852 9436 19908 9492
rect 19628 8540 19684 8596
rect 19516 8204 19572 8260
rect 19516 7532 19572 7588
rect 19180 6412 19236 6468
rect 19292 5794 19348 5796
rect 19292 5742 19294 5794
rect 19294 5742 19346 5794
rect 19346 5742 19348 5794
rect 19292 5740 19348 5742
rect 18956 5180 19012 5236
rect 18508 4732 18564 4788
rect 18732 4338 18788 4340
rect 18732 4286 18734 4338
rect 18734 4286 18786 4338
rect 18786 4286 18788 4338
rect 18732 4284 18788 4286
rect 19404 4338 19460 4340
rect 19404 4286 19406 4338
rect 19406 4286 19458 4338
rect 19458 4286 19460 4338
rect 19404 4284 19460 4286
rect 19964 8988 20020 9044
rect 20532 9434 20588 9436
rect 20532 9382 20534 9434
rect 20534 9382 20586 9434
rect 20586 9382 20588 9434
rect 20532 9380 20588 9382
rect 20636 9434 20692 9436
rect 20636 9382 20638 9434
rect 20638 9382 20690 9434
rect 20690 9382 20692 9434
rect 20636 9380 20692 9382
rect 20740 9434 20796 9436
rect 20740 9382 20742 9434
rect 20742 9382 20794 9434
rect 20794 9382 20796 9434
rect 20740 9380 20796 9382
rect 20412 8764 20468 8820
rect 20748 9100 20804 9156
rect 21756 10780 21812 10836
rect 21756 10108 21812 10164
rect 21868 9938 21924 9940
rect 21868 9886 21870 9938
rect 21870 9886 21922 9938
rect 21922 9886 21924 9938
rect 21868 9884 21924 9886
rect 22204 12066 22260 12068
rect 22204 12014 22206 12066
rect 22206 12014 22258 12066
rect 22258 12014 22260 12066
rect 22204 12012 22260 12014
rect 22204 11564 22260 11620
rect 22988 18956 23044 19012
rect 23100 18732 23156 18788
rect 23436 18956 23492 19012
rect 23436 18732 23492 18788
rect 23772 23548 23828 23604
rect 24220 29260 24276 29316
rect 24780 33458 24836 33460
rect 24780 33406 24782 33458
rect 24782 33406 24834 33458
rect 24834 33406 24836 33458
rect 24780 33404 24836 33406
rect 26236 36428 26292 36484
rect 26348 36988 26404 37044
rect 25340 36204 25396 36260
rect 25900 35756 25956 35812
rect 29148 36540 29204 36596
rect 27356 36482 27412 36484
rect 27356 36430 27358 36482
rect 27358 36430 27410 36482
rect 27410 36430 27412 36482
rect 27356 36428 27412 36430
rect 28252 36428 28308 36484
rect 27020 36370 27076 36372
rect 27020 36318 27022 36370
rect 27022 36318 27074 36370
rect 27074 36318 27076 36370
rect 27020 36316 27076 36318
rect 26348 35644 26404 35700
rect 25340 35084 25396 35140
rect 26572 35084 26628 35140
rect 27356 35084 27412 35140
rect 25340 34018 25396 34020
rect 25340 33966 25342 34018
rect 25342 33966 25394 34018
rect 25394 33966 25396 34018
rect 25340 33964 25396 33966
rect 25564 33964 25620 34020
rect 25228 33068 25284 33124
rect 25116 32844 25172 32900
rect 25228 32396 25284 32452
rect 25564 33292 25620 33348
rect 27132 34690 27188 34692
rect 27132 34638 27134 34690
rect 27134 34638 27186 34690
rect 27186 34638 27188 34690
rect 27132 34636 27188 34638
rect 27468 34524 27524 34580
rect 25900 34130 25956 34132
rect 25900 34078 25902 34130
rect 25902 34078 25954 34130
rect 25954 34078 25956 34130
rect 25900 34076 25956 34078
rect 26684 33346 26740 33348
rect 26684 33294 26686 33346
rect 26686 33294 26738 33346
rect 26738 33294 26740 33346
rect 26684 33292 26740 33294
rect 25452 32562 25508 32564
rect 25452 32510 25454 32562
rect 25454 32510 25506 32562
rect 25506 32510 25508 32562
rect 25452 32508 25508 32510
rect 25452 31948 25508 32004
rect 24668 31836 24724 31892
rect 25004 31724 25060 31780
rect 25004 31052 25060 31108
rect 26348 33122 26404 33124
rect 26348 33070 26350 33122
rect 26350 33070 26402 33122
rect 26402 33070 26404 33122
rect 26348 33068 26404 33070
rect 26684 32732 26740 32788
rect 27468 32844 27524 32900
rect 26348 32620 26404 32676
rect 24668 30828 24724 30884
rect 24892 30322 24948 30324
rect 24892 30270 24894 30322
rect 24894 30270 24946 30322
rect 24946 30270 24948 30322
rect 24892 30268 24948 30270
rect 25116 29820 25172 29876
rect 26124 32562 26180 32564
rect 26124 32510 26126 32562
rect 26126 32510 26178 32562
rect 26178 32510 26180 32562
rect 26124 32508 26180 32510
rect 27356 32562 27412 32564
rect 27356 32510 27358 32562
rect 27358 32510 27410 32562
rect 27410 32510 27412 32562
rect 27356 32508 27412 32510
rect 26572 32450 26628 32452
rect 26572 32398 26574 32450
rect 26574 32398 26626 32450
rect 26626 32398 26628 32450
rect 26572 32396 26628 32398
rect 25564 30828 25620 30884
rect 25228 29260 25284 29316
rect 24892 28700 24948 28756
rect 24556 28418 24612 28420
rect 24556 28366 24558 28418
rect 24558 28366 24610 28418
rect 24610 28366 24612 28418
rect 24556 28364 24612 28366
rect 24556 28082 24612 28084
rect 24556 28030 24558 28082
rect 24558 28030 24610 28082
rect 24610 28030 24612 28082
rect 24556 28028 24612 28030
rect 24332 27916 24388 27972
rect 24444 27468 24500 27524
rect 24556 26962 24612 26964
rect 24556 26910 24558 26962
rect 24558 26910 24610 26962
rect 24610 26910 24612 26962
rect 24556 26908 24612 26910
rect 24220 25564 24276 25620
rect 24444 24668 24500 24724
rect 23884 21868 23940 21924
rect 24108 21980 24164 22036
rect 24108 21810 24164 21812
rect 24108 21758 24110 21810
rect 24110 21758 24162 21810
rect 24162 21758 24164 21810
rect 24108 21756 24164 21758
rect 24332 21698 24388 21700
rect 24332 21646 24334 21698
rect 24334 21646 24386 21698
rect 24386 21646 24388 21698
rect 24332 21644 24388 21646
rect 23772 21586 23828 21588
rect 23772 21534 23774 21586
rect 23774 21534 23826 21586
rect 23826 21534 23828 21586
rect 23772 21532 23828 21534
rect 23884 21420 23940 21476
rect 23772 20860 23828 20916
rect 23996 19906 24052 19908
rect 23996 19854 23998 19906
rect 23998 19854 24050 19906
rect 24050 19854 24052 19906
rect 23996 19852 24052 19854
rect 24668 21532 24724 21588
rect 24668 21196 24724 21252
rect 23996 19404 24052 19460
rect 24668 20300 24724 20356
rect 24220 18844 24276 18900
rect 23772 18620 23828 18676
rect 23324 18284 23380 18340
rect 23996 18060 24052 18116
rect 23100 17778 23156 17780
rect 23100 17726 23102 17778
rect 23102 17726 23154 17778
rect 23154 17726 23156 17778
rect 23100 17724 23156 17726
rect 23100 17164 23156 17220
rect 23212 17276 23268 17332
rect 22876 16940 22932 16996
rect 22876 15372 22932 15428
rect 23100 13858 23156 13860
rect 23100 13806 23102 13858
rect 23102 13806 23154 13858
rect 23154 13806 23156 13858
rect 23100 13804 23156 13806
rect 24108 17276 24164 17332
rect 24556 17442 24612 17444
rect 24556 17390 24558 17442
rect 24558 17390 24610 17442
rect 24610 17390 24612 17442
rect 24556 17388 24612 17390
rect 24668 17276 24724 17332
rect 24332 17106 24388 17108
rect 24332 17054 24334 17106
rect 24334 17054 24386 17106
rect 24386 17054 24388 17106
rect 24332 17052 24388 17054
rect 23660 16604 23716 16660
rect 23548 15596 23604 15652
rect 24444 16994 24500 16996
rect 24444 16942 24446 16994
rect 24446 16942 24498 16994
rect 24498 16942 24500 16994
rect 24444 16940 24500 16942
rect 23996 15372 24052 15428
rect 23324 13804 23380 13860
rect 23436 15260 23492 15316
rect 23660 15314 23716 15316
rect 23660 15262 23662 15314
rect 23662 15262 23714 15314
rect 23714 15262 23716 15314
rect 23660 15260 23716 15262
rect 24332 16604 24388 16660
rect 22988 13580 23044 13636
rect 23772 14924 23828 14980
rect 22876 13468 22932 13524
rect 22652 12796 22708 12852
rect 22540 11282 22596 11284
rect 22540 11230 22542 11282
rect 22542 11230 22594 11282
rect 22594 11230 22596 11282
rect 22540 11228 22596 11230
rect 22316 10892 22372 10948
rect 22204 10610 22260 10612
rect 22204 10558 22206 10610
rect 22206 10558 22258 10610
rect 22258 10558 22260 10610
rect 22204 10556 22260 10558
rect 22092 9660 22148 9716
rect 20076 8258 20132 8260
rect 20076 8206 20078 8258
rect 20078 8206 20130 8258
rect 20130 8206 20132 8258
rect 20076 8204 20132 8206
rect 21756 8204 21812 8260
rect 21980 8258 22036 8260
rect 21980 8206 21982 8258
rect 21982 8206 22034 8258
rect 22034 8206 22036 8258
rect 21980 8204 22036 8206
rect 20532 7866 20588 7868
rect 20532 7814 20534 7866
rect 20534 7814 20586 7866
rect 20586 7814 20588 7866
rect 20532 7812 20588 7814
rect 20636 7866 20692 7868
rect 20636 7814 20638 7866
rect 20638 7814 20690 7866
rect 20690 7814 20692 7866
rect 20636 7812 20692 7814
rect 20740 7866 20796 7868
rect 20740 7814 20742 7866
rect 20742 7814 20794 7866
rect 20794 7814 20796 7866
rect 20740 7812 20796 7814
rect 20188 7420 20244 7476
rect 20188 6972 20244 7028
rect 19740 6524 19796 6580
rect 19740 6130 19796 6132
rect 19740 6078 19742 6130
rect 19742 6078 19794 6130
rect 19794 6078 19796 6130
rect 19740 6076 19796 6078
rect 19964 5964 20020 6020
rect 20300 6748 20356 6804
rect 20412 6578 20468 6580
rect 20412 6526 20414 6578
rect 20414 6526 20466 6578
rect 20466 6526 20468 6578
rect 20412 6524 20468 6526
rect 20532 6298 20588 6300
rect 20532 6246 20534 6298
rect 20534 6246 20586 6298
rect 20586 6246 20588 6298
rect 20532 6244 20588 6246
rect 20636 6298 20692 6300
rect 20636 6246 20638 6298
rect 20638 6246 20690 6298
rect 20690 6246 20692 6298
rect 20636 6244 20692 6246
rect 20740 6298 20796 6300
rect 20740 6246 20742 6298
rect 20742 6246 20794 6298
rect 20794 6246 20796 6298
rect 20740 6244 20796 6246
rect 20412 6018 20468 6020
rect 20412 5966 20414 6018
rect 20414 5966 20466 6018
rect 20466 5966 20468 6018
rect 20412 5964 20468 5966
rect 20748 5628 20804 5684
rect 20532 4730 20588 4732
rect 20532 4678 20534 4730
rect 20534 4678 20586 4730
rect 20586 4678 20588 4730
rect 20532 4676 20588 4678
rect 20636 4730 20692 4732
rect 20636 4678 20638 4730
rect 20638 4678 20690 4730
rect 20690 4678 20692 4730
rect 20636 4676 20692 4678
rect 20740 4730 20796 4732
rect 20740 4678 20742 4730
rect 20742 4678 20794 4730
rect 20794 4678 20796 4730
rect 20740 4676 20796 4678
rect 20188 3612 20244 3668
rect 19628 3276 19684 3332
rect 19740 3500 19796 3556
rect 20300 3554 20356 3556
rect 20300 3502 20302 3554
rect 20302 3502 20354 3554
rect 20354 3502 20356 3554
rect 20300 3500 20356 3502
rect 21308 6748 21364 6804
rect 22988 12962 23044 12964
rect 22988 12910 22990 12962
rect 22990 12910 23042 12962
rect 23042 12910 23044 12962
rect 22988 12908 23044 12910
rect 22764 11394 22820 11396
rect 22764 11342 22766 11394
rect 22766 11342 22818 11394
rect 22818 11342 22820 11394
rect 22764 11340 22820 11342
rect 22876 11170 22932 11172
rect 22876 11118 22878 11170
rect 22878 11118 22930 11170
rect 22930 11118 22932 11170
rect 22876 11116 22932 11118
rect 22428 6972 22484 7028
rect 21644 6578 21700 6580
rect 21644 6526 21646 6578
rect 21646 6526 21698 6578
rect 21698 6526 21700 6578
rect 21644 6524 21700 6526
rect 22428 5682 22484 5684
rect 22428 5630 22430 5682
rect 22430 5630 22482 5682
rect 22482 5630 22484 5682
rect 22428 5628 22484 5630
rect 22652 10722 22708 10724
rect 22652 10670 22654 10722
rect 22654 10670 22706 10722
rect 22706 10670 22708 10722
rect 22652 10668 22708 10670
rect 22764 10444 22820 10500
rect 22876 10108 22932 10164
rect 21756 4508 21812 4564
rect 23212 12460 23268 12516
rect 23548 13522 23604 13524
rect 23548 13470 23550 13522
rect 23550 13470 23602 13522
rect 23602 13470 23604 13522
rect 23548 13468 23604 13470
rect 24220 14140 24276 14196
rect 23996 13858 24052 13860
rect 23996 13806 23998 13858
rect 23998 13806 24050 13858
rect 24050 13806 24052 13858
rect 23996 13804 24052 13806
rect 24108 13580 24164 13636
rect 23772 12738 23828 12740
rect 23772 12686 23774 12738
rect 23774 12686 23826 12738
rect 23826 12686 23828 12738
rect 23772 12684 23828 12686
rect 23660 12572 23716 12628
rect 23884 12236 23940 12292
rect 23660 11676 23716 11732
rect 23884 11564 23940 11620
rect 24444 16156 24500 16212
rect 24332 13132 24388 13188
rect 24556 15314 24612 15316
rect 24556 15262 24558 15314
rect 24558 15262 24610 15314
rect 24610 15262 24612 15314
rect 24556 15260 24612 15262
rect 25228 28140 25284 28196
rect 25004 27244 25060 27300
rect 25116 27186 25172 27188
rect 25116 27134 25118 27186
rect 25118 27134 25170 27186
rect 25170 27134 25172 27186
rect 25116 27132 25172 27134
rect 25004 25506 25060 25508
rect 25004 25454 25006 25506
rect 25006 25454 25058 25506
rect 25058 25454 25060 25506
rect 25004 25452 25060 25454
rect 25228 24220 25284 24276
rect 25004 21980 25060 22036
rect 25452 30156 25508 30212
rect 26460 31500 26516 31556
rect 26236 31052 26292 31108
rect 26012 30828 26068 30884
rect 26012 30156 26068 30212
rect 27356 31666 27412 31668
rect 27356 31614 27358 31666
rect 27358 31614 27410 31666
rect 27410 31614 27412 31666
rect 27356 31612 27412 31614
rect 27132 31554 27188 31556
rect 27132 31502 27134 31554
rect 27134 31502 27186 31554
rect 27186 31502 27188 31554
rect 27132 31500 27188 31502
rect 26684 30380 26740 30436
rect 26796 30044 26852 30100
rect 25564 28028 25620 28084
rect 25900 27692 25956 27748
rect 25900 27468 25956 27524
rect 25788 27132 25844 27188
rect 25564 26908 25620 26964
rect 26124 29538 26180 29540
rect 26124 29486 26126 29538
rect 26126 29486 26178 29538
rect 26178 29486 26180 29538
rect 26124 29484 26180 29486
rect 26460 29372 26516 29428
rect 26236 28700 26292 28756
rect 26460 28530 26516 28532
rect 26460 28478 26462 28530
rect 26462 28478 26514 28530
rect 26514 28478 26516 28530
rect 26460 28476 26516 28478
rect 26796 29484 26852 29540
rect 27132 29372 27188 29428
rect 26684 29260 26740 29316
rect 26572 28252 26628 28308
rect 26348 28028 26404 28084
rect 26908 28252 26964 28308
rect 26796 27746 26852 27748
rect 26796 27694 26798 27746
rect 26798 27694 26850 27746
rect 26850 27694 26852 27746
rect 26796 27692 26852 27694
rect 26684 27356 26740 27412
rect 26572 27244 26628 27300
rect 26796 27132 26852 27188
rect 29596 36988 29652 37044
rect 28812 36316 28868 36372
rect 28700 36258 28756 36260
rect 28700 36206 28702 36258
rect 28702 36206 28754 36258
rect 28754 36206 28756 36258
rect 28700 36204 28756 36206
rect 28924 36258 28980 36260
rect 28924 36206 28926 36258
rect 28926 36206 28978 36258
rect 28978 36206 28980 36258
rect 28924 36204 28980 36206
rect 29372 36204 29428 36260
rect 27804 34972 27860 35028
rect 27692 34636 27748 34692
rect 27692 30156 27748 30212
rect 28364 34636 28420 34692
rect 28700 35420 28756 35476
rect 29148 35420 29204 35476
rect 29260 35532 29316 35588
rect 29036 35308 29092 35364
rect 28364 34300 28420 34356
rect 28028 34018 28084 34020
rect 28028 33966 28030 34018
rect 28030 33966 28082 34018
rect 28082 33966 28084 34018
rect 28028 33964 28084 33966
rect 28252 33346 28308 33348
rect 28252 33294 28254 33346
rect 28254 33294 28306 33346
rect 28306 33294 28308 33346
rect 28252 33292 28308 33294
rect 28140 33180 28196 33236
rect 28588 34188 28644 34244
rect 28700 35196 28756 35252
rect 28924 34860 28980 34916
rect 28812 34748 28868 34804
rect 27916 31948 27972 32004
rect 28588 33404 28644 33460
rect 28588 31612 28644 31668
rect 28252 31388 28308 31444
rect 28140 30492 28196 30548
rect 28028 29314 28084 29316
rect 28028 29262 28030 29314
rect 28030 29262 28082 29314
rect 28082 29262 28084 29314
rect 28028 29260 28084 29262
rect 27580 28476 27636 28532
rect 27468 28252 27524 28308
rect 27132 28028 27188 28084
rect 27804 28082 27860 28084
rect 27804 28030 27806 28082
rect 27806 28030 27858 28082
rect 27858 28030 27860 28082
rect 27804 28028 27860 28030
rect 27020 27692 27076 27748
rect 27132 27580 27188 27636
rect 27020 27074 27076 27076
rect 27020 27022 27022 27074
rect 27022 27022 27074 27074
rect 27074 27022 27076 27074
rect 27020 27020 27076 27022
rect 27356 27132 27412 27188
rect 27468 27020 27524 27076
rect 26236 26402 26292 26404
rect 26236 26350 26238 26402
rect 26238 26350 26290 26402
rect 26290 26350 26292 26402
rect 26236 26348 26292 26350
rect 25900 25340 25956 25396
rect 26012 24220 26068 24276
rect 25452 23548 25508 23604
rect 25228 20972 25284 21028
rect 24892 19404 24948 19460
rect 25004 20524 25060 20580
rect 25228 19852 25284 19908
rect 25228 19010 25284 19012
rect 25228 18958 25230 19010
rect 25230 18958 25282 19010
rect 25282 18958 25284 19010
rect 25228 18956 25284 18958
rect 25004 17836 25060 17892
rect 25340 17106 25396 17108
rect 25340 17054 25342 17106
rect 25342 17054 25394 17106
rect 25394 17054 25396 17106
rect 25340 17052 25396 17054
rect 25004 16380 25060 16436
rect 24780 14924 24836 14980
rect 24892 13804 24948 13860
rect 24220 12850 24276 12852
rect 24220 12798 24222 12850
rect 24222 12798 24274 12850
rect 24274 12798 24276 12850
rect 24220 12796 24276 12798
rect 25340 15314 25396 15316
rect 25340 15262 25342 15314
rect 25342 15262 25394 15314
rect 25394 15262 25396 15314
rect 25340 15260 25396 15262
rect 25676 23548 25732 23604
rect 25564 23436 25620 23492
rect 25676 23154 25732 23156
rect 25676 23102 25678 23154
rect 25678 23102 25730 23154
rect 25730 23102 25732 23154
rect 25676 23100 25732 23102
rect 26348 25564 26404 25620
rect 26348 23826 26404 23828
rect 26348 23774 26350 23826
rect 26350 23774 26402 23826
rect 26402 23774 26404 23826
rect 26348 23772 26404 23774
rect 26124 23436 26180 23492
rect 26684 26236 26740 26292
rect 26908 25564 26964 25620
rect 26908 25394 26964 25396
rect 26908 25342 26910 25394
rect 26910 25342 26962 25394
rect 26962 25342 26964 25394
rect 26908 25340 26964 25342
rect 26684 23436 26740 23492
rect 26460 23324 26516 23380
rect 28588 30994 28644 30996
rect 28588 30942 28590 30994
rect 28590 30942 28642 30994
rect 28642 30942 28644 30994
rect 28588 30940 28644 30942
rect 28252 30210 28308 30212
rect 28252 30158 28254 30210
rect 28254 30158 28306 30210
rect 28306 30158 28308 30210
rect 28252 30156 28308 30158
rect 28364 29932 28420 29988
rect 28028 28082 28084 28084
rect 28028 28030 28030 28082
rect 28030 28030 28082 28082
rect 28082 28030 28084 28082
rect 28028 28028 28084 28030
rect 27132 26290 27188 26292
rect 27132 26238 27134 26290
rect 27134 26238 27186 26290
rect 27186 26238 27188 26290
rect 27132 26236 27188 26238
rect 27692 26348 27748 26404
rect 27468 25506 27524 25508
rect 27468 25454 27470 25506
rect 27470 25454 27522 25506
rect 27522 25454 27524 25506
rect 27468 25452 27524 25454
rect 27244 25116 27300 25172
rect 26012 23042 26068 23044
rect 26012 22990 26014 23042
rect 26014 22990 26066 23042
rect 26066 22990 26068 23042
rect 26012 22988 26068 22990
rect 26348 22594 26404 22596
rect 26348 22542 26350 22594
rect 26350 22542 26402 22594
rect 26402 22542 26404 22594
rect 26348 22540 26404 22542
rect 25788 22428 25844 22484
rect 26572 22428 26628 22484
rect 25676 21868 25732 21924
rect 26012 22146 26068 22148
rect 26012 22094 26014 22146
rect 26014 22094 26066 22146
rect 26066 22094 26068 22146
rect 26012 22092 26068 22094
rect 25900 21756 25956 21812
rect 25564 21474 25620 21476
rect 25564 21422 25566 21474
rect 25566 21422 25618 21474
rect 25618 21422 25620 21474
rect 25564 21420 25620 21422
rect 25788 21420 25844 21476
rect 26124 21586 26180 21588
rect 26124 21534 26126 21586
rect 26126 21534 26178 21586
rect 26178 21534 26180 21586
rect 26124 21532 26180 21534
rect 26572 22204 26628 22260
rect 26460 21586 26516 21588
rect 26460 21534 26462 21586
rect 26462 21534 26514 21586
rect 26514 21534 26516 21586
rect 26460 21532 26516 21534
rect 26236 20748 26292 20804
rect 25900 20524 25956 20580
rect 26796 21868 26852 21924
rect 27244 23548 27300 23604
rect 27468 24780 27524 24836
rect 27244 23378 27300 23380
rect 27244 23326 27246 23378
rect 27246 23326 27298 23378
rect 27298 23326 27300 23378
rect 27244 23324 27300 23326
rect 27020 21756 27076 21812
rect 27244 21756 27300 21812
rect 26908 20076 26964 20132
rect 27580 21756 27636 21812
rect 27804 26236 27860 26292
rect 28140 27858 28196 27860
rect 28140 27806 28142 27858
rect 28142 27806 28194 27858
rect 28194 27806 28196 27858
rect 28140 27804 28196 27806
rect 28364 28140 28420 28196
rect 28588 29314 28644 29316
rect 28588 29262 28590 29314
rect 28590 29262 28642 29314
rect 28642 29262 28644 29314
rect 28588 29260 28644 29262
rect 28700 28082 28756 28084
rect 28700 28030 28702 28082
rect 28702 28030 28754 28082
rect 28754 28030 28756 28082
rect 28700 28028 28756 28030
rect 28252 26348 28308 26404
rect 28028 25900 28084 25956
rect 28588 26684 28644 26740
rect 28588 25788 28644 25844
rect 28700 25900 28756 25956
rect 28140 25228 28196 25284
rect 27804 24780 27860 24836
rect 28476 25452 28532 25508
rect 27916 24722 27972 24724
rect 27916 24670 27918 24722
rect 27918 24670 27970 24722
rect 27970 24670 27972 24722
rect 27916 24668 27972 24670
rect 28140 24834 28196 24836
rect 28140 24782 28142 24834
rect 28142 24782 28194 24834
rect 28194 24782 28196 24834
rect 28140 24780 28196 24782
rect 28588 24668 28644 24724
rect 28700 25228 28756 25284
rect 28476 23884 28532 23940
rect 27916 23436 27972 23492
rect 27804 22764 27860 22820
rect 27804 22428 27860 22484
rect 28028 22764 28084 22820
rect 28364 23548 28420 23604
rect 28364 23266 28420 23268
rect 28364 23214 28366 23266
rect 28366 23214 28418 23266
rect 28418 23214 28420 23266
rect 28364 23212 28420 23214
rect 28252 23100 28308 23156
rect 28140 22092 28196 22148
rect 27804 21532 27860 21588
rect 29484 35868 29540 35924
rect 29484 35698 29540 35700
rect 29484 35646 29486 35698
rect 29486 35646 29538 35698
rect 29538 35646 29540 35698
rect 29484 35644 29540 35646
rect 30192 36874 30248 36876
rect 30192 36822 30194 36874
rect 30194 36822 30246 36874
rect 30246 36822 30248 36874
rect 30192 36820 30248 36822
rect 30296 36874 30352 36876
rect 30296 36822 30298 36874
rect 30298 36822 30350 36874
rect 30350 36822 30352 36874
rect 30296 36820 30352 36822
rect 30400 36874 30456 36876
rect 30400 36822 30402 36874
rect 30402 36822 30454 36874
rect 30454 36822 30456 36874
rect 30400 36820 30456 36822
rect 31164 36594 31220 36596
rect 31164 36542 31166 36594
rect 31166 36542 31218 36594
rect 31218 36542 31220 36594
rect 31164 36540 31220 36542
rect 34972 37212 35028 37268
rect 31612 36594 31668 36596
rect 31612 36542 31614 36594
rect 31614 36542 31666 36594
rect 31666 36542 31668 36594
rect 31612 36540 31668 36542
rect 32844 36540 32900 36596
rect 29820 36370 29876 36372
rect 29820 36318 29822 36370
rect 29822 36318 29874 36370
rect 29874 36318 29876 36370
rect 29820 36316 29876 36318
rect 30156 35532 30212 35588
rect 29596 35420 29652 35476
rect 29372 35308 29428 35364
rect 29484 34914 29540 34916
rect 29484 34862 29486 34914
rect 29486 34862 29538 34914
rect 29538 34862 29540 34914
rect 29484 34860 29540 34862
rect 29708 34802 29764 34804
rect 29708 34750 29710 34802
rect 29710 34750 29762 34802
rect 29762 34750 29764 34802
rect 29708 34748 29764 34750
rect 30492 35474 30548 35476
rect 30492 35422 30494 35474
rect 30494 35422 30546 35474
rect 30546 35422 30548 35474
rect 30492 35420 30548 35422
rect 30192 35306 30248 35308
rect 30192 35254 30194 35306
rect 30194 35254 30246 35306
rect 30246 35254 30248 35306
rect 30192 35252 30248 35254
rect 30296 35306 30352 35308
rect 30296 35254 30298 35306
rect 30298 35254 30350 35306
rect 30350 35254 30352 35306
rect 30296 35252 30352 35254
rect 30400 35306 30456 35308
rect 30400 35254 30402 35306
rect 30402 35254 30454 35306
rect 30454 35254 30456 35306
rect 30400 35252 30456 35254
rect 29820 34524 29876 34580
rect 30604 34860 30660 34916
rect 31276 35698 31332 35700
rect 31276 35646 31278 35698
rect 31278 35646 31330 35698
rect 31330 35646 31332 35698
rect 31276 35644 31332 35646
rect 31948 35586 32004 35588
rect 31948 35534 31950 35586
rect 31950 35534 32002 35586
rect 32002 35534 32004 35586
rect 31948 35532 32004 35534
rect 30828 34748 30884 34804
rect 30716 34524 30772 34580
rect 30044 34300 30100 34356
rect 29932 34188 29988 34244
rect 29260 33234 29316 33236
rect 29260 33182 29262 33234
rect 29262 33182 29314 33234
rect 29314 33182 29316 33234
rect 29260 33180 29316 33182
rect 29484 31948 29540 32004
rect 29820 33122 29876 33124
rect 29820 33070 29822 33122
rect 29822 33070 29874 33122
rect 29874 33070 29876 33122
rect 29820 33068 29876 33070
rect 30192 33738 30248 33740
rect 30192 33686 30194 33738
rect 30194 33686 30246 33738
rect 30246 33686 30248 33738
rect 30192 33684 30248 33686
rect 30296 33738 30352 33740
rect 30296 33686 30298 33738
rect 30298 33686 30350 33738
rect 30350 33686 30352 33738
rect 30296 33684 30352 33686
rect 30400 33738 30456 33740
rect 30400 33686 30402 33738
rect 30402 33686 30454 33738
rect 30454 33686 30456 33738
rect 30400 33684 30456 33686
rect 30380 33346 30436 33348
rect 30380 33294 30382 33346
rect 30382 33294 30434 33346
rect 30434 33294 30436 33346
rect 30380 33292 30436 33294
rect 30828 32562 30884 32564
rect 30828 32510 30830 32562
rect 30830 32510 30882 32562
rect 30882 32510 30884 32562
rect 30828 32508 30884 32510
rect 30192 32170 30248 32172
rect 30192 32118 30194 32170
rect 30194 32118 30246 32170
rect 30246 32118 30248 32170
rect 30192 32116 30248 32118
rect 30296 32170 30352 32172
rect 30296 32118 30298 32170
rect 30298 32118 30350 32170
rect 30350 32118 30352 32170
rect 30296 32116 30352 32118
rect 30400 32170 30456 32172
rect 30400 32118 30402 32170
rect 30402 32118 30454 32170
rect 30454 32118 30456 32170
rect 30400 32116 30456 32118
rect 30156 31778 30212 31780
rect 30156 31726 30158 31778
rect 30158 31726 30210 31778
rect 30210 31726 30212 31778
rect 30156 31724 30212 31726
rect 30604 31948 30660 32004
rect 30380 31666 30436 31668
rect 30380 31614 30382 31666
rect 30382 31614 30434 31666
rect 30434 31614 30436 31666
rect 30380 31612 30436 31614
rect 29596 31500 29652 31556
rect 30492 31500 30548 31556
rect 30156 31106 30212 31108
rect 30156 31054 30158 31106
rect 30158 31054 30210 31106
rect 30210 31054 30212 31106
rect 30156 31052 30212 31054
rect 28924 28028 28980 28084
rect 29148 30156 29204 30212
rect 29036 27858 29092 27860
rect 29036 27806 29038 27858
rect 29038 27806 29090 27858
rect 29090 27806 29092 27858
rect 29036 27804 29092 27806
rect 28924 25228 28980 25284
rect 28924 25004 28980 25060
rect 29036 24892 29092 24948
rect 29036 24722 29092 24724
rect 29036 24670 29038 24722
rect 29038 24670 29090 24722
rect 29090 24670 29092 24722
rect 29036 24668 29092 24670
rect 28924 24498 28980 24500
rect 28924 24446 28926 24498
rect 28926 24446 28978 24498
rect 28978 24446 28980 24498
rect 28924 24444 28980 24446
rect 28812 22988 28868 23044
rect 29372 30156 29428 30212
rect 29260 29986 29316 29988
rect 29260 29934 29262 29986
rect 29262 29934 29314 29986
rect 29314 29934 29316 29986
rect 29260 29932 29316 29934
rect 29372 29596 29428 29652
rect 29596 30268 29652 30324
rect 31164 33234 31220 33236
rect 31164 33182 31166 33234
rect 31166 33182 31218 33234
rect 31218 33182 31220 33234
rect 31164 33180 31220 33182
rect 31500 34524 31556 34580
rect 31948 34300 32004 34356
rect 32172 35420 32228 35476
rect 31500 34076 31556 34132
rect 32060 34130 32116 34132
rect 32060 34078 32062 34130
rect 32062 34078 32114 34130
rect 32114 34078 32116 34130
rect 32060 34076 32116 34078
rect 31948 34018 32004 34020
rect 31948 33966 31950 34018
rect 31950 33966 32002 34018
rect 32002 33966 32004 34018
rect 31948 33964 32004 33966
rect 31388 33458 31444 33460
rect 31388 33406 31390 33458
rect 31390 33406 31442 33458
rect 31442 33406 31444 33458
rect 31388 33404 31444 33406
rect 31836 33404 31892 33460
rect 32060 33234 32116 33236
rect 32060 33182 32062 33234
rect 32062 33182 32114 33234
rect 32114 33182 32116 33234
rect 32060 33180 32116 33182
rect 31388 32060 31444 32116
rect 31836 32396 31892 32452
rect 31836 31948 31892 32004
rect 31388 31890 31444 31892
rect 31388 31838 31390 31890
rect 31390 31838 31442 31890
rect 31442 31838 31444 31890
rect 31388 31836 31444 31838
rect 31500 31778 31556 31780
rect 31500 31726 31502 31778
rect 31502 31726 31554 31778
rect 31554 31726 31556 31778
rect 31500 31724 31556 31726
rect 31052 31500 31108 31556
rect 31388 31612 31444 31668
rect 30940 31388 30996 31444
rect 31276 31276 31332 31332
rect 30192 30602 30248 30604
rect 30192 30550 30194 30602
rect 30194 30550 30246 30602
rect 30246 30550 30248 30602
rect 30192 30548 30248 30550
rect 30296 30602 30352 30604
rect 30296 30550 30298 30602
rect 30298 30550 30350 30602
rect 30350 30550 30352 30602
rect 30296 30548 30352 30550
rect 30400 30602 30456 30604
rect 30400 30550 30402 30602
rect 30402 30550 30454 30602
rect 30454 30550 30456 30602
rect 30400 30548 30456 30550
rect 30716 30604 30772 30660
rect 29932 30156 29988 30212
rect 29708 30098 29764 30100
rect 29708 30046 29710 30098
rect 29710 30046 29762 30098
rect 29762 30046 29764 30098
rect 29708 30044 29764 30046
rect 29708 29484 29764 29540
rect 29932 29650 29988 29652
rect 29932 29598 29934 29650
rect 29934 29598 29986 29650
rect 29986 29598 29988 29650
rect 29932 29596 29988 29598
rect 30156 29650 30212 29652
rect 30156 29598 30158 29650
rect 30158 29598 30210 29650
rect 30210 29598 30212 29650
rect 30156 29596 30212 29598
rect 30044 29484 30100 29540
rect 30192 29034 30248 29036
rect 30192 28982 30194 29034
rect 30194 28982 30246 29034
rect 30246 28982 30248 29034
rect 30192 28980 30248 28982
rect 30296 29034 30352 29036
rect 30296 28982 30298 29034
rect 30298 28982 30350 29034
rect 30350 28982 30352 29034
rect 30296 28980 30352 28982
rect 30400 29034 30456 29036
rect 30400 28982 30402 29034
rect 30402 28982 30454 29034
rect 30454 28982 30456 29034
rect 30400 28980 30456 28982
rect 30380 28812 30436 28868
rect 30492 27858 30548 27860
rect 30492 27806 30494 27858
rect 30494 27806 30546 27858
rect 30546 27806 30548 27858
rect 30492 27804 30548 27806
rect 30828 29708 30884 29764
rect 31052 29596 31108 29652
rect 30940 28530 30996 28532
rect 30940 28478 30942 28530
rect 30942 28478 30994 28530
rect 30994 28478 30996 28530
rect 30940 28476 30996 28478
rect 31164 28252 31220 28308
rect 30716 27916 30772 27972
rect 30492 27580 30548 27636
rect 30828 27634 30884 27636
rect 30828 27582 30830 27634
rect 30830 27582 30882 27634
rect 30882 27582 30884 27634
rect 30828 27580 30884 27582
rect 30192 27466 30248 27468
rect 30192 27414 30194 27466
rect 30194 27414 30246 27466
rect 30246 27414 30248 27466
rect 30192 27412 30248 27414
rect 30296 27466 30352 27468
rect 30296 27414 30298 27466
rect 30298 27414 30350 27466
rect 30350 27414 30352 27466
rect 30296 27412 30352 27414
rect 30400 27466 30456 27468
rect 30400 27414 30402 27466
rect 30402 27414 30454 27466
rect 30454 27414 30456 27466
rect 30400 27412 30456 27414
rect 31164 27244 31220 27300
rect 29820 27020 29876 27076
rect 30380 26962 30436 26964
rect 30380 26910 30382 26962
rect 30382 26910 30434 26962
rect 30434 26910 30436 26962
rect 30380 26908 30436 26910
rect 29708 26572 29764 26628
rect 30716 26348 30772 26404
rect 29372 26290 29428 26292
rect 29372 26238 29374 26290
rect 29374 26238 29426 26290
rect 29426 26238 29428 26290
rect 29372 26236 29428 26238
rect 29260 25564 29316 25620
rect 29596 25340 29652 25396
rect 30192 25898 30248 25900
rect 30192 25846 30194 25898
rect 30194 25846 30246 25898
rect 30246 25846 30248 25898
rect 30192 25844 30248 25846
rect 30296 25898 30352 25900
rect 30296 25846 30298 25898
rect 30298 25846 30350 25898
rect 30350 25846 30352 25898
rect 30296 25844 30352 25846
rect 30400 25898 30456 25900
rect 30400 25846 30402 25898
rect 30402 25846 30454 25898
rect 30454 25846 30456 25898
rect 30400 25844 30456 25846
rect 30268 25618 30324 25620
rect 30268 25566 30270 25618
rect 30270 25566 30322 25618
rect 30322 25566 30324 25618
rect 30268 25564 30324 25566
rect 29820 25340 29876 25396
rect 29596 24892 29652 24948
rect 29708 25228 29764 25284
rect 29932 25004 29988 25060
rect 30156 25228 30212 25284
rect 30044 24892 30100 24948
rect 29372 24668 29428 24724
rect 29820 24050 29876 24052
rect 29820 23998 29822 24050
rect 29822 23998 29874 24050
rect 29874 23998 29876 24050
rect 29820 23996 29876 23998
rect 29708 23938 29764 23940
rect 29708 23886 29710 23938
rect 29710 23886 29762 23938
rect 29762 23886 29764 23938
rect 29708 23884 29764 23886
rect 29260 23212 29316 23268
rect 29036 22876 29092 22932
rect 29148 22764 29204 22820
rect 28364 21868 28420 21924
rect 27356 20524 27412 20580
rect 27132 20018 27188 20020
rect 27132 19966 27134 20018
rect 27134 19966 27186 20018
rect 27186 19966 27188 20018
rect 27132 19964 27188 19966
rect 27468 19964 27524 20020
rect 27244 19740 27300 19796
rect 26236 19404 26292 19460
rect 26124 19234 26180 19236
rect 26124 19182 26126 19234
rect 26126 19182 26178 19234
rect 26178 19182 26180 19234
rect 26124 19180 26180 19182
rect 25676 19010 25732 19012
rect 25676 18958 25678 19010
rect 25678 18958 25730 19010
rect 25730 18958 25732 19010
rect 25676 18956 25732 18958
rect 26124 18620 26180 18676
rect 25676 17836 25732 17892
rect 25564 17442 25620 17444
rect 25564 17390 25566 17442
rect 25566 17390 25618 17442
rect 25618 17390 25620 17442
rect 25564 17388 25620 17390
rect 25676 17164 25732 17220
rect 25564 16380 25620 16436
rect 25788 16994 25844 16996
rect 25788 16942 25790 16994
rect 25790 16942 25842 16994
rect 25842 16942 25844 16994
rect 25788 16940 25844 16942
rect 25788 15932 25844 15988
rect 25788 15314 25844 15316
rect 25788 15262 25790 15314
rect 25790 15262 25842 15314
rect 25842 15262 25844 15314
rect 25788 15260 25844 15262
rect 25564 13804 25620 13860
rect 25004 13244 25060 13300
rect 25228 13692 25284 13748
rect 24892 13020 24948 13076
rect 25116 13074 25172 13076
rect 25116 13022 25118 13074
rect 25118 13022 25170 13074
rect 25170 13022 25172 13074
rect 25116 13020 25172 13022
rect 25452 13692 25508 13748
rect 25340 13634 25396 13636
rect 25340 13582 25342 13634
rect 25342 13582 25394 13634
rect 25394 13582 25396 13634
rect 25340 13580 25396 13582
rect 25452 13356 25508 13412
rect 25228 12962 25284 12964
rect 25228 12910 25230 12962
rect 25230 12910 25282 12962
rect 25282 12910 25284 12962
rect 25228 12908 25284 12910
rect 25340 13244 25396 13300
rect 23436 11340 23492 11396
rect 23548 10892 23604 10948
rect 23660 11228 23716 11284
rect 23660 10668 23716 10724
rect 24108 12738 24164 12740
rect 24108 12686 24110 12738
rect 24110 12686 24162 12738
rect 24162 12686 24164 12738
rect 24108 12684 24164 12686
rect 24444 12684 24500 12740
rect 24108 11900 24164 11956
rect 24332 12178 24388 12180
rect 24332 12126 24334 12178
rect 24334 12126 24386 12178
rect 24386 12126 24388 12178
rect 24332 12124 24388 12126
rect 25452 12738 25508 12740
rect 25452 12686 25454 12738
rect 25454 12686 25506 12738
rect 25506 12686 25508 12738
rect 25452 12684 25508 12686
rect 24780 12572 24836 12628
rect 24668 12460 24724 12516
rect 24220 11676 24276 11732
rect 23996 11340 24052 11396
rect 24108 11282 24164 11284
rect 24108 11230 24110 11282
rect 24110 11230 24162 11282
rect 24162 11230 24164 11282
rect 24108 11228 24164 11230
rect 23996 10892 24052 10948
rect 24220 11116 24276 11172
rect 24444 11564 24500 11620
rect 24556 11282 24612 11284
rect 24556 11230 24558 11282
rect 24558 11230 24610 11282
rect 24610 11230 24612 11282
rect 24556 11228 24612 11230
rect 24108 10610 24164 10612
rect 24108 10558 24110 10610
rect 24110 10558 24162 10610
rect 24162 10558 24164 10610
rect 24556 10780 24612 10836
rect 25900 14140 25956 14196
rect 25788 13916 25844 13972
rect 26012 13804 26068 13860
rect 27020 19404 27076 19460
rect 26572 19234 26628 19236
rect 26572 19182 26574 19234
rect 26574 19182 26626 19234
rect 26626 19182 26628 19234
rect 26572 19180 26628 19182
rect 27132 19180 27188 19236
rect 27356 19234 27412 19236
rect 27356 19182 27358 19234
rect 27358 19182 27410 19234
rect 27410 19182 27412 19234
rect 27356 19180 27412 19182
rect 27244 18732 27300 18788
rect 28140 20690 28196 20692
rect 28140 20638 28142 20690
rect 28142 20638 28194 20690
rect 28194 20638 28196 20690
rect 28140 20636 28196 20638
rect 27916 20076 27972 20132
rect 27804 20018 27860 20020
rect 27804 19966 27806 20018
rect 27806 19966 27858 20018
rect 27858 19966 27860 20018
rect 27804 19964 27860 19966
rect 27916 19180 27972 19236
rect 28140 19852 28196 19908
rect 28028 19068 28084 19124
rect 28028 18844 28084 18900
rect 26796 17554 26852 17556
rect 26796 17502 26798 17554
rect 26798 17502 26850 17554
rect 26850 17502 26852 17554
rect 26796 17500 26852 17502
rect 26684 16882 26740 16884
rect 26684 16830 26686 16882
rect 26686 16830 26738 16882
rect 26738 16830 26740 16882
rect 26684 16828 26740 16830
rect 27132 17052 27188 17108
rect 27692 18172 27748 18228
rect 28588 21474 28644 21476
rect 28588 21422 28590 21474
rect 28590 21422 28642 21474
rect 28642 21422 28644 21474
rect 28588 21420 28644 21422
rect 28700 20412 28756 20468
rect 28588 19404 28644 19460
rect 28588 19180 28644 19236
rect 29596 21810 29652 21812
rect 29596 21758 29598 21810
rect 29598 21758 29650 21810
rect 29650 21758 29652 21810
rect 29596 21756 29652 21758
rect 29372 21532 29428 21588
rect 29148 21420 29204 21476
rect 29596 21532 29652 21588
rect 29932 22092 29988 22148
rect 29932 21810 29988 21812
rect 29932 21758 29934 21810
rect 29934 21758 29986 21810
rect 29986 21758 29988 21810
rect 29932 21756 29988 21758
rect 29596 21308 29652 21364
rect 29820 21532 29876 21588
rect 29260 20524 29316 20580
rect 29036 19852 29092 19908
rect 29372 19964 29428 20020
rect 29036 19234 29092 19236
rect 29036 19182 29038 19234
rect 29038 19182 29090 19234
rect 29090 19182 29092 19234
rect 29036 19180 29092 19182
rect 29820 20748 29876 20804
rect 29708 20412 29764 20468
rect 29820 20188 29876 20244
rect 29708 19234 29764 19236
rect 29708 19182 29710 19234
rect 29710 19182 29762 19234
rect 29762 19182 29764 19234
rect 29708 19180 29764 19182
rect 29708 18956 29764 19012
rect 28252 18396 28308 18452
rect 29036 18450 29092 18452
rect 29036 18398 29038 18450
rect 29038 18398 29090 18450
rect 29090 18398 29092 18450
rect 29036 18396 29092 18398
rect 29484 18338 29540 18340
rect 29484 18286 29486 18338
rect 29486 18286 29538 18338
rect 29538 18286 29540 18338
rect 29484 18284 29540 18286
rect 29484 18060 29540 18116
rect 27692 16940 27748 16996
rect 27804 17276 27860 17332
rect 26348 16156 26404 16212
rect 26348 15036 26404 15092
rect 26124 13580 26180 13636
rect 26236 13692 26292 13748
rect 26012 13244 26068 13300
rect 26236 13020 26292 13076
rect 27020 15986 27076 15988
rect 27020 15934 27022 15986
rect 27022 15934 27074 15986
rect 27074 15934 27076 15986
rect 27020 15932 27076 15934
rect 27468 15986 27524 15988
rect 27468 15934 27470 15986
rect 27470 15934 27522 15986
rect 27522 15934 27524 15986
rect 27468 15932 27524 15934
rect 27132 15260 27188 15316
rect 27132 14252 27188 14308
rect 26460 13580 26516 13636
rect 26684 13634 26740 13636
rect 26684 13582 26686 13634
rect 26686 13582 26738 13634
rect 26738 13582 26740 13634
rect 26684 13580 26740 13582
rect 26908 13522 26964 13524
rect 26908 13470 26910 13522
rect 26910 13470 26962 13522
rect 26962 13470 26964 13522
rect 26908 13468 26964 13470
rect 26460 13020 26516 13076
rect 25676 12178 25732 12180
rect 25676 12126 25678 12178
rect 25678 12126 25730 12178
rect 25730 12126 25732 12178
rect 25676 12124 25732 12126
rect 25452 12012 25508 12068
rect 25340 11564 25396 11620
rect 24892 11340 24948 11396
rect 24108 10556 24164 10558
rect 23996 10332 24052 10388
rect 23772 10220 23828 10276
rect 23324 10108 23380 10164
rect 24108 10108 24164 10164
rect 23884 8092 23940 8148
rect 24892 10108 24948 10164
rect 25116 9996 25172 10052
rect 25676 11900 25732 11956
rect 25564 11452 25620 11508
rect 25452 10892 25508 10948
rect 25340 10332 25396 10388
rect 25788 11452 25844 11508
rect 25788 11228 25844 11284
rect 25788 10892 25844 10948
rect 25564 10108 25620 10164
rect 25788 10220 25844 10276
rect 24668 8092 24724 8148
rect 24220 7644 24276 7700
rect 23996 7586 24052 7588
rect 23996 7534 23998 7586
rect 23998 7534 24050 7586
rect 24050 7534 24052 7586
rect 23996 7532 24052 7534
rect 23212 4956 23268 5012
rect 23548 5740 23604 5796
rect 24220 5794 24276 5796
rect 24220 5742 24222 5794
rect 24222 5742 24274 5794
rect 24274 5742 24276 5794
rect 24220 5740 24276 5742
rect 25004 7644 25060 7700
rect 25340 7980 25396 8036
rect 26236 12012 26292 12068
rect 26124 11900 26180 11956
rect 26124 8204 26180 8260
rect 26012 8034 26068 8036
rect 26012 7982 26014 8034
rect 26014 7982 26066 8034
rect 26066 7982 26068 8034
rect 26012 7980 26068 7982
rect 25900 7868 25956 7924
rect 25340 7698 25396 7700
rect 25340 7646 25342 7698
rect 25342 7646 25394 7698
rect 25394 7646 25396 7698
rect 25340 7644 25396 7646
rect 26124 7644 26180 7700
rect 25900 7586 25956 7588
rect 25900 7534 25902 7586
rect 25902 7534 25954 7586
rect 25954 7534 25956 7586
rect 25900 7532 25956 7534
rect 25340 6466 25396 6468
rect 25340 6414 25342 6466
rect 25342 6414 25394 6466
rect 25394 6414 25396 6466
rect 25340 6412 25396 6414
rect 25116 6076 25172 6132
rect 25676 6076 25732 6132
rect 25004 5740 25060 5796
rect 23548 4620 23604 4676
rect 23324 4562 23380 4564
rect 23324 4510 23326 4562
rect 23326 4510 23378 4562
rect 23378 4510 23380 4562
rect 23324 4508 23380 4510
rect 24556 4956 24612 5012
rect 24444 4620 24500 4676
rect 23884 4284 23940 4340
rect 20972 3554 21028 3556
rect 20972 3502 20974 3554
rect 20974 3502 21026 3554
rect 21026 3502 21028 3554
rect 20972 3500 21028 3502
rect 20532 3162 20588 3164
rect 20532 3110 20534 3162
rect 20534 3110 20586 3162
rect 20586 3110 20588 3162
rect 20532 3108 20588 3110
rect 20636 3162 20692 3164
rect 20636 3110 20638 3162
rect 20638 3110 20690 3162
rect 20690 3110 20692 3162
rect 20636 3108 20692 3110
rect 20740 3162 20796 3164
rect 20740 3110 20742 3162
rect 20742 3110 20794 3162
rect 20794 3110 20796 3162
rect 20740 3108 20796 3110
rect 26012 6130 26068 6132
rect 26012 6078 26014 6130
rect 26014 6078 26066 6130
rect 26066 6078 26068 6130
rect 26012 6076 26068 6078
rect 26348 11170 26404 11172
rect 26348 11118 26350 11170
rect 26350 11118 26402 11170
rect 26402 11118 26404 11170
rect 26348 11116 26404 11118
rect 26796 13132 26852 13188
rect 27356 15260 27412 15316
rect 27356 13132 27412 13188
rect 28028 17164 28084 17220
rect 28812 17106 28868 17108
rect 28812 17054 28814 17106
rect 28814 17054 28866 17106
rect 28866 17054 28868 17106
rect 28812 17052 28868 17054
rect 28252 16940 28308 16996
rect 29260 16828 29316 16884
rect 29372 17724 29428 17780
rect 28476 16604 28532 16660
rect 28476 15820 28532 15876
rect 28140 15148 28196 15204
rect 28364 15260 28420 15316
rect 27804 13634 27860 13636
rect 27804 13582 27806 13634
rect 27806 13582 27858 13634
rect 27858 13582 27860 13634
rect 27804 13580 27860 13582
rect 27580 13074 27636 13076
rect 27580 13022 27582 13074
rect 27582 13022 27634 13074
rect 27634 13022 27636 13074
rect 27580 13020 27636 13022
rect 27468 12908 27524 12964
rect 26572 11788 26628 11844
rect 26796 12012 26852 12068
rect 28588 14700 28644 14756
rect 29932 19852 29988 19908
rect 30192 24330 30248 24332
rect 30192 24278 30194 24330
rect 30194 24278 30246 24330
rect 30246 24278 30248 24330
rect 30192 24276 30248 24278
rect 30296 24330 30352 24332
rect 30296 24278 30298 24330
rect 30298 24278 30350 24330
rect 30350 24278 30352 24330
rect 30296 24276 30352 24278
rect 30400 24330 30456 24332
rect 30400 24278 30402 24330
rect 30402 24278 30454 24330
rect 30454 24278 30456 24330
rect 30400 24276 30456 24278
rect 30492 23884 30548 23940
rect 30604 23826 30660 23828
rect 30604 23774 30606 23826
rect 30606 23774 30658 23826
rect 30658 23774 30660 23826
rect 30604 23772 30660 23774
rect 30380 23266 30436 23268
rect 30380 23214 30382 23266
rect 30382 23214 30434 23266
rect 30434 23214 30436 23266
rect 30380 23212 30436 23214
rect 30716 23154 30772 23156
rect 30716 23102 30718 23154
rect 30718 23102 30770 23154
rect 30770 23102 30772 23154
rect 30716 23100 30772 23102
rect 30192 22762 30248 22764
rect 30192 22710 30194 22762
rect 30194 22710 30246 22762
rect 30246 22710 30248 22762
rect 30192 22708 30248 22710
rect 30296 22762 30352 22764
rect 30296 22710 30298 22762
rect 30298 22710 30350 22762
rect 30350 22710 30352 22762
rect 30296 22708 30352 22710
rect 30400 22762 30456 22764
rect 30400 22710 30402 22762
rect 30402 22710 30454 22762
rect 30454 22710 30456 22762
rect 30400 22708 30456 22710
rect 31164 26402 31220 26404
rect 31164 26350 31166 26402
rect 31166 26350 31218 26402
rect 31218 26350 31220 26402
rect 31164 26348 31220 26350
rect 31276 26962 31332 26964
rect 31276 26910 31278 26962
rect 31278 26910 31330 26962
rect 31330 26910 31332 26962
rect 31276 26908 31332 26910
rect 31052 25452 31108 25508
rect 30940 23996 30996 24052
rect 33068 35308 33124 35364
rect 32396 33964 32452 34020
rect 32508 33740 32564 33796
rect 32396 33068 32452 33124
rect 32284 31948 32340 32004
rect 32172 31778 32228 31780
rect 32172 31726 32174 31778
rect 32174 31726 32226 31778
rect 32226 31726 32228 31778
rect 32172 31724 32228 31726
rect 31612 31052 31668 31108
rect 31724 30210 31780 30212
rect 31724 30158 31726 30210
rect 31726 30158 31778 30210
rect 31778 30158 31780 30210
rect 31724 30156 31780 30158
rect 32284 31612 32340 31668
rect 31500 29372 31556 29428
rect 31500 28812 31556 28868
rect 31612 28588 31668 28644
rect 32172 29372 32228 29428
rect 32396 31500 32452 31556
rect 33292 35698 33348 35700
rect 33292 35646 33294 35698
rect 33294 35646 33346 35698
rect 33346 35646 33348 35698
rect 33292 35644 33348 35646
rect 33516 35474 33572 35476
rect 33516 35422 33518 35474
rect 33518 35422 33570 35474
rect 33570 35422 33572 35474
rect 33516 35420 33572 35422
rect 33628 35308 33684 35364
rect 33292 34354 33348 34356
rect 33292 34302 33294 34354
rect 33294 34302 33346 34354
rect 33346 34302 33348 34354
rect 33292 34300 33348 34302
rect 33180 33404 33236 33460
rect 33180 33068 33236 33124
rect 33516 33404 33572 33460
rect 33180 31612 33236 31668
rect 32396 31276 32452 31332
rect 32060 28700 32116 28756
rect 31724 27804 31780 27860
rect 31836 27916 31892 27972
rect 31724 27074 31780 27076
rect 31724 27022 31726 27074
rect 31726 27022 31778 27074
rect 31778 27022 31780 27074
rect 31724 27020 31780 27022
rect 31836 26348 31892 26404
rect 31948 24556 32004 24612
rect 32620 30716 32676 30772
rect 32396 29036 32452 29092
rect 32396 28642 32452 28644
rect 32396 28590 32398 28642
rect 32398 28590 32450 28642
rect 32450 28590 32452 28642
rect 32396 28588 32452 28590
rect 32172 27916 32228 27972
rect 32172 27580 32228 27636
rect 33628 32284 33684 32340
rect 33404 32060 33460 32116
rect 34076 34076 34132 34132
rect 33852 33964 33908 34020
rect 34300 33740 34356 33796
rect 33964 33628 34020 33684
rect 34524 33628 34580 33684
rect 33852 33180 33908 33236
rect 33740 31836 33796 31892
rect 33404 31724 33460 31780
rect 33516 31500 33572 31556
rect 33740 31164 33796 31220
rect 34188 32396 34244 32452
rect 32844 29596 32900 29652
rect 33180 29538 33236 29540
rect 33180 29486 33182 29538
rect 33182 29486 33234 29538
rect 33234 29486 33236 29538
rect 33180 29484 33236 29486
rect 33292 29372 33348 29428
rect 33068 29036 33124 29092
rect 33180 28700 33236 28756
rect 33516 30268 33572 30324
rect 34076 31948 34132 32004
rect 33404 29260 33460 29316
rect 33292 28588 33348 28644
rect 34076 30044 34132 30100
rect 33740 28476 33796 28532
rect 33628 28364 33684 28420
rect 34748 34914 34804 34916
rect 34748 34862 34750 34914
rect 34750 34862 34802 34914
rect 34802 34862 34804 34914
rect 34748 34860 34804 34862
rect 34748 33180 34804 33236
rect 34748 32060 34804 32116
rect 34524 30322 34580 30324
rect 34524 30270 34526 30322
rect 34526 30270 34578 30322
rect 34578 30270 34580 30322
rect 34524 30268 34580 30270
rect 34188 29708 34244 29764
rect 34300 29260 34356 29316
rect 34860 29932 34916 29988
rect 39564 37548 39620 37604
rect 35420 34860 35476 34916
rect 35644 34412 35700 34468
rect 36204 34914 36260 34916
rect 36204 34862 36206 34914
rect 36206 34862 36258 34914
rect 36258 34862 36260 34914
rect 36204 34860 36260 34862
rect 35756 31724 35812 31780
rect 36204 33458 36260 33460
rect 36204 33406 36206 33458
rect 36206 33406 36258 33458
rect 36258 33406 36260 33458
rect 36204 33404 36260 33406
rect 36540 35420 36596 35476
rect 36764 35196 36820 35252
rect 36428 34412 36484 34468
rect 36540 34300 36596 34356
rect 36540 34130 36596 34132
rect 36540 34078 36542 34130
rect 36542 34078 36594 34130
rect 36594 34078 36596 34130
rect 36540 34076 36596 34078
rect 36652 33292 36708 33348
rect 36428 33234 36484 33236
rect 36428 33182 36430 33234
rect 36430 33182 36482 33234
rect 36482 33182 36484 33234
rect 36428 33180 36484 33182
rect 35644 31218 35700 31220
rect 35644 31166 35646 31218
rect 35646 31166 35698 31218
rect 35698 31166 35700 31218
rect 35644 31164 35700 31166
rect 36428 32844 36484 32900
rect 36092 30434 36148 30436
rect 36092 30382 36094 30434
rect 36094 30382 36146 30434
rect 36146 30382 36148 30434
rect 36092 30380 36148 30382
rect 35084 30044 35140 30100
rect 36540 31724 36596 31780
rect 36540 30940 36596 30996
rect 36652 30882 36708 30884
rect 36652 30830 36654 30882
rect 36654 30830 36706 30882
rect 36706 30830 36708 30882
rect 36652 30828 36708 30830
rect 36652 30380 36708 30436
rect 35868 29596 35924 29652
rect 36428 30156 36484 30212
rect 34860 29260 34916 29316
rect 34748 28418 34804 28420
rect 34748 28366 34750 28418
rect 34750 28366 34802 28418
rect 34802 28366 34804 28418
rect 34748 28364 34804 28366
rect 34412 28252 34468 28308
rect 33852 27804 33908 27860
rect 32620 26348 32676 26404
rect 32732 26850 32788 26852
rect 32732 26798 32734 26850
rect 32734 26798 32786 26850
rect 32786 26798 32788 26850
rect 32732 26796 32788 26798
rect 33068 26290 33124 26292
rect 33068 26238 33070 26290
rect 33070 26238 33122 26290
rect 33122 26238 33124 26290
rect 33068 26236 33124 26238
rect 33292 26236 33348 26292
rect 32732 25452 32788 25508
rect 31724 24108 31780 24164
rect 31164 23772 31220 23828
rect 31500 23436 31556 23492
rect 30380 21586 30436 21588
rect 30380 21534 30382 21586
rect 30382 21534 30434 21586
rect 30434 21534 30436 21586
rect 30380 21532 30436 21534
rect 30604 22258 30660 22260
rect 30604 22206 30606 22258
rect 30606 22206 30658 22258
rect 30658 22206 30660 22258
rect 30604 22204 30660 22206
rect 31052 22204 31108 22260
rect 30940 21868 30996 21924
rect 31164 21644 31220 21700
rect 30268 21308 30324 21364
rect 30192 21194 30248 21196
rect 30192 21142 30194 21194
rect 30194 21142 30246 21194
rect 30246 21142 30248 21194
rect 30192 21140 30248 21142
rect 30296 21194 30352 21196
rect 30296 21142 30298 21194
rect 30298 21142 30350 21194
rect 30350 21142 30352 21194
rect 30296 21140 30352 21142
rect 30400 21194 30456 21196
rect 30400 21142 30402 21194
rect 30402 21142 30454 21194
rect 30454 21142 30456 21194
rect 30400 21140 30456 21142
rect 30268 20578 30324 20580
rect 30268 20526 30270 20578
rect 30270 20526 30322 20578
rect 30322 20526 30324 20578
rect 30268 20524 30324 20526
rect 30828 20802 30884 20804
rect 30828 20750 30830 20802
rect 30830 20750 30882 20802
rect 30882 20750 30884 20802
rect 30828 20748 30884 20750
rect 31164 21308 31220 21364
rect 31276 21980 31332 22036
rect 31164 20914 31220 20916
rect 31164 20862 31166 20914
rect 31166 20862 31218 20914
rect 31218 20862 31220 20914
rect 31164 20860 31220 20862
rect 31388 20748 31444 20804
rect 31164 20524 31220 20580
rect 30156 20300 30212 20356
rect 30192 19626 30248 19628
rect 30192 19574 30194 19626
rect 30194 19574 30246 19626
rect 30246 19574 30248 19626
rect 30192 19572 30248 19574
rect 30296 19626 30352 19628
rect 30296 19574 30298 19626
rect 30298 19574 30350 19626
rect 30350 19574 30352 19626
rect 30296 19572 30352 19574
rect 30400 19626 30456 19628
rect 30400 19574 30402 19626
rect 30402 19574 30454 19626
rect 30454 19574 30456 19626
rect 30400 19572 30456 19574
rect 30716 19516 30772 19572
rect 30268 19068 30324 19124
rect 30716 18956 30772 19012
rect 30044 18396 30100 18452
rect 30492 18450 30548 18452
rect 30492 18398 30494 18450
rect 30494 18398 30546 18450
rect 30546 18398 30548 18450
rect 30492 18396 30548 18398
rect 30192 18058 30248 18060
rect 30192 18006 30194 18058
rect 30194 18006 30246 18058
rect 30246 18006 30248 18058
rect 30192 18004 30248 18006
rect 30296 18058 30352 18060
rect 30296 18006 30298 18058
rect 30298 18006 30350 18058
rect 30350 18006 30352 18058
rect 30296 18004 30352 18006
rect 30400 18058 30456 18060
rect 30400 18006 30402 18058
rect 30402 18006 30454 18058
rect 30454 18006 30456 18058
rect 30400 18004 30456 18006
rect 29820 17612 29876 17668
rect 30940 20076 30996 20132
rect 30940 19068 30996 19124
rect 31052 18284 31108 18340
rect 30380 17500 30436 17556
rect 30604 16882 30660 16884
rect 30604 16830 30606 16882
rect 30606 16830 30658 16882
rect 30658 16830 30660 16882
rect 30604 16828 30660 16830
rect 29708 15596 29764 15652
rect 29932 15260 29988 15316
rect 30192 16490 30248 16492
rect 30192 16438 30194 16490
rect 30194 16438 30246 16490
rect 30246 16438 30248 16490
rect 30192 16436 30248 16438
rect 30296 16490 30352 16492
rect 30296 16438 30298 16490
rect 30298 16438 30350 16490
rect 30350 16438 30352 16490
rect 30296 16436 30352 16438
rect 30400 16490 30456 16492
rect 30400 16438 30402 16490
rect 30402 16438 30454 16490
rect 30454 16438 30456 16490
rect 30400 16436 30456 16438
rect 31612 23378 31668 23380
rect 31612 23326 31614 23378
rect 31614 23326 31666 23378
rect 31666 23326 31668 23378
rect 31612 23324 31668 23326
rect 32060 23324 32116 23380
rect 31948 23212 32004 23268
rect 33068 24556 33124 24612
rect 32396 23826 32452 23828
rect 32396 23774 32398 23826
rect 32398 23774 32450 23826
rect 32450 23774 32452 23826
rect 32396 23772 32452 23774
rect 32620 23436 32676 23492
rect 33180 23324 33236 23380
rect 33404 25340 33460 25396
rect 33628 24780 33684 24836
rect 34188 27692 34244 27748
rect 34300 27020 34356 27076
rect 33740 24668 33796 24724
rect 33628 24444 33684 24500
rect 33852 24050 33908 24052
rect 33852 23998 33854 24050
rect 33854 23998 33906 24050
rect 33906 23998 33908 24050
rect 33852 23996 33908 23998
rect 33404 23938 33460 23940
rect 33404 23886 33406 23938
rect 33406 23886 33458 23938
rect 33458 23886 33460 23938
rect 33404 23884 33460 23886
rect 33404 23548 33460 23604
rect 34076 24780 34132 24836
rect 34188 24108 34244 24164
rect 33628 23492 33684 23548
rect 33292 23212 33348 23268
rect 32508 23154 32564 23156
rect 32508 23102 32510 23154
rect 32510 23102 32562 23154
rect 32562 23102 32564 23154
rect 32508 23100 32564 23102
rect 31948 21868 32004 21924
rect 32732 21644 32788 21700
rect 31612 21532 31668 21588
rect 31500 18396 31556 18452
rect 31276 17554 31332 17556
rect 31276 17502 31278 17554
rect 31278 17502 31330 17554
rect 31330 17502 31332 17554
rect 31276 17500 31332 17502
rect 30828 16268 30884 16324
rect 29596 15148 29652 15204
rect 28588 14530 28644 14532
rect 28588 14478 28590 14530
rect 28590 14478 28642 14530
rect 28642 14478 28644 14530
rect 28588 14476 28644 14478
rect 28812 14700 28868 14756
rect 28812 14364 28868 14420
rect 28252 13746 28308 13748
rect 28252 13694 28254 13746
rect 28254 13694 28306 13746
rect 28306 13694 28308 13746
rect 28252 13692 28308 13694
rect 28140 12290 28196 12292
rect 28140 12238 28142 12290
rect 28142 12238 28194 12290
rect 28194 12238 28196 12290
rect 28140 12236 28196 12238
rect 27244 11506 27300 11508
rect 27244 11454 27246 11506
rect 27246 11454 27298 11506
rect 27298 11454 27300 11506
rect 27244 11452 27300 11454
rect 27804 11116 27860 11172
rect 28028 11564 28084 11620
rect 28140 11394 28196 11396
rect 28140 11342 28142 11394
rect 28142 11342 28194 11394
rect 28194 11342 28196 11394
rect 28140 11340 28196 11342
rect 28028 11004 28084 11060
rect 27468 10668 27524 10724
rect 26460 9436 26516 9492
rect 27356 8876 27412 8932
rect 26796 8258 26852 8260
rect 26796 8206 26798 8258
rect 26798 8206 26850 8258
rect 26850 8206 26852 8258
rect 26796 8204 26852 8206
rect 27468 8258 27524 8260
rect 27468 8206 27470 8258
rect 27470 8206 27522 8258
rect 27522 8206 27524 8258
rect 27468 8204 27524 8206
rect 26908 7644 26964 7700
rect 27468 7084 27524 7140
rect 26908 6748 26964 6804
rect 28252 10108 28308 10164
rect 29036 13746 29092 13748
rect 29036 13694 29038 13746
rect 29038 13694 29090 13746
rect 29090 13694 29092 13746
rect 29036 13692 29092 13694
rect 28924 13020 28980 13076
rect 28700 12962 28756 12964
rect 28700 12910 28702 12962
rect 28702 12910 28754 12962
rect 28754 12910 28756 12962
rect 28700 12908 28756 12910
rect 28700 12290 28756 12292
rect 28700 12238 28702 12290
rect 28702 12238 28754 12290
rect 28754 12238 28756 12290
rect 28700 12236 28756 12238
rect 28588 12124 28644 12180
rect 28140 8258 28196 8260
rect 28140 8206 28142 8258
rect 28142 8206 28194 8258
rect 28194 8206 28196 8258
rect 28140 8204 28196 8206
rect 26572 6076 26628 6132
rect 27020 6412 27076 6468
rect 26348 5906 26404 5908
rect 26348 5854 26350 5906
rect 26350 5854 26402 5906
rect 26402 5854 26404 5906
rect 26348 5852 26404 5854
rect 26684 5794 26740 5796
rect 26684 5742 26686 5794
rect 26686 5742 26738 5794
rect 26738 5742 26740 5794
rect 26684 5740 26740 5742
rect 26236 5516 26292 5572
rect 27468 6412 27524 6468
rect 27916 6412 27972 6468
rect 28140 5740 28196 5796
rect 27916 5404 27972 5460
rect 28476 11116 28532 11172
rect 29932 14700 29988 14756
rect 30192 14922 30248 14924
rect 30192 14870 30194 14922
rect 30194 14870 30246 14922
rect 30246 14870 30248 14922
rect 30192 14868 30248 14870
rect 30296 14922 30352 14924
rect 30296 14870 30298 14922
rect 30298 14870 30350 14922
rect 30350 14870 30352 14922
rect 30296 14868 30352 14870
rect 30400 14922 30456 14924
rect 30400 14870 30402 14922
rect 30402 14870 30454 14922
rect 30454 14870 30456 14922
rect 30400 14868 30456 14870
rect 30268 14700 30324 14756
rect 29484 14252 29540 14308
rect 30828 14588 30884 14644
rect 30268 14530 30324 14532
rect 30268 14478 30270 14530
rect 30270 14478 30322 14530
rect 30322 14478 30324 14530
rect 30268 14476 30324 14478
rect 30044 13970 30100 13972
rect 30044 13918 30046 13970
rect 30046 13918 30098 13970
rect 30098 13918 30100 13970
rect 30044 13916 30100 13918
rect 29484 13634 29540 13636
rect 29484 13582 29486 13634
rect 29486 13582 29538 13634
rect 29538 13582 29540 13634
rect 29484 13580 29540 13582
rect 30192 13354 30248 13356
rect 30192 13302 30194 13354
rect 30194 13302 30246 13354
rect 30246 13302 30248 13354
rect 30192 13300 30248 13302
rect 30296 13354 30352 13356
rect 30296 13302 30298 13354
rect 30298 13302 30350 13354
rect 30350 13302 30352 13354
rect 30296 13300 30352 13302
rect 30400 13354 30456 13356
rect 30400 13302 30402 13354
rect 30402 13302 30454 13354
rect 30454 13302 30456 13354
rect 30400 13300 30456 13302
rect 29260 12908 29316 12964
rect 29036 12796 29092 12852
rect 29036 11900 29092 11956
rect 30192 11786 30248 11788
rect 30192 11734 30194 11786
rect 30194 11734 30246 11786
rect 30246 11734 30248 11786
rect 30192 11732 30248 11734
rect 30296 11786 30352 11788
rect 30296 11734 30298 11786
rect 30298 11734 30350 11786
rect 30350 11734 30352 11786
rect 30296 11732 30352 11734
rect 30400 11786 30456 11788
rect 30400 11734 30402 11786
rect 30402 11734 30454 11786
rect 30454 11734 30456 11786
rect 30400 11732 30456 11734
rect 29260 11564 29316 11620
rect 29260 11394 29316 11396
rect 29260 11342 29262 11394
rect 29262 11342 29314 11394
rect 29314 11342 29316 11394
rect 29260 11340 29316 11342
rect 30716 13580 30772 13636
rect 30828 12348 30884 12404
rect 30716 11228 30772 11284
rect 30156 11170 30212 11172
rect 30156 11118 30158 11170
rect 30158 11118 30210 11170
rect 30210 11118 30212 11170
rect 30156 11116 30212 11118
rect 29708 11004 29764 11060
rect 28588 10780 28644 10836
rect 28588 10610 28644 10612
rect 28588 10558 28590 10610
rect 28590 10558 28642 10610
rect 28642 10558 28644 10610
rect 28588 10556 28644 10558
rect 28476 9660 28532 9716
rect 29036 8930 29092 8932
rect 29036 8878 29038 8930
rect 29038 8878 29090 8930
rect 29090 8878 29092 8930
rect 29036 8876 29092 8878
rect 30192 10218 30248 10220
rect 30192 10166 30194 10218
rect 30194 10166 30246 10218
rect 30246 10166 30248 10218
rect 30192 10164 30248 10166
rect 30296 10218 30352 10220
rect 30296 10166 30298 10218
rect 30298 10166 30350 10218
rect 30350 10166 30352 10218
rect 30296 10164 30352 10166
rect 30400 10218 30456 10220
rect 30400 10166 30402 10218
rect 30402 10166 30454 10218
rect 30454 10166 30456 10218
rect 30400 10164 30456 10166
rect 30492 9996 30548 10052
rect 30492 9660 30548 9716
rect 31052 16268 31108 16324
rect 31388 16044 31444 16100
rect 31164 15932 31220 15988
rect 32284 21308 32340 21364
rect 33180 21474 33236 21476
rect 33180 21422 33182 21474
rect 33182 21422 33234 21474
rect 33234 21422 33236 21474
rect 33180 21420 33236 21422
rect 32732 20860 32788 20916
rect 32172 20130 32228 20132
rect 32172 20078 32174 20130
rect 32174 20078 32226 20130
rect 32226 20078 32228 20130
rect 32172 20076 32228 20078
rect 33292 20690 33348 20692
rect 33292 20638 33294 20690
rect 33294 20638 33346 20690
rect 33346 20638 33348 20690
rect 33292 20636 33348 20638
rect 32844 20188 32900 20244
rect 32508 20130 32564 20132
rect 32508 20078 32510 20130
rect 32510 20078 32562 20130
rect 32562 20078 32564 20130
rect 32508 20076 32564 20078
rect 32396 19180 32452 19236
rect 32620 17612 32676 17668
rect 31836 16940 31892 16996
rect 32060 16828 32116 16884
rect 32172 16716 32228 16772
rect 31612 15932 31668 15988
rect 31724 15708 31780 15764
rect 31276 15596 31332 15652
rect 31052 13692 31108 13748
rect 31164 14028 31220 14084
rect 31164 13580 31220 13636
rect 31836 15932 31892 15988
rect 31724 15314 31780 15316
rect 31724 15262 31726 15314
rect 31726 15262 31778 15314
rect 31778 15262 31780 15314
rect 31724 15260 31780 15262
rect 31388 13804 31444 13860
rect 31500 13746 31556 13748
rect 31500 13694 31502 13746
rect 31502 13694 31554 13746
rect 31554 13694 31556 13746
rect 31500 13692 31556 13694
rect 31836 13468 31892 13524
rect 31612 13132 31668 13188
rect 32060 15820 32116 15876
rect 32284 16268 32340 16324
rect 32284 15538 32340 15540
rect 32284 15486 32286 15538
rect 32286 15486 32338 15538
rect 32338 15486 32340 15538
rect 32284 15484 32340 15486
rect 32508 15932 32564 15988
rect 31948 12684 32004 12740
rect 32396 14140 32452 14196
rect 31724 12572 31780 12628
rect 32508 13692 32564 13748
rect 32732 16828 32788 16884
rect 33404 20076 33460 20132
rect 33516 21756 33572 21812
rect 35196 28866 35252 28868
rect 35196 28814 35198 28866
rect 35198 28814 35250 28866
rect 35250 28814 35252 28866
rect 35196 28812 35252 28814
rect 35532 29538 35588 29540
rect 35532 29486 35534 29538
rect 35534 29486 35586 29538
rect 35586 29486 35588 29538
rect 35532 29484 35588 29486
rect 35756 29314 35812 29316
rect 35756 29262 35758 29314
rect 35758 29262 35810 29314
rect 35810 29262 35812 29314
rect 35756 29260 35812 29262
rect 35420 28812 35476 28868
rect 35308 28642 35364 28644
rect 35308 28590 35310 28642
rect 35310 28590 35362 28642
rect 35362 28590 35364 28642
rect 35308 28588 35364 28590
rect 36204 29426 36260 29428
rect 36204 29374 36206 29426
rect 36206 29374 36258 29426
rect 36258 29374 36260 29426
rect 36204 29372 36260 29374
rect 35084 28252 35140 28308
rect 35644 28476 35700 28532
rect 35420 28082 35476 28084
rect 35420 28030 35422 28082
rect 35422 28030 35474 28082
rect 35474 28030 35476 28082
rect 35420 28028 35476 28030
rect 34860 27970 34916 27972
rect 34860 27918 34862 27970
rect 34862 27918 34914 27970
rect 34914 27918 34916 27970
rect 34860 27916 34916 27918
rect 34972 27858 35028 27860
rect 34972 27806 34974 27858
rect 34974 27806 35026 27858
rect 35026 27806 35028 27858
rect 34972 27804 35028 27806
rect 34412 25564 34468 25620
rect 34524 27580 34580 27636
rect 34412 24668 34468 24724
rect 34524 23884 34580 23940
rect 34748 27020 34804 27076
rect 34636 23154 34692 23156
rect 34636 23102 34638 23154
rect 34638 23102 34690 23154
rect 34690 23102 34692 23154
rect 34636 23100 34692 23102
rect 34188 22876 34244 22932
rect 34412 22930 34468 22932
rect 34412 22878 34414 22930
rect 34414 22878 34466 22930
rect 34466 22878 34468 22930
rect 34412 22876 34468 22878
rect 34300 21474 34356 21476
rect 34300 21422 34302 21474
rect 34302 21422 34354 21474
rect 34354 21422 34356 21474
rect 34300 21420 34356 21422
rect 34636 22258 34692 22260
rect 34636 22206 34638 22258
rect 34638 22206 34690 22258
rect 34690 22206 34692 22258
rect 34636 22204 34692 22206
rect 35420 27692 35476 27748
rect 35084 27132 35140 27188
rect 35532 26684 35588 26740
rect 35308 26572 35364 26628
rect 35196 25676 35252 25732
rect 35532 25564 35588 25620
rect 35308 25004 35364 25060
rect 35868 27356 35924 27412
rect 35756 27244 35812 27300
rect 35756 26908 35812 26964
rect 35756 25618 35812 25620
rect 35756 25566 35758 25618
rect 35758 25566 35810 25618
rect 35810 25566 35812 25618
rect 35756 25564 35812 25566
rect 35532 23996 35588 24052
rect 34860 23436 34916 23492
rect 35420 23100 35476 23156
rect 36092 28812 36148 28868
rect 36092 28364 36148 28420
rect 36428 28364 36484 28420
rect 36652 28588 36708 28644
rect 37548 35532 37604 35588
rect 36876 35084 36932 35140
rect 36988 35420 37044 35476
rect 36876 34300 36932 34356
rect 37100 34860 37156 34916
rect 36876 32956 36932 33012
rect 37436 34018 37492 34020
rect 37436 33966 37438 34018
rect 37438 33966 37490 34018
rect 37490 33966 37492 34018
rect 37436 33964 37492 33966
rect 37212 33404 37268 33460
rect 37772 35586 37828 35588
rect 37772 35534 37774 35586
rect 37774 35534 37826 35586
rect 37826 35534 37828 35586
rect 37772 35532 37828 35534
rect 37884 35196 37940 35252
rect 38444 35196 38500 35252
rect 38444 34914 38500 34916
rect 38444 34862 38446 34914
rect 38446 34862 38498 34914
rect 38498 34862 38500 34914
rect 38444 34860 38500 34862
rect 38780 35196 38836 35252
rect 38892 35084 38948 35140
rect 37548 33292 37604 33348
rect 37772 33404 37828 33460
rect 37324 33180 37380 33236
rect 37996 33234 38052 33236
rect 37996 33182 37998 33234
rect 37998 33182 38050 33234
rect 38050 33182 38052 33234
rect 37996 33180 38052 33182
rect 37212 32844 37268 32900
rect 37324 32508 37380 32564
rect 37212 32396 37268 32452
rect 37436 31948 37492 32004
rect 36988 31724 37044 31780
rect 36988 31218 37044 31220
rect 36988 31166 36990 31218
rect 36990 31166 37042 31218
rect 37042 31166 37044 31218
rect 36988 31164 37044 31166
rect 37436 30994 37492 30996
rect 37436 30942 37438 30994
rect 37438 30942 37490 30994
rect 37490 30942 37492 30994
rect 37436 30940 37492 30942
rect 37212 30828 37268 30884
rect 36988 29484 37044 29540
rect 36764 28028 36820 28084
rect 36316 26684 36372 26740
rect 36652 26514 36708 26516
rect 36652 26462 36654 26514
rect 36654 26462 36706 26514
rect 36706 26462 36708 26514
rect 36652 26460 36708 26462
rect 36988 29260 37044 29316
rect 37100 28924 37156 28980
rect 37100 27916 37156 27972
rect 37100 27356 37156 27412
rect 38444 33068 38500 33124
rect 38556 32844 38612 32900
rect 39228 35308 39284 35364
rect 39116 35084 39172 35140
rect 38892 33292 38948 33348
rect 38892 32508 38948 32564
rect 38444 32450 38500 32452
rect 38444 32398 38446 32450
rect 38446 32398 38498 32450
rect 38498 32398 38500 32450
rect 38444 32396 38500 32398
rect 39340 34076 39396 34132
rect 39452 33346 39508 33348
rect 39452 33294 39454 33346
rect 39454 33294 39506 33346
rect 39506 33294 39508 33346
rect 39452 33292 39508 33294
rect 39452 32732 39508 32788
rect 39452 32396 39508 32452
rect 39452 31836 39508 31892
rect 39004 31612 39060 31668
rect 37660 30380 37716 30436
rect 37436 30156 37492 30212
rect 37660 30210 37716 30212
rect 37660 30158 37662 30210
rect 37662 30158 37714 30210
rect 37714 30158 37716 30210
rect 37660 30156 37716 30158
rect 37324 30098 37380 30100
rect 37324 30046 37326 30098
rect 37326 30046 37378 30098
rect 37378 30046 37380 30098
rect 37324 30044 37380 30046
rect 37996 30828 38052 30884
rect 37772 30044 37828 30100
rect 37884 30492 37940 30548
rect 37324 28364 37380 28420
rect 37996 30156 38052 30212
rect 38220 30940 38276 30996
rect 38892 30940 38948 30996
rect 38108 29986 38164 29988
rect 38108 29934 38110 29986
rect 38110 29934 38162 29986
rect 38162 29934 38164 29986
rect 38108 29932 38164 29934
rect 38444 29538 38500 29540
rect 38444 29486 38446 29538
rect 38446 29486 38498 29538
rect 38498 29486 38500 29538
rect 38444 29484 38500 29486
rect 38668 29372 38724 29428
rect 39116 31500 39172 31556
rect 39452 30604 39508 30660
rect 39452 30156 39508 30212
rect 39340 29932 39396 29988
rect 38444 29260 38500 29316
rect 37436 27804 37492 27860
rect 37548 28140 37604 28196
rect 37436 27468 37492 27524
rect 37212 25004 37268 25060
rect 36316 24444 36372 24500
rect 35980 23548 36036 23604
rect 36316 24162 36372 24164
rect 36316 24110 36318 24162
rect 36318 24110 36370 24162
rect 36370 24110 36372 24162
rect 36316 24108 36372 24110
rect 36540 23436 36596 23492
rect 34076 20188 34132 20244
rect 33180 19234 33236 19236
rect 33180 19182 33182 19234
rect 33182 19182 33234 19234
rect 33234 19182 33236 19234
rect 33180 19180 33236 19182
rect 33628 19404 33684 19460
rect 33964 20130 34020 20132
rect 33964 20078 33966 20130
rect 33966 20078 34018 20130
rect 34018 20078 34020 20130
rect 33964 20076 34020 20078
rect 33516 18620 33572 18676
rect 33404 17778 33460 17780
rect 33404 17726 33406 17778
rect 33406 17726 33458 17778
rect 33458 17726 33460 17778
rect 33404 17724 33460 17726
rect 32956 16322 33012 16324
rect 32956 16270 32958 16322
rect 32958 16270 33010 16322
rect 33010 16270 33012 16322
rect 32956 16268 33012 16270
rect 33628 17554 33684 17556
rect 33628 17502 33630 17554
rect 33630 17502 33682 17554
rect 33682 17502 33684 17554
rect 33628 17500 33684 17502
rect 33292 16828 33348 16884
rect 33516 16716 33572 16772
rect 33628 16268 33684 16324
rect 33068 16044 33124 16100
rect 33068 15708 33124 15764
rect 33628 15596 33684 15652
rect 33068 14140 33124 14196
rect 33068 13858 33124 13860
rect 33068 13806 33070 13858
rect 33070 13806 33122 13858
rect 33122 13806 33124 13858
rect 33068 13804 33124 13806
rect 34524 20076 34580 20132
rect 34636 19740 34692 19796
rect 34300 18450 34356 18452
rect 34300 18398 34302 18450
rect 34302 18398 34354 18450
rect 34354 18398 34356 18450
rect 34300 18396 34356 18398
rect 34972 18562 35028 18564
rect 34972 18510 34974 18562
rect 34974 18510 35026 18562
rect 35026 18510 35028 18562
rect 34972 18508 35028 18510
rect 34748 17948 34804 18004
rect 34972 17836 35028 17892
rect 34636 17666 34692 17668
rect 34636 17614 34638 17666
rect 34638 17614 34690 17666
rect 34690 17614 34692 17666
rect 34636 17612 34692 17614
rect 34188 17164 34244 17220
rect 34748 17388 34804 17444
rect 34412 16770 34468 16772
rect 34412 16718 34414 16770
rect 34414 16718 34466 16770
rect 34466 16718 34468 16770
rect 34412 16716 34468 16718
rect 33852 16604 33908 16660
rect 34300 16268 34356 16324
rect 33852 15596 33908 15652
rect 33964 15820 34020 15876
rect 33404 14140 33460 14196
rect 33628 13916 33684 13972
rect 33852 13916 33908 13972
rect 33180 13580 33236 13636
rect 34524 15596 34580 15652
rect 34188 15036 34244 15092
rect 34188 14476 34244 14532
rect 34524 14140 34580 14196
rect 34076 13804 34132 13860
rect 34076 13634 34132 13636
rect 34076 13582 34078 13634
rect 34078 13582 34130 13634
rect 34130 13582 34132 13634
rect 34076 13580 34132 13582
rect 33292 13132 33348 13188
rect 32732 12908 32788 12964
rect 31388 12236 31444 12292
rect 31724 11228 31780 11284
rect 30192 8650 30248 8652
rect 30192 8598 30194 8650
rect 30194 8598 30246 8650
rect 30246 8598 30248 8650
rect 30192 8596 30248 8598
rect 30296 8650 30352 8652
rect 30296 8598 30298 8650
rect 30298 8598 30350 8650
rect 30350 8598 30352 8650
rect 30296 8596 30352 8598
rect 30400 8650 30456 8652
rect 30400 8598 30402 8650
rect 30402 8598 30454 8650
rect 30454 8598 30456 8650
rect 30400 8596 30456 8598
rect 29484 6748 29540 6804
rect 29372 6466 29428 6468
rect 29372 6414 29374 6466
rect 29374 6414 29426 6466
rect 29426 6414 29428 6466
rect 29372 6412 29428 6414
rect 28476 5628 28532 5684
rect 27020 4620 27076 4676
rect 25788 4450 25844 4452
rect 25788 4398 25790 4450
rect 25790 4398 25842 4450
rect 25842 4398 25844 4450
rect 25788 4396 25844 4398
rect 25452 4338 25508 4340
rect 25452 4286 25454 4338
rect 25454 4286 25506 4338
rect 25506 4286 25508 4338
rect 25452 4284 25508 4286
rect 28700 4956 28756 5012
rect 27804 4620 27860 4676
rect 28028 4338 28084 4340
rect 28028 4286 28030 4338
rect 28030 4286 28082 4338
rect 28082 4286 28084 4338
rect 28028 4284 28084 4286
rect 25788 4172 25844 4228
rect 25004 2492 25060 2548
rect 29484 5628 29540 5684
rect 30192 7082 30248 7084
rect 30192 7030 30194 7082
rect 30194 7030 30246 7082
rect 30246 7030 30248 7082
rect 30192 7028 30248 7030
rect 30296 7082 30352 7084
rect 30296 7030 30298 7082
rect 30298 7030 30350 7082
rect 30350 7030 30352 7082
rect 30296 7028 30352 7030
rect 30400 7082 30456 7084
rect 30400 7030 30402 7082
rect 30402 7030 30454 7082
rect 30454 7030 30456 7082
rect 30400 7028 30456 7030
rect 30192 5514 30248 5516
rect 30192 5462 30194 5514
rect 30194 5462 30246 5514
rect 30246 5462 30248 5514
rect 30192 5460 30248 5462
rect 30296 5514 30352 5516
rect 30296 5462 30298 5514
rect 30298 5462 30350 5514
rect 30350 5462 30352 5514
rect 30296 5460 30352 5462
rect 30400 5514 30456 5516
rect 30400 5462 30402 5514
rect 30402 5462 30454 5514
rect 30454 5462 30456 5514
rect 30400 5460 30456 5462
rect 29708 5068 29764 5124
rect 31500 9714 31556 9716
rect 31500 9662 31502 9714
rect 31502 9662 31554 9714
rect 31554 9662 31556 9714
rect 31500 9660 31556 9662
rect 31388 8540 31444 8596
rect 32508 11116 32564 11172
rect 32956 12684 33012 12740
rect 32732 12572 32788 12628
rect 32396 9996 32452 10052
rect 32396 9714 32452 9716
rect 32396 9662 32398 9714
rect 32398 9662 32450 9714
rect 32450 9662 32452 9714
rect 32396 9660 32452 9662
rect 33740 12962 33796 12964
rect 33740 12910 33742 12962
rect 33742 12910 33794 12962
rect 33794 12910 33796 12962
rect 33740 12908 33796 12910
rect 33516 12402 33572 12404
rect 33516 12350 33518 12402
rect 33518 12350 33570 12402
rect 33570 12350 33572 12402
rect 33516 12348 33572 12350
rect 33292 12290 33348 12292
rect 33292 12238 33294 12290
rect 33294 12238 33346 12290
rect 33346 12238 33348 12290
rect 33292 12236 33348 12238
rect 33068 11900 33124 11956
rect 32956 8428 33012 8484
rect 31724 6972 31780 7028
rect 31948 5122 32004 5124
rect 31948 5070 31950 5122
rect 31950 5070 32002 5122
rect 32002 5070 32004 5122
rect 31948 5068 32004 5070
rect 30268 4956 30324 5012
rect 31612 5010 31668 5012
rect 31612 4958 31614 5010
rect 31614 4958 31666 5010
rect 31666 4958 31668 5010
rect 31612 4956 31668 4958
rect 32284 4284 32340 4340
rect 30192 3946 30248 3948
rect 30192 3894 30194 3946
rect 30194 3894 30246 3946
rect 30246 3894 30248 3946
rect 30192 3892 30248 3894
rect 30296 3946 30352 3948
rect 30296 3894 30298 3946
rect 30298 3894 30350 3946
rect 30350 3894 30352 3946
rect 30296 3892 30352 3894
rect 30400 3946 30456 3948
rect 30400 3894 30402 3946
rect 30402 3894 30454 3946
rect 30454 3894 30456 3946
rect 30400 3892 30456 3894
rect 29372 2604 29428 2660
rect 33180 8540 33236 8596
rect 32620 6972 32676 7028
rect 33852 12402 33908 12404
rect 33852 12350 33854 12402
rect 33854 12350 33906 12402
rect 33906 12350 33908 12402
rect 33852 12348 33908 12350
rect 34860 13970 34916 13972
rect 34860 13918 34862 13970
rect 34862 13918 34914 13970
rect 34914 13918 34916 13970
rect 34860 13916 34916 13918
rect 34636 13468 34692 13524
rect 34748 13692 34804 13748
rect 34972 13692 35028 13748
rect 34636 12962 34692 12964
rect 34636 12910 34638 12962
rect 34638 12910 34690 12962
rect 34690 12910 34692 12962
rect 34636 12908 34692 12910
rect 34524 12402 34580 12404
rect 34524 12350 34526 12402
rect 34526 12350 34578 12402
rect 34578 12350 34580 12402
rect 34524 12348 34580 12350
rect 33404 11676 33460 11732
rect 34188 11676 34244 11732
rect 34188 11228 34244 11284
rect 34076 8540 34132 8596
rect 33740 7308 33796 7364
rect 34412 7362 34468 7364
rect 34412 7310 34414 7362
rect 34414 7310 34466 7362
rect 34466 7310 34468 7362
rect 34412 7308 34468 7310
rect 33292 6300 33348 6356
rect 34188 6860 34244 6916
rect 33628 5906 33684 5908
rect 33628 5854 33630 5906
rect 33630 5854 33682 5906
rect 33682 5854 33684 5906
rect 33628 5852 33684 5854
rect 33292 4956 33348 5012
rect 34300 5906 34356 5908
rect 34300 5854 34302 5906
rect 34302 5854 34354 5906
rect 34354 5854 34356 5906
rect 34300 5852 34356 5854
rect 35308 21756 35364 21812
rect 35980 21980 36036 22036
rect 36428 23324 36484 23380
rect 36652 23266 36708 23268
rect 36652 23214 36654 23266
rect 36654 23214 36706 23266
rect 36706 23214 36708 23266
rect 36652 23212 36708 23214
rect 36540 21980 36596 22036
rect 37212 23996 37268 24052
rect 37100 23548 37156 23604
rect 36764 22876 36820 22932
rect 38220 28588 38276 28644
rect 38668 28588 38724 28644
rect 38108 28140 38164 28196
rect 37996 27692 38052 27748
rect 38780 28364 38836 28420
rect 39004 29484 39060 29540
rect 39340 29372 39396 29428
rect 39004 28700 39060 28756
rect 39116 28588 39172 28644
rect 38892 28140 38948 28196
rect 38668 27916 38724 27972
rect 37660 27020 37716 27076
rect 37884 27074 37940 27076
rect 37884 27022 37886 27074
rect 37886 27022 37938 27074
rect 37938 27022 37940 27074
rect 37884 27020 37940 27022
rect 38332 27356 38388 27412
rect 38556 27580 38612 27636
rect 37548 25900 37604 25956
rect 37996 25788 38052 25844
rect 38108 25900 38164 25956
rect 38108 25340 38164 25396
rect 41580 37436 41636 37492
rect 39852 36090 39908 36092
rect 39852 36038 39854 36090
rect 39854 36038 39906 36090
rect 39906 36038 39908 36090
rect 39852 36036 39908 36038
rect 39956 36090 40012 36092
rect 39956 36038 39958 36090
rect 39958 36038 40010 36090
rect 40010 36038 40012 36090
rect 39956 36036 40012 36038
rect 40060 36090 40116 36092
rect 40060 36038 40062 36090
rect 40062 36038 40114 36090
rect 40114 36038 40116 36090
rect 40060 36036 40116 36038
rect 40012 34860 40068 34916
rect 40236 35196 40292 35252
rect 40572 35532 40628 35588
rect 40460 35084 40516 35140
rect 40348 34748 40404 34804
rect 39852 34522 39908 34524
rect 39852 34470 39854 34522
rect 39854 34470 39906 34522
rect 39906 34470 39908 34522
rect 39852 34468 39908 34470
rect 39956 34522 40012 34524
rect 39956 34470 39958 34522
rect 39958 34470 40010 34522
rect 40010 34470 40012 34522
rect 39956 34468 40012 34470
rect 40060 34522 40116 34524
rect 40060 34470 40062 34522
rect 40062 34470 40114 34522
rect 40114 34470 40116 34522
rect 40060 34468 40116 34470
rect 39676 34018 39732 34020
rect 39676 33966 39678 34018
rect 39678 33966 39730 34018
rect 39730 33966 39732 34018
rect 39676 33964 39732 33966
rect 39852 32954 39908 32956
rect 39852 32902 39854 32954
rect 39854 32902 39906 32954
rect 39906 32902 39908 32954
rect 39852 32900 39908 32902
rect 39956 32954 40012 32956
rect 39956 32902 39958 32954
rect 39958 32902 40010 32954
rect 40010 32902 40012 32954
rect 39956 32900 40012 32902
rect 40060 32954 40116 32956
rect 40060 32902 40062 32954
rect 40062 32902 40114 32954
rect 40114 32902 40116 32954
rect 40060 32900 40116 32902
rect 39676 32562 39732 32564
rect 39676 32510 39678 32562
rect 39678 32510 39730 32562
rect 39730 32510 39732 32562
rect 39676 32508 39732 32510
rect 39900 32620 39956 32676
rect 40236 32620 40292 32676
rect 39788 31836 39844 31892
rect 39852 31386 39908 31388
rect 39852 31334 39854 31386
rect 39854 31334 39906 31386
rect 39906 31334 39908 31386
rect 39852 31332 39908 31334
rect 39956 31386 40012 31388
rect 39956 31334 39958 31386
rect 39958 31334 40010 31386
rect 40010 31334 40012 31386
rect 39956 31332 40012 31334
rect 40060 31386 40116 31388
rect 40060 31334 40062 31386
rect 40062 31334 40114 31386
rect 40114 31334 40116 31386
rect 40060 31332 40116 31334
rect 40012 31218 40068 31220
rect 40012 31166 40014 31218
rect 40014 31166 40066 31218
rect 40066 31166 40068 31218
rect 40012 31164 40068 31166
rect 39788 30994 39844 30996
rect 39788 30942 39790 30994
rect 39790 30942 39842 30994
rect 39842 30942 39844 30994
rect 39788 30940 39844 30942
rect 40236 29932 40292 29988
rect 39852 29818 39908 29820
rect 39852 29766 39854 29818
rect 39854 29766 39906 29818
rect 39906 29766 39908 29818
rect 39852 29764 39908 29766
rect 39956 29818 40012 29820
rect 39956 29766 39958 29818
rect 39958 29766 40010 29818
rect 40010 29766 40012 29818
rect 39956 29764 40012 29766
rect 40060 29818 40116 29820
rect 40060 29766 40062 29818
rect 40062 29766 40114 29818
rect 40114 29766 40116 29818
rect 40060 29764 40116 29766
rect 40012 29650 40068 29652
rect 40012 29598 40014 29650
rect 40014 29598 40066 29650
rect 40066 29598 40068 29650
rect 40012 29596 40068 29598
rect 39564 28588 39620 28644
rect 39788 29372 39844 29428
rect 39228 28028 39284 28084
rect 39564 27916 39620 27972
rect 40124 28812 40180 28868
rect 39788 28700 39844 28756
rect 40348 29372 40404 29428
rect 40460 28588 40516 28644
rect 39900 28418 39956 28420
rect 39900 28366 39902 28418
rect 39902 28366 39954 28418
rect 39954 28366 39956 28418
rect 39900 28364 39956 28366
rect 39852 28250 39908 28252
rect 39852 28198 39854 28250
rect 39854 28198 39906 28250
rect 39906 28198 39908 28250
rect 39852 28196 39908 28198
rect 39956 28250 40012 28252
rect 39956 28198 39958 28250
rect 39958 28198 40010 28250
rect 40010 28198 40012 28250
rect 39956 28196 40012 28198
rect 40060 28250 40116 28252
rect 40060 28198 40062 28250
rect 40062 28198 40114 28250
rect 40114 28198 40116 28250
rect 40060 28196 40116 28198
rect 39900 28028 39956 28084
rect 38780 27804 38836 27860
rect 38668 26572 38724 26628
rect 38444 25788 38500 25844
rect 38780 26684 38836 26740
rect 39340 27746 39396 27748
rect 39340 27694 39342 27746
rect 39342 27694 39394 27746
rect 39394 27694 39396 27746
rect 39340 27692 39396 27694
rect 39004 27468 39060 27524
rect 39116 27356 39172 27412
rect 39340 27468 39396 27524
rect 39676 27468 39732 27524
rect 40124 27634 40180 27636
rect 40124 27582 40126 27634
rect 40126 27582 40178 27634
rect 40178 27582 40180 27634
rect 40124 27580 40180 27582
rect 39340 27074 39396 27076
rect 39340 27022 39342 27074
rect 39342 27022 39394 27074
rect 39394 27022 39396 27074
rect 39340 27020 39396 27022
rect 39340 26850 39396 26852
rect 39340 26798 39342 26850
rect 39342 26798 39394 26850
rect 39394 26798 39396 26850
rect 39340 26796 39396 26798
rect 38556 25340 38612 25396
rect 38668 25900 38724 25956
rect 38220 25282 38276 25284
rect 38220 25230 38222 25282
rect 38222 25230 38274 25282
rect 38274 25230 38276 25282
rect 38220 25228 38276 25230
rect 38444 24780 38500 24836
rect 37436 24444 37492 24500
rect 37884 24444 37940 24500
rect 38220 24668 38276 24724
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 38108 23772 38164 23828
rect 38108 23548 38164 23604
rect 36204 21756 36260 21812
rect 36428 21586 36484 21588
rect 36428 21534 36430 21586
rect 36430 21534 36482 21586
rect 36482 21534 36484 21586
rect 36428 21532 36484 21534
rect 36204 21196 36260 21252
rect 36316 21420 36372 21476
rect 35420 20636 35476 20692
rect 36428 20860 36484 20916
rect 36428 20636 36484 20692
rect 36316 20524 36372 20580
rect 35420 19740 35476 19796
rect 35308 19628 35364 19684
rect 35196 17388 35252 17444
rect 36988 22258 37044 22260
rect 36988 22206 36990 22258
rect 36990 22206 37042 22258
rect 37042 22206 37044 22258
rect 36988 22204 37044 22206
rect 36764 19852 36820 19908
rect 36428 19234 36484 19236
rect 36428 19182 36430 19234
rect 36430 19182 36482 19234
rect 36482 19182 36484 19234
rect 36428 19180 36484 19182
rect 35532 17500 35588 17556
rect 37100 21532 37156 21588
rect 36988 21420 37044 21476
rect 36876 18732 36932 18788
rect 35644 17724 35700 17780
rect 35420 17052 35476 17108
rect 35532 16770 35588 16772
rect 35532 16718 35534 16770
rect 35534 16718 35586 16770
rect 35586 16718 35588 16770
rect 35532 16716 35588 16718
rect 35308 16380 35364 16436
rect 35196 15820 35252 15876
rect 35196 13692 35252 13748
rect 35420 16156 35476 16212
rect 35644 16044 35700 16100
rect 35868 17948 35924 18004
rect 36092 17836 36148 17892
rect 36204 17500 36260 17556
rect 36540 17836 36596 17892
rect 36316 16268 36372 16324
rect 36428 17164 36484 17220
rect 35980 15874 36036 15876
rect 35980 15822 35982 15874
rect 35982 15822 36034 15874
rect 36034 15822 36036 15874
rect 35980 15820 36036 15822
rect 37548 20300 37604 20356
rect 37324 18508 37380 18564
rect 37436 18732 37492 18788
rect 37660 18732 37716 18788
rect 36988 17948 37044 18004
rect 37212 17612 37268 17668
rect 36652 15932 36708 15988
rect 36764 16828 36820 16884
rect 37548 17276 37604 17332
rect 36988 16716 37044 16772
rect 37436 16716 37492 16772
rect 36764 15202 36820 15204
rect 36764 15150 36766 15202
rect 36766 15150 36818 15202
rect 36818 15150 36820 15202
rect 36764 15148 36820 15150
rect 35644 14530 35700 14532
rect 35644 14478 35646 14530
rect 35646 14478 35698 14530
rect 35698 14478 35700 14530
rect 35644 14476 35700 14478
rect 36204 14530 36260 14532
rect 36204 14478 36206 14530
rect 36206 14478 36258 14530
rect 36258 14478 36260 14530
rect 36204 14476 36260 14478
rect 37100 14028 37156 14084
rect 35308 13132 35364 13188
rect 35420 13804 35476 13860
rect 35308 12962 35364 12964
rect 35308 12910 35310 12962
rect 35310 12910 35362 12962
rect 35362 12910 35364 12962
rect 35308 12908 35364 12910
rect 35644 13858 35700 13860
rect 35644 13806 35646 13858
rect 35646 13806 35698 13858
rect 35698 13806 35700 13858
rect 35644 13804 35700 13806
rect 35644 12684 35700 12740
rect 34860 9772 34916 9828
rect 34972 9212 35028 9268
rect 35084 12124 35140 12180
rect 34972 8540 35028 8596
rect 34860 7196 34916 7252
rect 34748 6860 34804 6916
rect 35196 6860 35252 6916
rect 35084 6412 35140 6468
rect 32508 4284 32564 4340
rect 33628 4338 33684 4340
rect 33628 4286 33630 4338
rect 33630 4286 33682 4338
rect 33682 4286 33684 4338
rect 33628 4284 33684 4286
rect 35420 5122 35476 5124
rect 35420 5070 35422 5122
rect 35422 5070 35474 5122
rect 35474 5070 35476 5122
rect 35420 5068 35476 5070
rect 35644 9042 35700 9044
rect 35644 8990 35646 9042
rect 35646 8990 35698 9042
rect 35698 8990 35700 9042
rect 35644 8988 35700 8990
rect 35644 8092 35700 8148
rect 37100 13468 37156 13524
rect 36316 13132 36372 13188
rect 35980 12684 36036 12740
rect 37212 13074 37268 13076
rect 37212 13022 37214 13074
rect 37214 13022 37266 13074
rect 37266 13022 37268 13074
rect 37212 13020 37268 13022
rect 36428 12460 36484 12516
rect 36092 12348 36148 12404
rect 36204 11788 36260 11844
rect 36428 11170 36484 11172
rect 36428 11118 36430 11170
rect 36430 11118 36482 11170
rect 36482 11118 36484 11170
rect 36428 11116 36484 11118
rect 36988 11004 37044 11060
rect 35868 9772 35924 9828
rect 36204 9042 36260 9044
rect 36204 8990 36206 9042
rect 36206 8990 36258 9042
rect 36258 8990 36260 9042
rect 36204 8988 36260 8990
rect 37436 15596 37492 15652
rect 37772 15148 37828 15204
rect 37548 13970 37604 13972
rect 37548 13918 37550 13970
rect 37550 13918 37602 13970
rect 37602 13918 37604 13970
rect 37548 13916 37604 13918
rect 39004 25900 39060 25956
rect 38780 25788 38836 25844
rect 38780 25452 38836 25508
rect 38892 25394 38948 25396
rect 38892 25342 38894 25394
rect 38894 25342 38946 25394
rect 38946 25342 38948 25394
rect 38892 25340 38948 25342
rect 39116 25394 39172 25396
rect 39116 25342 39118 25394
rect 39118 25342 39170 25394
rect 39170 25342 39172 25394
rect 39116 25340 39172 25342
rect 38556 24108 38612 24164
rect 38780 23938 38836 23940
rect 38780 23886 38782 23938
rect 38782 23886 38834 23938
rect 38834 23886 38836 23938
rect 38780 23884 38836 23886
rect 38780 23212 38836 23268
rect 39116 23884 39172 23940
rect 38892 22988 38948 23044
rect 39004 22876 39060 22932
rect 38444 21698 38500 21700
rect 38444 21646 38446 21698
rect 38446 21646 38498 21698
rect 38498 21646 38500 21698
rect 38444 21644 38500 21646
rect 38780 21810 38836 21812
rect 38780 21758 38782 21810
rect 38782 21758 38834 21810
rect 38834 21758 38836 21810
rect 38780 21756 38836 21758
rect 38220 19404 38276 19460
rect 38108 19010 38164 19012
rect 38108 18958 38110 19010
rect 38110 18958 38162 19010
rect 38162 18958 38164 19010
rect 38108 18956 38164 18958
rect 37996 18450 38052 18452
rect 37996 18398 37998 18450
rect 37998 18398 38050 18450
rect 38050 18398 38052 18450
rect 37996 18396 38052 18398
rect 38220 16098 38276 16100
rect 38220 16046 38222 16098
rect 38222 16046 38274 16098
rect 38274 16046 38276 16098
rect 38220 16044 38276 16046
rect 38332 15596 38388 15652
rect 38108 14700 38164 14756
rect 37996 14642 38052 14644
rect 37996 14590 37998 14642
rect 37998 14590 38050 14642
rect 38050 14590 38052 14642
rect 37996 14588 38052 14590
rect 37772 13132 37828 13188
rect 37324 11676 37380 11732
rect 37324 11170 37380 11172
rect 37324 11118 37326 11170
rect 37326 11118 37378 11170
rect 37378 11118 37380 11170
rect 37324 11116 37380 11118
rect 36988 8316 37044 8372
rect 37324 9772 37380 9828
rect 37772 12124 37828 12180
rect 38892 21420 38948 21476
rect 39340 24668 39396 24724
rect 39900 26962 39956 26964
rect 39900 26910 39902 26962
rect 39902 26910 39954 26962
rect 39954 26910 39956 26962
rect 39900 26908 39956 26910
rect 39788 26850 39844 26852
rect 39788 26798 39790 26850
rect 39790 26798 39842 26850
rect 39842 26798 39844 26850
rect 39788 26796 39844 26798
rect 39676 26684 39732 26740
rect 39852 26682 39908 26684
rect 39564 26572 39620 26628
rect 39852 26630 39854 26682
rect 39854 26630 39906 26682
rect 39906 26630 39908 26682
rect 39852 26628 39908 26630
rect 39956 26682 40012 26684
rect 39956 26630 39958 26682
rect 39958 26630 40010 26682
rect 40010 26630 40012 26682
rect 39956 26628 40012 26630
rect 40060 26682 40116 26684
rect 40060 26630 40062 26682
rect 40062 26630 40114 26682
rect 40114 26630 40116 26682
rect 40060 26628 40116 26630
rect 39676 26236 39732 26292
rect 39564 25788 39620 25844
rect 39228 23772 39284 23828
rect 39340 23436 39396 23492
rect 39340 23212 39396 23268
rect 38780 20412 38836 20468
rect 39228 21420 39284 21476
rect 38556 17388 38612 17444
rect 38892 18396 38948 18452
rect 38668 17164 38724 17220
rect 38892 16828 38948 16884
rect 38668 16492 38724 16548
rect 38556 14754 38612 14756
rect 38556 14702 38558 14754
rect 38558 14702 38610 14754
rect 38610 14702 38612 14754
rect 38556 14700 38612 14702
rect 39116 19068 39172 19124
rect 39340 20972 39396 21028
rect 39452 22204 39508 22260
rect 39452 19180 39508 19236
rect 39340 17554 39396 17556
rect 39340 17502 39342 17554
rect 39342 17502 39394 17554
rect 39394 17502 39396 17554
rect 39340 17500 39396 17502
rect 39116 16098 39172 16100
rect 39116 16046 39118 16098
rect 39118 16046 39170 16098
rect 39170 16046 39172 16098
rect 39116 16044 39172 16046
rect 40124 26460 40180 26516
rect 39788 25452 39844 25508
rect 40012 26012 40068 26068
rect 41244 34860 41300 34916
rect 41132 34748 41188 34804
rect 41244 34354 41300 34356
rect 41244 34302 41246 34354
rect 41246 34302 41298 34354
rect 41298 34302 41300 34354
rect 41244 34300 41300 34302
rect 41132 33852 41188 33908
rect 41468 33964 41524 34020
rect 41356 32508 41412 32564
rect 40796 31276 40852 31332
rect 40684 28866 40740 28868
rect 40684 28814 40686 28866
rect 40686 28814 40738 28866
rect 40738 28814 40740 28866
rect 40684 28812 40740 28814
rect 40348 26012 40404 26068
rect 40348 25340 40404 25396
rect 39852 25114 39908 25116
rect 39852 25062 39854 25114
rect 39854 25062 39906 25114
rect 39906 25062 39908 25114
rect 39852 25060 39908 25062
rect 39956 25114 40012 25116
rect 39956 25062 39958 25114
rect 39958 25062 40010 25114
rect 40010 25062 40012 25114
rect 39956 25060 40012 25062
rect 40060 25114 40116 25116
rect 40060 25062 40062 25114
rect 40062 25062 40114 25114
rect 40114 25062 40116 25114
rect 40060 25060 40116 25062
rect 39676 24722 39732 24724
rect 39676 24670 39678 24722
rect 39678 24670 39730 24722
rect 39730 24670 39732 24722
rect 39676 24668 39732 24670
rect 40012 24834 40068 24836
rect 40012 24782 40014 24834
rect 40014 24782 40066 24834
rect 40066 24782 40068 24834
rect 40012 24780 40068 24782
rect 41244 31164 41300 31220
rect 41020 30994 41076 30996
rect 41020 30942 41022 30994
rect 41022 30942 41074 30994
rect 41074 30942 41076 30994
rect 41020 30940 41076 30942
rect 42476 37324 42532 37380
rect 42140 35308 42196 35364
rect 41916 34354 41972 34356
rect 41916 34302 41918 34354
rect 41918 34302 41970 34354
rect 41970 34302 41972 34354
rect 41916 34300 41972 34302
rect 42028 33964 42084 34020
rect 41692 32620 41748 32676
rect 42364 32396 42420 32452
rect 42364 31836 42420 31892
rect 42252 30828 42308 30884
rect 44380 37212 44436 37268
rect 43036 36482 43092 36484
rect 43036 36430 43038 36482
rect 43038 36430 43090 36482
rect 43090 36430 43092 36482
rect 43036 36428 43092 36430
rect 43260 35532 43316 35588
rect 43036 35026 43092 35028
rect 43036 34974 43038 35026
rect 43038 34974 43090 35026
rect 43090 34974 43092 35026
rect 43036 34972 43092 34974
rect 42588 34802 42644 34804
rect 42588 34750 42590 34802
rect 42590 34750 42642 34802
rect 42642 34750 42644 34802
rect 42588 34748 42644 34750
rect 42588 33740 42644 33796
rect 43036 33404 43092 33460
rect 42700 32732 42756 32788
rect 43036 32786 43092 32788
rect 43036 32734 43038 32786
rect 43038 32734 43090 32786
rect 43090 32734 43092 32786
rect 43036 32732 43092 32734
rect 42700 32450 42756 32452
rect 42700 32398 42702 32450
rect 42702 32398 42754 32450
rect 42754 32398 42756 32450
rect 42700 32396 42756 32398
rect 42476 30940 42532 30996
rect 41804 30268 41860 30324
rect 41580 30156 41636 30212
rect 41468 29596 41524 29652
rect 41916 29708 41972 29764
rect 41020 28588 41076 28644
rect 39900 24108 39956 24164
rect 39852 23546 39908 23548
rect 39852 23494 39854 23546
rect 39854 23494 39906 23546
rect 39906 23494 39908 23546
rect 39852 23492 39908 23494
rect 39956 23546 40012 23548
rect 39956 23494 39958 23546
rect 39958 23494 40010 23546
rect 40010 23494 40012 23546
rect 39956 23492 40012 23494
rect 40060 23546 40116 23548
rect 40060 23494 40062 23546
rect 40062 23494 40114 23546
rect 40114 23494 40116 23546
rect 40060 23492 40116 23494
rect 40460 23884 40516 23940
rect 39676 23266 39732 23268
rect 39676 23214 39678 23266
rect 39678 23214 39730 23266
rect 39730 23214 39732 23266
rect 39676 23212 39732 23214
rect 40124 23154 40180 23156
rect 40124 23102 40126 23154
rect 40126 23102 40178 23154
rect 40178 23102 40180 23154
rect 40124 23100 40180 23102
rect 39788 22876 39844 22932
rect 39900 22988 39956 23044
rect 39676 22540 39732 22596
rect 39900 22370 39956 22372
rect 39900 22318 39902 22370
rect 39902 22318 39954 22370
rect 39954 22318 39956 22370
rect 39900 22316 39956 22318
rect 39788 22204 39844 22260
rect 39852 21978 39908 21980
rect 39852 21926 39854 21978
rect 39854 21926 39906 21978
rect 39906 21926 39908 21978
rect 39852 21924 39908 21926
rect 39956 21978 40012 21980
rect 39956 21926 39958 21978
rect 39958 21926 40010 21978
rect 40010 21926 40012 21978
rect 39956 21924 40012 21926
rect 40060 21978 40116 21980
rect 40060 21926 40062 21978
rect 40062 21926 40114 21978
rect 40114 21926 40116 21978
rect 40060 21924 40116 21926
rect 40348 21756 40404 21812
rect 40460 21868 40516 21924
rect 40124 21420 40180 21476
rect 40236 20860 40292 20916
rect 40124 20690 40180 20692
rect 40124 20638 40126 20690
rect 40126 20638 40178 20690
rect 40178 20638 40180 20690
rect 40124 20636 40180 20638
rect 39852 20410 39908 20412
rect 39852 20358 39854 20410
rect 39854 20358 39906 20410
rect 39906 20358 39908 20410
rect 39852 20356 39908 20358
rect 39956 20410 40012 20412
rect 39956 20358 39958 20410
rect 39958 20358 40010 20410
rect 40010 20358 40012 20410
rect 39956 20356 40012 20358
rect 40060 20410 40116 20412
rect 40060 20358 40062 20410
rect 40062 20358 40114 20410
rect 40114 20358 40116 20410
rect 40060 20356 40116 20358
rect 40460 20076 40516 20132
rect 39852 18842 39908 18844
rect 39852 18790 39854 18842
rect 39854 18790 39906 18842
rect 39906 18790 39908 18842
rect 39852 18788 39908 18790
rect 39956 18842 40012 18844
rect 39956 18790 39958 18842
rect 39958 18790 40010 18842
rect 40010 18790 40012 18842
rect 39956 18788 40012 18790
rect 40060 18842 40116 18844
rect 40060 18790 40062 18842
rect 40062 18790 40114 18842
rect 40114 18790 40116 18842
rect 40060 18788 40116 18790
rect 40012 18450 40068 18452
rect 40012 18398 40014 18450
rect 40014 18398 40066 18450
rect 40066 18398 40068 18450
rect 40012 18396 40068 18398
rect 40684 27692 40740 27748
rect 40796 27356 40852 27412
rect 41692 28812 41748 28868
rect 41580 28754 41636 28756
rect 41580 28702 41582 28754
rect 41582 28702 41634 28754
rect 41634 28702 41636 28754
rect 41580 28700 41636 28702
rect 41804 29036 41860 29092
rect 41468 27858 41524 27860
rect 41468 27806 41470 27858
rect 41470 27806 41522 27858
rect 41522 27806 41524 27858
rect 41468 27804 41524 27806
rect 41356 27244 41412 27300
rect 41356 27020 41412 27076
rect 40684 26460 40740 26516
rect 40684 26236 40740 26292
rect 40908 25340 40964 25396
rect 40908 25116 40964 25172
rect 40908 24780 40964 24836
rect 40908 24444 40964 24500
rect 40684 23772 40740 23828
rect 40908 24108 40964 24164
rect 40796 23324 40852 23380
rect 40796 22540 40852 22596
rect 40684 22316 40740 22372
rect 40684 21756 40740 21812
rect 41020 23100 41076 23156
rect 41692 26962 41748 26964
rect 41692 26910 41694 26962
rect 41694 26910 41746 26962
rect 41746 26910 41748 26962
rect 41692 26908 41748 26910
rect 42252 30604 42308 30660
rect 42476 30268 42532 30324
rect 42588 30210 42644 30212
rect 42588 30158 42590 30210
rect 42590 30158 42642 30210
rect 42642 30158 42644 30210
rect 42588 30156 42644 30158
rect 44268 35586 44324 35588
rect 44268 35534 44270 35586
rect 44270 35534 44322 35586
rect 44322 35534 44324 35586
rect 44268 35532 44324 35534
rect 44156 35308 44212 35364
rect 43708 34914 43764 34916
rect 43708 34862 43710 34914
rect 43710 34862 43762 34914
rect 43762 34862 43764 34914
rect 43708 34860 43764 34862
rect 43484 34802 43540 34804
rect 43484 34750 43486 34802
rect 43486 34750 43538 34802
rect 43538 34750 43540 34802
rect 43484 34748 43540 34750
rect 44044 34802 44100 34804
rect 44044 34750 44046 34802
rect 44046 34750 44098 34802
rect 44098 34750 44100 34802
rect 44044 34748 44100 34750
rect 44380 35196 44436 35252
rect 44268 34972 44324 35028
rect 44156 34354 44212 34356
rect 44156 34302 44158 34354
rect 44158 34302 44210 34354
rect 44210 34302 44212 34354
rect 44156 34300 44212 34302
rect 43484 34242 43540 34244
rect 43484 34190 43486 34242
rect 43486 34190 43538 34242
rect 43538 34190 43540 34242
rect 43484 34188 43540 34190
rect 43484 33458 43540 33460
rect 43484 33406 43486 33458
rect 43486 33406 43538 33458
rect 43538 33406 43540 33458
rect 43484 33404 43540 33406
rect 43932 32732 43988 32788
rect 43484 31666 43540 31668
rect 43484 31614 43486 31666
rect 43486 31614 43538 31666
rect 43538 31614 43540 31666
rect 43484 31612 43540 31614
rect 43708 31500 43764 31556
rect 43932 31554 43988 31556
rect 43932 31502 43934 31554
rect 43934 31502 43986 31554
rect 43986 31502 43988 31554
rect 43932 31500 43988 31502
rect 43820 30994 43876 30996
rect 43820 30942 43822 30994
rect 43822 30942 43874 30994
rect 43874 30942 43876 30994
rect 43820 30940 43876 30942
rect 44268 30994 44324 30996
rect 44268 30942 44270 30994
rect 44270 30942 44322 30994
rect 44322 30942 44324 30994
rect 44268 30940 44324 30942
rect 43148 30716 43204 30772
rect 43148 30044 43204 30100
rect 43596 30098 43652 30100
rect 43596 30046 43598 30098
rect 43598 30046 43650 30098
rect 43650 30046 43652 30098
rect 43596 30044 43652 30046
rect 43820 30098 43876 30100
rect 43820 30046 43822 30098
rect 43822 30046 43874 30098
rect 43874 30046 43876 30098
rect 43820 30044 43876 30046
rect 44044 29986 44100 29988
rect 44044 29934 44046 29986
rect 44046 29934 44098 29986
rect 44098 29934 44100 29986
rect 44044 29932 44100 29934
rect 43260 29820 43316 29876
rect 43820 29820 43876 29876
rect 42588 29372 42644 29428
rect 42364 28812 42420 28868
rect 43484 28364 43540 28420
rect 43260 28140 43316 28196
rect 42476 27858 42532 27860
rect 42476 27806 42478 27858
rect 42478 27806 42530 27858
rect 42530 27806 42532 27858
rect 42476 27804 42532 27806
rect 41916 25788 41972 25844
rect 41356 25564 41412 25620
rect 41692 25116 41748 25172
rect 41356 24498 41412 24500
rect 41356 24446 41358 24498
rect 41358 24446 41410 24498
rect 41410 24446 41412 24498
rect 41356 24444 41412 24446
rect 41804 24332 41860 24388
rect 41468 24220 41524 24276
rect 41692 23938 41748 23940
rect 41692 23886 41694 23938
rect 41694 23886 41746 23938
rect 41746 23886 41748 23938
rect 41692 23884 41748 23886
rect 41244 23772 41300 23828
rect 41468 23378 41524 23380
rect 41468 23326 41470 23378
rect 41470 23326 41522 23378
rect 41522 23326 41524 23378
rect 41468 23324 41524 23326
rect 41244 22988 41300 23044
rect 41356 21644 41412 21700
rect 41916 23042 41972 23044
rect 41916 22990 41918 23042
rect 41918 22990 41970 23042
rect 41970 22990 41972 23042
rect 41916 22988 41972 22990
rect 40460 19292 40516 19348
rect 40572 19404 40628 19460
rect 40348 18338 40404 18340
rect 40348 18286 40350 18338
rect 40350 18286 40402 18338
rect 40402 18286 40404 18338
rect 40348 18284 40404 18286
rect 40348 18060 40404 18116
rect 40236 17836 40292 17892
rect 39852 17274 39908 17276
rect 39852 17222 39854 17274
rect 39854 17222 39906 17274
rect 39906 17222 39908 17274
rect 39852 17220 39908 17222
rect 39956 17274 40012 17276
rect 39956 17222 39958 17274
rect 39958 17222 40010 17274
rect 40010 17222 40012 17274
rect 39956 17220 40012 17222
rect 40060 17274 40116 17276
rect 40060 17222 40062 17274
rect 40062 17222 40114 17274
rect 40114 17222 40116 17274
rect 40060 17220 40116 17222
rect 40684 18956 40740 19012
rect 42140 22370 42196 22372
rect 42140 22318 42142 22370
rect 42142 22318 42194 22370
rect 42194 22318 42196 22370
rect 42140 22316 42196 22318
rect 41916 21868 41972 21924
rect 41804 21756 41860 21812
rect 42140 20972 42196 21028
rect 41356 20076 41412 20132
rect 41132 19516 41188 19572
rect 40684 18060 40740 18116
rect 40796 18284 40852 18340
rect 40684 17890 40740 17892
rect 40684 17838 40686 17890
rect 40686 17838 40738 17890
rect 40738 17838 40740 17890
rect 40684 17836 40740 17838
rect 40572 17276 40628 17332
rect 38668 14140 38724 14196
rect 39676 16156 39732 16212
rect 39852 15706 39908 15708
rect 39852 15654 39854 15706
rect 39854 15654 39906 15706
rect 39906 15654 39908 15706
rect 39852 15652 39908 15654
rect 39956 15706 40012 15708
rect 39956 15654 39958 15706
rect 39958 15654 40010 15706
rect 40010 15654 40012 15706
rect 39956 15652 40012 15654
rect 40060 15706 40116 15708
rect 40060 15654 40062 15706
rect 40062 15654 40114 15706
rect 40114 15654 40116 15706
rect 40060 15652 40116 15654
rect 40012 15484 40068 15540
rect 38668 13916 38724 13972
rect 38444 13634 38500 13636
rect 38444 13582 38446 13634
rect 38446 13582 38498 13634
rect 38498 13582 38500 13634
rect 38444 13580 38500 13582
rect 38220 13132 38276 13188
rect 37660 10556 37716 10612
rect 38108 12572 38164 12628
rect 37212 8988 37268 9044
rect 37548 8652 37604 8708
rect 37212 8316 37268 8372
rect 37324 8428 37380 8484
rect 37100 8146 37156 8148
rect 37100 8094 37102 8146
rect 37102 8094 37154 8146
rect 37154 8094 37156 8146
rect 37100 8092 37156 8094
rect 35644 6300 35700 6356
rect 37436 7308 37492 7364
rect 36092 6748 36148 6804
rect 36204 6524 36260 6580
rect 35868 6188 35924 6244
rect 36204 6130 36260 6132
rect 36204 6078 36206 6130
rect 36206 6078 36258 6130
rect 36258 6078 36260 6130
rect 36204 6076 36260 6078
rect 37100 6130 37156 6132
rect 37100 6078 37102 6130
rect 37102 6078 37154 6130
rect 37154 6078 37156 6130
rect 37100 6076 37156 6078
rect 37436 6076 37492 6132
rect 35756 5964 35812 6020
rect 35644 5180 35700 5236
rect 35308 4172 35364 4228
rect 35644 4898 35700 4900
rect 35644 4846 35646 4898
rect 35646 4846 35698 4898
rect 35698 4846 35700 4898
rect 35644 4844 35700 4846
rect 32508 3442 32564 3444
rect 32508 3390 32510 3442
rect 32510 3390 32562 3442
rect 32562 3390 32564 3442
rect 32508 3388 32564 3390
rect 32284 2828 32340 2884
rect 36204 5292 36260 5348
rect 36652 5292 36708 5348
rect 36428 4060 36484 4116
rect 35420 2380 35476 2436
rect 37436 5234 37492 5236
rect 37436 5182 37438 5234
rect 37438 5182 37490 5234
rect 37490 5182 37492 5234
rect 37436 5180 37492 5182
rect 37100 5122 37156 5124
rect 37100 5070 37102 5122
rect 37102 5070 37154 5122
rect 37154 5070 37156 5122
rect 37100 5068 37156 5070
rect 37996 11340 38052 11396
rect 37884 11228 37940 11284
rect 38220 11228 38276 11284
rect 38668 11900 38724 11956
rect 38668 11676 38724 11732
rect 38668 10498 38724 10500
rect 38668 10446 38670 10498
rect 38670 10446 38722 10498
rect 38722 10446 38724 10498
rect 38668 10444 38724 10446
rect 38556 10332 38612 10388
rect 37884 9996 37940 10052
rect 37996 8652 38052 8708
rect 38332 8428 38388 8484
rect 38220 7868 38276 7924
rect 38108 6860 38164 6916
rect 37996 6130 38052 6132
rect 37996 6078 37998 6130
rect 37998 6078 38050 6130
rect 38050 6078 38052 6130
rect 37996 6076 38052 6078
rect 37772 4956 37828 5012
rect 38892 14306 38948 14308
rect 38892 14254 38894 14306
rect 38894 14254 38946 14306
rect 38946 14254 38948 14306
rect 38892 14252 38948 14254
rect 39228 13970 39284 13972
rect 39228 13918 39230 13970
rect 39230 13918 39282 13970
rect 39282 13918 39284 13970
rect 39228 13916 39284 13918
rect 39900 14530 39956 14532
rect 39900 14478 39902 14530
rect 39902 14478 39954 14530
rect 39954 14478 39956 14530
rect 39900 14476 39956 14478
rect 39852 14138 39908 14140
rect 39852 14086 39854 14138
rect 39854 14086 39906 14138
rect 39906 14086 39908 14138
rect 39852 14084 39908 14086
rect 39956 14138 40012 14140
rect 39956 14086 39958 14138
rect 39958 14086 40010 14138
rect 40010 14086 40012 14138
rect 39956 14084 40012 14086
rect 40060 14138 40116 14140
rect 40060 14086 40062 14138
rect 40062 14086 40114 14138
rect 40114 14086 40116 14138
rect 40060 14084 40116 14086
rect 40348 15202 40404 15204
rect 40348 15150 40350 15202
rect 40350 15150 40402 15202
rect 40402 15150 40404 15202
rect 40348 15148 40404 15150
rect 38444 6748 38500 6804
rect 38220 5122 38276 5124
rect 38220 5070 38222 5122
rect 38222 5070 38274 5122
rect 38274 5070 38276 5122
rect 38220 5068 38276 5070
rect 37660 4844 37716 4900
rect 38780 7868 38836 7924
rect 38780 7084 38836 7140
rect 39116 13074 39172 13076
rect 39116 13022 39118 13074
rect 39118 13022 39170 13074
rect 39170 13022 39172 13074
rect 39116 13020 39172 13022
rect 39340 13020 39396 13076
rect 39340 12572 39396 12628
rect 39452 12908 39508 12964
rect 40012 12684 40068 12740
rect 39852 12570 39908 12572
rect 39852 12518 39854 12570
rect 39854 12518 39906 12570
rect 39906 12518 39908 12570
rect 39852 12516 39908 12518
rect 39956 12570 40012 12572
rect 39956 12518 39958 12570
rect 39958 12518 40010 12570
rect 40010 12518 40012 12570
rect 39956 12516 40012 12518
rect 40060 12570 40116 12572
rect 40060 12518 40062 12570
rect 40062 12518 40114 12570
rect 40114 12518 40116 12570
rect 40060 12516 40116 12518
rect 39900 12348 39956 12404
rect 39004 12012 39060 12068
rect 39004 11506 39060 11508
rect 39004 11454 39006 11506
rect 39006 11454 39058 11506
rect 39058 11454 39060 11506
rect 39004 11452 39060 11454
rect 40124 11452 40180 11508
rect 40348 12236 40404 12292
rect 39340 11228 39396 11284
rect 39452 11004 39508 11060
rect 39852 11002 39908 11004
rect 39852 10950 39854 11002
rect 39854 10950 39906 11002
rect 39906 10950 39908 11002
rect 39852 10948 39908 10950
rect 39956 11002 40012 11004
rect 39956 10950 39958 11002
rect 39958 10950 40010 11002
rect 40010 10950 40012 11002
rect 39956 10948 40012 10950
rect 40060 11002 40116 11004
rect 40060 10950 40062 11002
rect 40062 10950 40114 11002
rect 40114 10950 40116 11002
rect 40060 10948 40116 10950
rect 39340 10668 39396 10724
rect 40012 10722 40068 10724
rect 40012 10670 40014 10722
rect 40014 10670 40066 10722
rect 40066 10670 40068 10722
rect 40012 10668 40068 10670
rect 39676 10444 39732 10500
rect 39852 9434 39908 9436
rect 39852 9382 39854 9434
rect 39854 9382 39906 9434
rect 39906 9382 39908 9434
rect 39852 9380 39908 9382
rect 39956 9434 40012 9436
rect 39956 9382 39958 9434
rect 39958 9382 40010 9434
rect 40010 9382 40012 9434
rect 39956 9380 40012 9382
rect 40060 9434 40116 9436
rect 40060 9382 40062 9434
rect 40062 9382 40114 9434
rect 40114 9382 40116 9434
rect 40060 9380 40116 9382
rect 39452 7474 39508 7476
rect 39452 7422 39454 7474
rect 39454 7422 39506 7474
rect 39506 7422 39508 7474
rect 39452 7420 39508 7422
rect 40796 16940 40852 16996
rect 41020 18060 41076 18116
rect 41244 17948 41300 18004
rect 41020 17276 41076 17332
rect 41020 16994 41076 16996
rect 41020 16942 41022 16994
rect 41022 16942 41074 16994
rect 41074 16942 41076 16994
rect 41020 16940 41076 16942
rect 40460 8092 40516 8148
rect 40684 16268 40740 16324
rect 41020 15820 41076 15876
rect 41580 19010 41636 19012
rect 41580 18958 41582 19010
rect 41582 18958 41634 19010
rect 41634 18958 41636 19010
rect 41580 18956 41636 18958
rect 42028 19740 42084 19796
rect 41692 19292 41748 19348
rect 41468 18396 41524 18452
rect 41020 14530 41076 14532
rect 41020 14478 41022 14530
rect 41022 14478 41074 14530
rect 41074 14478 41076 14530
rect 41020 14476 41076 14478
rect 39852 7866 39908 7868
rect 39852 7814 39854 7866
rect 39854 7814 39906 7866
rect 39906 7814 39908 7866
rect 39852 7812 39908 7814
rect 39956 7866 40012 7868
rect 39956 7814 39958 7866
rect 39958 7814 40010 7866
rect 40010 7814 40012 7866
rect 39956 7812 40012 7814
rect 40060 7866 40116 7868
rect 40060 7814 40062 7866
rect 40062 7814 40114 7866
rect 40114 7814 40116 7866
rect 40060 7812 40116 7814
rect 40124 7586 40180 7588
rect 40124 7534 40126 7586
rect 40126 7534 40178 7586
rect 40178 7534 40180 7586
rect 40124 7532 40180 7534
rect 40684 14364 40740 14420
rect 40236 6972 40292 7028
rect 38892 6636 38948 6692
rect 39852 6298 39908 6300
rect 39852 6246 39854 6298
rect 39854 6246 39906 6298
rect 39906 6246 39908 6298
rect 39852 6244 39908 6246
rect 39956 6298 40012 6300
rect 39956 6246 39958 6298
rect 39958 6246 40010 6298
rect 40010 6246 40012 6298
rect 39956 6244 40012 6246
rect 40060 6298 40116 6300
rect 40060 6246 40062 6298
rect 40062 6246 40114 6298
rect 40114 6246 40116 6298
rect 40060 6244 40116 6246
rect 39004 5852 39060 5908
rect 38668 5068 38724 5124
rect 40908 13858 40964 13860
rect 40908 13806 40910 13858
rect 40910 13806 40962 13858
rect 40962 13806 40964 13858
rect 40908 13804 40964 13806
rect 42028 18450 42084 18452
rect 42028 18398 42030 18450
rect 42030 18398 42082 18450
rect 42082 18398 42084 18450
rect 42028 18396 42084 18398
rect 42700 26514 42756 26516
rect 42700 26462 42702 26514
rect 42702 26462 42754 26514
rect 42754 26462 42756 26514
rect 42700 26460 42756 26462
rect 43484 27074 43540 27076
rect 43484 27022 43486 27074
rect 43486 27022 43538 27074
rect 43538 27022 43540 27074
rect 43484 27020 43540 27022
rect 43372 26962 43428 26964
rect 43372 26910 43374 26962
rect 43374 26910 43426 26962
rect 43426 26910 43428 26962
rect 43372 26908 43428 26910
rect 42476 24722 42532 24724
rect 42476 24670 42478 24722
rect 42478 24670 42530 24722
rect 42530 24670 42532 24722
rect 42476 24668 42532 24670
rect 42700 24220 42756 24276
rect 42588 24108 42644 24164
rect 43372 25900 43428 25956
rect 43484 25564 43540 25620
rect 43932 29372 43988 29428
rect 43932 28082 43988 28084
rect 43932 28030 43934 28082
rect 43934 28030 43986 28082
rect 43986 28030 43988 28082
rect 43932 28028 43988 28030
rect 44268 29260 44324 29316
rect 45836 36428 45892 36484
rect 44940 35026 44996 35028
rect 44940 34974 44942 35026
rect 44942 34974 44994 35026
rect 44994 34974 44996 35026
rect 44940 34972 44996 34974
rect 45164 35420 45220 35476
rect 45164 34636 45220 34692
rect 44716 34242 44772 34244
rect 44716 34190 44718 34242
rect 44718 34190 44770 34242
rect 44770 34190 44772 34242
rect 44716 34188 44772 34190
rect 44828 33458 44884 33460
rect 44828 33406 44830 33458
rect 44830 33406 44882 33458
rect 44882 33406 44884 33458
rect 44828 33404 44884 33406
rect 44604 31106 44660 31108
rect 44604 31054 44606 31106
rect 44606 31054 44658 31106
rect 44658 31054 44660 31106
rect 44604 31052 44660 31054
rect 45388 35026 45444 35028
rect 45388 34974 45390 35026
rect 45390 34974 45442 35026
rect 45442 34974 45444 35026
rect 45388 34972 45444 34974
rect 45388 33458 45444 33460
rect 45388 33406 45390 33458
rect 45390 33406 45442 33458
rect 45442 33406 45444 33458
rect 45388 33404 45444 33406
rect 45276 32732 45332 32788
rect 44828 32396 44884 32452
rect 45164 32396 45220 32452
rect 45612 35196 45668 35252
rect 45724 34972 45780 35028
rect 45612 34748 45668 34804
rect 46284 36204 46340 36260
rect 46284 35868 46340 35924
rect 46844 35868 46900 35924
rect 48188 35810 48244 35812
rect 48188 35758 48190 35810
rect 48190 35758 48242 35810
rect 48242 35758 48244 35810
rect 48188 35756 48244 35758
rect 45948 34914 46004 34916
rect 45948 34862 45950 34914
rect 45950 34862 46002 34914
rect 46002 34862 46004 34914
rect 45948 34860 46004 34862
rect 45836 34748 45892 34804
rect 47628 35698 47684 35700
rect 47628 35646 47630 35698
rect 47630 35646 47682 35698
rect 47682 35646 47684 35698
rect 47628 35644 47684 35646
rect 46172 35308 46228 35364
rect 45724 34300 45780 34356
rect 45836 34242 45892 34244
rect 45836 34190 45838 34242
rect 45838 34190 45890 34242
rect 45890 34190 45892 34242
rect 45836 34188 45892 34190
rect 45836 33346 45892 33348
rect 45836 33294 45838 33346
rect 45838 33294 45890 33346
rect 45890 33294 45892 33346
rect 45836 33292 45892 33294
rect 45612 32786 45668 32788
rect 45612 32734 45614 32786
rect 45614 32734 45666 32786
rect 45666 32734 45668 32786
rect 45612 32732 45668 32734
rect 46396 35026 46452 35028
rect 46396 34974 46398 35026
rect 46398 34974 46450 35026
rect 46450 34974 46452 35026
rect 46396 34972 46452 34974
rect 46732 34860 46788 34916
rect 47628 34972 47684 35028
rect 46284 32786 46340 32788
rect 46284 32734 46286 32786
rect 46286 32734 46338 32786
rect 46338 32734 46340 32786
rect 46284 32732 46340 32734
rect 45052 31612 45108 31668
rect 44940 31500 44996 31556
rect 44940 29820 44996 29876
rect 44716 29426 44772 29428
rect 44716 29374 44718 29426
rect 44718 29374 44770 29426
rect 44770 29374 44772 29426
rect 44716 29372 44772 29374
rect 44940 29148 44996 29204
rect 44940 28700 44996 28756
rect 44380 28082 44436 28084
rect 44380 28030 44382 28082
rect 44382 28030 44434 28082
rect 44434 28030 44436 28082
rect 44380 28028 44436 28030
rect 44492 27692 44548 27748
rect 44492 27356 44548 27412
rect 43932 26124 43988 26180
rect 43820 25900 43876 25956
rect 44268 25452 44324 25508
rect 43036 24668 43092 24724
rect 43260 24220 43316 24276
rect 43036 23884 43092 23940
rect 43372 23548 43428 23604
rect 42476 23212 42532 23268
rect 42812 23378 42868 23380
rect 42812 23326 42814 23378
rect 42814 23326 42866 23378
rect 42866 23326 42868 23378
rect 42812 23324 42868 23326
rect 43372 22540 43428 22596
rect 43260 22370 43316 22372
rect 43260 22318 43262 22370
rect 43262 22318 43314 22370
rect 43314 22318 43316 22370
rect 43260 22316 43316 22318
rect 42364 21810 42420 21812
rect 42364 21758 42366 21810
rect 42366 21758 42418 21810
rect 42418 21758 42420 21810
rect 42364 21756 42420 21758
rect 42812 21586 42868 21588
rect 42812 21534 42814 21586
rect 42814 21534 42866 21586
rect 42866 21534 42868 21586
rect 42812 21532 42868 21534
rect 43372 21586 43428 21588
rect 43372 21534 43374 21586
rect 43374 21534 43426 21586
rect 43426 21534 43428 21586
rect 43372 21532 43428 21534
rect 43708 23938 43764 23940
rect 43708 23886 43710 23938
rect 43710 23886 43762 23938
rect 43762 23886 43764 23938
rect 43708 23884 43764 23886
rect 43596 23826 43652 23828
rect 43596 23774 43598 23826
rect 43598 23774 43650 23826
rect 43650 23774 43652 23826
rect 43596 23772 43652 23774
rect 43820 23042 43876 23044
rect 43820 22990 43822 23042
rect 43822 22990 43874 23042
rect 43874 22990 43876 23042
rect 43820 22988 43876 22990
rect 43708 22146 43764 22148
rect 43708 22094 43710 22146
rect 43710 22094 43762 22146
rect 43762 22094 43764 22146
rect 43708 22092 43764 22094
rect 42700 20972 42756 21028
rect 44156 25116 44212 25172
rect 44044 24610 44100 24612
rect 44044 24558 44046 24610
rect 44046 24558 44098 24610
rect 44098 24558 44100 24610
rect 44044 24556 44100 24558
rect 44044 23996 44100 24052
rect 44156 23548 44212 23604
rect 44828 26962 44884 26964
rect 44828 26910 44830 26962
rect 44830 26910 44882 26962
rect 44882 26910 44884 26962
rect 44828 26908 44884 26910
rect 44828 26684 44884 26740
rect 46172 31890 46228 31892
rect 46172 31838 46174 31890
rect 46174 31838 46226 31890
rect 46226 31838 46228 31890
rect 46172 31836 46228 31838
rect 45388 31554 45444 31556
rect 45388 31502 45390 31554
rect 45390 31502 45442 31554
rect 45442 31502 45444 31554
rect 45388 31500 45444 31502
rect 45388 31164 45444 31220
rect 45724 29820 45780 29876
rect 46060 29932 46116 29988
rect 45276 29484 45332 29540
rect 45948 29314 46004 29316
rect 45948 29262 45950 29314
rect 45950 29262 46002 29314
rect 46002 29262 46004 29314
rect 45948 29260 46004 29262
rect 46172 29538 46228 29540
rect 46172 29486 46174 29538
rect 46174 29486 46226 29538
rect 46226 29486 46228 29538
rect 46172 29484 46228 29486
rect 45164 27356 45220 27412
rect 45388 27746 45444 27748
rect 45388 27694 45390 27746
rect 45390 27694 45442 27746
rect 45442 27694 45444 27746
rect 45388 27692 45444 27694
rect 45500 26962 45556 26964
rect 45500 26910 45502 26962
rect 45502 26910 45554 26962
rect 45554 26910 45556 26962
rect 45500 26908 45556 26910
rect 45836 26962 45892 26964
rect 45836 26910 45838 26962
rect 45838 26910 45890 26962
rect 45890 26910 45892 26962
rect 45836 26908 45892 26910
rect 46172 27916 46228 27972
rect 46620 31724 46676 31780
rect 46732 31554 46788 31556
rect 46732 31502 46734 31554
rect 46734 31502 46786 31554
rect 46786 31502 46788 31554
rect 46732 31500 46788 31502
rect 47964 35420 48020 35476
rect 49512 36874 49568 36876
rect 49512 36822 49514 36874
rect 49514 36822 49566 36874
rect 49566 36822 49568 36874
rect 49512 36820 49568 36822
rect 49616 36874 49672 36876
rect 49616 36822 49618 36874
rect 49618 36822 49670 36874
rect 49670 36822 49672 36874
rect 49616 36820 49672 36822
rect 49720 36874 49776 36876
rect 49720 36822 49722 36874
rect 49722 36822 49774 36874
rect 49774 36822 49776 36874
rect 49720 36820 49776 36822
rect 48972 35810 49028 35812
rect 48972 35758 48974 35810
rect 48974 35758 49026 35810
rect 49026 35758 49028 35810
rect 48972 35756 49028 35758
rect 49084 35698 49140 35700
rect 49084 35646 49086 35698
rect 49086 35646 49138 35698
rect 49138 35646 49140 35698
rect 49084 35644 49140 35646
rect 48860 35420 48916 35476
rect 48412 35084 48468 35140
rect 49196 34636 49252 34692
rect 48076 34412 48132 34468
rect 47740 33516 47796 33572
rect 48524 31948 48580 32004
rect 47964 31836 48020 31892
rect 47516 31500 47572 31556
rect 46844 30940 46900 30996
rect 47964 30882 48020 30884
rect 47964 30830 47966 30882
rect 47966 30830 48018 30882
rect 48018 30830 48020 30882
rect 47964 30828 48020 30830
rect 46396 28588 46452 28644
rect 46284 27580 46340 27636
rect 46732 29372 46788 29428
rect 46956 29986 47012 29988
rect 46956 29934 46958 29986
rect 46958 29934 47010 29986
rect 47010 29934 47012 29986
rect 46956 29932 47012 29934
rect 46956 29260 47012 29316
rect 46844 28700 46900 28756
rect 46956 28924 47012 28980
rect 46956 28028 47012 28084
rect 46956 27580 47012 27636
rect 45052 25900 45108 25956
rect 44940 25788 44996 25844
rect 44828 25506 44884 25508
rect 44828 25454 44830 25506
rect 44830 25454 44882 25506
rect 44882 25454 44884 25506
rect 44828 25452 44884 25454
rect 46844 27020 46900 27076
rect 45724 26066 45780 26068
rect 45724 26014 45726 26066
rect 45726 26014 45778 26066
rect 45778 26014 45780 26066
rect 45724 26012 45780 26014
rect 45612 25788 45668 25844
rect 45948 25228 46004 25284
rect 44716 24556 44772 24612
rect 45276 24722 45332 24724
rect 45276 24670 45278 24722
rect 45278 24670 45330 24722
rect 45330 24670 45332 24722
rect 45276 24668 45332 24670
rect 44380 23324 44436 23380
rect 43932 21532 43988 21588
rect 43036 20524 43092 20580
rect 43932 20578 43988 20580
rect 43932 20526 43934 20578
rect 43934 20526 43986 20578
rect 43986 20526 43988 20578
rect 43932 20524 43988 20526
rect 42476 20130 42532 20132
rect 42476 20078 42478 20130
rect 42478 20078 42530 20130
rect 42530 20078 42532 20130
rect 42476 20076 42532 20078
rect 42700 20130 42756 20132
rect 42700 20078 42702 20130
rect 42702 20078 42754 20130
rect 42754 20078 42756 20130
rect 42700 20076 42756 20078
rect 42364 19516 42420 19572
rect 42252 19180 42308 19236
rect 42476 18956 42532 19012
rect 42476 17164 42532 17220
rect 42588 16940 42644 16996
rect 41804 16716 41860 16772
rect 42364 16882 42420 16884
rect 42364 16830 42366 16882
rect 42366 16830 42418 16882
rect 42418 16830 42420 16882
rect 42364 16828 42420 16830
rect 42700 18172 42756 18228
rect 43260 20130 43316 20132
rect 43260 20078 43262 20130
rect 43262 20078 43314 20130
rect 43314 20078 43316 20130
rect 43260 20076 43316 20078
rect 43708 19740 43764 19796
rect 43932 19068 43988 19124
rect 43036 18284 43092 18340
rect 42924 17500 42980 17556
rect 42812 16044 42868 16100
rect 42924 17164 42980 17220
rect 43484 18284 43540 18340
rect 44044 18396 44100 18452
rect 43596 17500 43652 17556
rect 43260 17164 43316 17220
rect 43372 17388 43428 17444
rect 43148 16940 43204 16996
rect 42364 15932 42420 15988
rect 42028 15484 42084 15540
rect 41692 14364 41748 14420
rect 41916 14476 41972 14532
rect 41580 14252 41636 14308
rect 41244 13916 41300 13972
rect 40796 11506 40852 11508
rect 40796 11454 40798 11506
rect 40798 11454 40850 11506
rect 40850 11454 40852 11506
rect 40796 11452 40852 11454
rect 40796 10892 40852 10948
rect 41692 13858 41748 13860
rect 41692 13806 41694 13858
rect 41694 13806 41746 13858
rect 41746 13806 41748 13858
rect 41692 13804 41748 13806
rect 41468 13468 41524 13524
rect 41692 13244 41748 13300
rect 41356 12796 41412 12852
rect 41132 12684 41188 12740
rect 43036 15820 43092 15876
rect 42924 15708 42980 15764
rect 42812 15484 42868 15540
rect 42700 15426 42756 15428
rect 42700 15374 42702 15426
rect 42702 15374 42754 15426
rect 42754 15374 42756 15426
rect 42700 15372 42756 15374
rect 43596 16882 43652 16884
rect 43596 16830 43598 16882
rect 43598 16830 43650 16882
rect 43650 16830 43652 16882
rect 43596 16828 43652 16830
rect 43484 16098 43540 16100
rect 43484 16046 43486 16098
rect 43486 16046 43538 16098
rect 43538 16046 43540 16098
rect 43484 16044 43540 16046
rect 43484 15708 43540 15764
rect 43708 15484 43764 15540
rect 43820 16940 43876 16996
rect 43932 16828 43988 16884
rect 44044 17164 44100 17220
rect 43372 15260 43428 15316
rect 43932 16492 43988 16548
rect 43932 16044 43988 16100
rect 44268 21308 44324 21364
rect 44492 21420 44548 21476
rect 44492 19516 44548 19572
rect 44268 17554 44324 17556
rect 44268 17502 44270 17554
rect 44270 17502 44322 17554
rect 44322 17502 44324 17554
rect 44268 17500 44324 17502
rect 44380 17442 44436 17444
rect 44380 17390 44382 17442
rect 44382 17390 44434 17442
rect 44434 17390 44436 17442
rect 44380 17388 44436 17390
rect 44156 16882 44212 16884
rect 44156 16830 44158 16882
rect 44158 16830 44210 16882
rect 44210 16830 44212 16882
rect 44156 16828 44212 16830
rect 44156 15708 44212 15764
rect 43932 15596 43988 15652
rect 42364 13804 42420 13860
rect 42140 13356 42196 13412
rect 42252 13132 42308 13188
rect 42364 12962 42420 12964
rect 42364 12910 42366 12962
rect 42366 12910 42418 12962
rect 42418 12910 42420 12962
rect 42364 12908 42420 12910
rect 42588 13916 42644 13972
rect 42588 13356 42644 13412
rect 41804 12290 41860 12292
rect 41804 12238 41806 12290
rect 41806 12238 41858 12290
rect 41858 12238 41860 12290
rect 41804 12236 41860 12238
rect 41692 12012 41748 12068
rect 41132 11228 41188 11284
rect 42140 11506 42196 11508
rect 42140 11454 42142 11506
rect 42142 11454 42194 11506
rect 42194 11454 42196 11506
rect 42140 11452 42196 11454
rect 41804 11282 41860 11284
rect 41804 11230 41806 11282
rect 41806 11230 41858 11282
rect 41858 11230 41860 11282
rect 41804 11228 41860 11230
rect 41356 11170 41412 11172
rect 41356 11118 41358 11170
rect 41358 11118 41410 11170
rect 41410 11118 41412 11170
rect 41356 11116 41412 11118
rect 41356 10892 41412 10948
rect 42364 12402 42420 12404
rect 42364 12350 42366 12402
rect 42366 12350 42418 12402
rect 42418 12350 42420 12402
rect 42364 12348 42420 12350
rect 42364 11676 42420 11732
rect 41580 10386 41636 10388
rect 41580 10334 41582 10386
rect 41582 10334 41634 10386
rect 41634 10334 41636 10386
rect 41580 10332 41636 10334
rect 40908 8204 40964 8260
rect 40796 7532 40852 7588
rect 41468 7420 41524 7476
rect 41468 6972 41524 7028
rect 41916 7532 41972 7588
rect 42028 6972 42084 7028
rect 39852 4730 39908 4732
rect 39852 4678 39854 4730
rect 39854 4678 39906 4730
rect 39906 4678 39908 4730
rect 39852 4676 39908 4678
rect 39956 4730 40012 4732
rect 39956 4678 39958 4730
rect 39958 4678 40010 4730
rect 40010 4678 40012 4730
rect 39956 4676 40012 4678
rect 40060 4730 40116 4732
rect 40060 4678 40062 4730
rect 40062 4678 40114 4730
rect 40114 4678 40116 4730
rect 40060 4676 40116 4678
rect 38668 4396 38724 4452
rect 40460 4732 40516 4788
rect 40348 4338 40404 4340
rect 40348 4286 40350 4338
rect 40350 4286 40402 4338
rect 40402 4286 40404 4338
rect 40348 4284 40404 4286
rect 40236 3948 40292 4004
rect 38556 3724 38612 3780
rect 41020 4338 41076 4340
rect 41020 4286 41022 4338
rect 41022 4286 41074 4338
rect 41074 4286 41076 4338
rect 41020 4284 41076 4286
rect 42476 11116 42532 11172
rect 42588 10892 42644 10948
rect 42364 10332 42420 10388
rect 42364 8092 42420 8148
rect 43036 13970 43092 13972
rect 43036 13918 43038 13970
rect 43038 13918 43090 13970
rect 43090 13918 43092 13970
rect 43036 13916 43092 13918
rect 42924 13746 42980 13748
rect 42924 13694 42926 13746
rect 42926 13694 42978 13746
rect 42978 13694 42980 13746
rect 42924 13692 42980 13694
rect 42812 13468 42868 13524
rect 43260 13858 43316 13860
rect 43260 13806 43262 13858
rect 43262 13806 43314 13858
rect 43314 13806 43316 13858
rect 43260 13804 43316 13806
rect 43820 13746 43876 13748
rect 43820 13694 43822 13746
rect 43822 13694 43874 13746
rect 43874 13694 43876 13746
rect 43820 13692 43876 13694
rect 44156 15538 44212 15540
rect 44156 15486 44158 15538
rect 44158 15486 44210 15538
rect 44210 15486 44212 15538
rect 44156 15484 44212 15486
rect 44044 15314 44100 15316
rect 44044 15262 44046 15314
rect 44046 15262 44098 15314
rect 44098 15262 44100 15314
rect 44044 15260 44100 15262
rect 44380 16770 44436 16772
rect 44380 16718 44382 16770
rect 44382 16718 44434 16770
rect 44434 16718 44436 16770
rect 44380 16716 44436 16718
rect 44380 15820 44436 15876
rect 44492 15596 44548 15652
rect 44268 13244 44324 13300
rect 42812 12012 42868 12068
rect 42812 11170 42868 11172
rect 42812 11118 42814 11170
rect 42814 11118 42866 11170
rect 42866 11118 42868 11170
rect 42812 11116 42868 11118
rect 44156 12908 44212 12964
rect 43484 12178 43540 12180
rect 43484 12126 43486 12178
rect 43486 12126 43538 12178
rect 43538 12126 43540 12178
rect 43484 12124 43540 12126
rect 43036 11900 43092 11956
rect 43148 11452 43204 11508
rect 43932 12066 43988 12068
rect 43932 12014 43934 12066
rect 43934 12014 43986 12066
rect 43986 12014 43988 12066
rect 43932 12012 43988 12014
rect 43484 11340 43540 11396
rect 43820 11394 43876 11396
rect 43820 11342 43822 11394
rect 43822 11342 43874 11394
rect 43874 11342 43876 11394
rect 43820 11340 43876 11342
rect 43148 10610 43204 10612
rect 43148 10558 43150 10610
rect 43150 10558 43202 10610
rect 43202 10558 43204 10610
rect 43148 10556 43204 10558
rect 43036 9996 43092 10052
rect 43260 9996 43316 10052
rect 43036 9436 43092 9492
rect 42812 9100 42868 9156
rect 42588 8316 42644 8372
rect 42588 7586 42644 7588
rect 42588 7534 42590 7586
rect 42590 7534 42642 7586
rect 42642 7534 42644 7586
rect 42588 7532 42644 7534
rect 42476 7196 42532 7252
rect 42364 4956 42420 5012
rect 42028 4338 42084 4340
rect 42028 4286 42030 4338
rect 42030 4286 42082 4338
rect 42082 4286 42084 4338
rect 42028 4284 42084 4286
rect 41916 4060 41972 4116
rect 42924 6972 42980 7028
rect 43260 7250 43316 7252
rect 43260 7198 43262 7250
rect 43262 7198 43314 7250
rect 43314 7198 43316 7250
rect 43260 7196 43316 7198
rect 43820 10610 43876 10612
rect 43820 10558 43822 10610
rect 43822 10558 43874 10610
rect 43874 10558 43876 10610
rect 43820 10556 43876 10558
rect 43484 10332 43540 10388
rect 44268 10498 44324 10500
rect 44268 10446 44270 10498
rect 44270 10446 44322 10498
rect 44322 10446 44324 10498
rect 44268 10444 44324 10446
rect 43484 8988 43540 9044
rect 45164 22652 45220 22708
rect 45388 24556 45444 24612
rect 45836 24556 45892 24612
rect 46172 24722 46228 24724
rect 46172 24670 46174 24722
rect 46174 24670 46226 24722
rect 46226 24670 46228 24722
rect 46172 24668 46228 24670
rect 46284 26012 46340 26068
rect 46620 24946 46676 24948
rect 46620 24894 46622 24946
rect 46622 24894 46674 24946
rect 46674 24894 46676 24946
rect 46620 24892 46676 24894
rect 48076 30210 48132 30212
rect 48076 30158 48078 30210
rect 48078 30158 48130 30210
rect 48130 30158 48132 30210
rect 48076 30156 48132 30158
rect 47180 29484 47236 29540
rect 47292 28700 47348 28756
rect 47740 29986 47796 29988
rect 47740 29934 47742 29986
rect 47742 29934 47794 29986
rect 47794 29934 47796 29986
rect 47740 29932 47796 29934
rect 47740 29484 47796 29540
rect 47852 29372 47908 29428
rect 47852 28642 47908 28644
rect 47852 28590 47854 28642
rect 47854 28590 47906 28642
rect 47906 28590 47908 28642
rect 47852 28588 47908 28590
rect 48412 29596 48468 29652
rect 48300 29484 48356 29540
rect 48636 31554 48692 31556
rect 48636 31502 48638 31554
rect 48638 31502 48690 31554
rect 48690 31502 48692 31554
rect 48636 31500 48692 31502
rect 49512 35306 49568 35308
rect 49512 35254 49514 35306
rect 49514 35254 49566 35306
rect 49566 35254 49568 35306
rect 49512 35252 49568 35254
rect 49616 35306 49672 35308
rect 49616 35254 49618 35306
rect 49618 35254 49670 35306
rect 49670 35254 49672 35306
rect 49616 35252 49672 35254
rect 49720 35306 49776 35308
rect 49720 35254 49722 35306
rect 49722 35254 49774 35306
rect 49774 35254 49776 35306
rect 49720 35252 49776 35254
rect 49420 34412 49476 34468
rect 50428 36258 50484 36260
rect 50428 36206 50430 36258
rect 50430 36206 50482 36258
rect 50482 36206 50484 36258
rect 50428 36204 50484 36206
rect 50428 35698 50484 35700
rect 50428 35646 50430 35698
rect 50430 35646 50482 35698
rect 50482 35646 50484 35698
rect 50428 35644 50484 35646
rect 49868 34076 49924 34132
rect 48860 33570 48916 33572
rect 48860 33518 48862 33570
rect 48862 33518 48914 33570
rect 48914 33518 48916 33570
rect 48860 33516 48916 33518
rect 49512 33738 49568 33740
rect 49512 33686 49514 33738
rect 49514 33686 49566 33738
rect 49566 33686 49568 33738
rect 49512 33684 49568 33686
rect 49616 33738 49672 33740
rect 49616 33686 49618 33738
rect 49618 33686 49670 33738
rect 49670 33686 49672 33738
rect 49616 33684 49672 33686
rect 49720 33738 49776 33740
rect 49720 33686 49722 33738
rect 49722 33686 49774 33738
rect 49774 33686 49776 33738
rect 49720 33684 49776 33686
rect 49196 33346 49252 33348
rect 49196 33294 49198 33346
rect 49198 33294 49250 33346
rect 49250 33294 49252 33346
rect 49196 33292 49252 33294
rect 49868 33068 49924 33124
rect 49512 32170 49568 32172
rect 49512 32118 49514 32170
rect 49514 32118 49566 32170
rect 49566 32118 49568 32170
rect 49512 32116 49568 32118
rect 49616 32170 49672 32172
rect 49616 32118 49618 32170
rect 49618 32118 49670 32170
rect 49670 32118 49672 32170
rect 49616 32116 49672 32118
rect 49720 32170 49776 32172
rect 49720 32118 49722 32170
rect 49722 32118 49774 32170
rect 49774 32118 49776 32170
rect 49720 32116 49776 32118
rect 48972 31836 49028 31892
rect 49644 31666 49700 31668
rect 49644 31614 49646 31666
rect 49646 31614 49698 31666
rect 49698 31614 49700 31666
rect 49644 31612 49700 31614
rect 48972 31554 49028 31556
rect 48972 31502 48974 31554
rect 48974 31502 49026 31554
rect 49026 31502 49028 31554
rect 48972 31500 49028 31502
rect 49420 31500 49476 31556
rect 50652 35196 50708 35252
rect 50652 34636 50708 34692
rect 52556 37100 52612 37156
rect 52444 36652 52500 36708
rect 52332 36428 52388 36484
rect 50988 35698 51044 35700
rect 50988 35646 50990 35698
rect 50990 35646 51042 35698
rect 51042 35646 51044 35698
rect 50988 35644 51044 35646
rect 51324 35196 51380 35252
rect 51548 34972 51604 35028
rect 50540 33180 50596 33236
rect 50652 33068 50708 33124
rect 50092 31836 50148 31892
rect 48748 30156 48804 30212
rect 48972 31106 49028 31108
rect 48972 31054 48974 31106
rect 48974 31054 49026 31106
rect 49026 31054 49028 31106
rect 48972 31052 49028 31054
rect 48636 29426 48692 29428
rect 48636 29374 48638 29426
rect 48638 29374 48690 29426
rect 48690 29374 48692 29426
rect 48636 29372 48692 29374
rect 49308 31106 49364 31108
rect 49308 31054 49310 31106
rect 49310 31054 49362 31106
rect 49362 31054 49364 31106
rect 49308 31052 49364 31054
rect 49512 30602 49568 30604
rect 49512 30550 49514 30602
rect 49514 30550 49566 30602
rect 49566 30550 49568 30602
rect 49512 30548 49568 30550
rect 49616 30602 49672 30604
rect 49616 30550 49618 30602
rect 49618 30550 49670 30602
rect 49670 30550 49672 30602
rect 49616 30548 49672 30550
rect 49720 30602 49776 30604
rect 49720 30550 49722 30602
rect 49722 30550 49774 30602
rect 49774 30550 49776 30602
rect 49720 30548 49776 30550
rect 48972 30156 49028 30212
rect 49084 29650 49140 29652
rect 49084 29598 49086 29650
rect 49086 29598 49138 29650
rect 49138 29598 49140 29650
rect 49084 29596 49140 29598
rect 49868 29596 49924 29652
rect 49756 29538 49812 29540
rect 49756 29486 49758 29538
rect 49758 29486 49810 29538
rect 49810 29486 49812 29538
rect 49756 29484 49812 29486
rect 49756 29202 49812 29204
rect 49756 29150 49758 29202
rect 49758 29150 49810 29202
rect 49810 29150 49812 29202
rect 49756 29148 49812 29150
rect 48860 28700 48916 28756
rect 48524 28476 48580 28532
rect 47404 27916 47460 27972
rect 46956 24668 47012 24724
rect 45612 23436 45668 23492
rect 45388 23324 45444 23380
rect 45500 23042 45556 23044
rect 45500 22990 45502 23042
rect 45502 22990 45554 23042
rect 45554 22990 45556 23042
rect 45500 22988 45556 22990
rect 46172 23378 46228 23380
rect 46172 23326 46174 23378
rect 46174 23326 46226 23378
rect 46226 23326 46228 23378
rect 46172 23324 46228 23326
rect 47292 26796 47348 26852
rect 47852 26684 47908 26740
rect 48412 26850 48468 26852
rect 48412 26798 48414 26850
rect 48414 26798 48466 26850
rect 48466 26798 48468 26850
rect 48412 26796 48468 26798
rect 47292 26572 47348 26628
rect 48188 26178 48244 26180
rect 48188 26126 48190 26178
rect 48190 26126 48242 26178
rect 48242 26126 48244 26178
rect 48188 26124 48244 26126
rect 47516 25676 47572 25732
rect 48412 26012 48468 26068
rect 47852 25676 47908 25732
rect 48972 28476 49028 28532
rect 49512 29034 49568 29036
rect 49512 28982 49514 29034
rect 49514 28982 49566 29034
rect 49566 28982 49568 29034
rect 49512 28980 49568 28982
rect 49616 29034 49672 29036
rect 49616 28982 49618 29034
rect 49618 28982 49670 29034
rect 49670 28982 49672 29034
rect 49616 28980 49672 28982
rect 49720 29034 49776 29036
rect 49720 28982 49722 29034
rect 49722 28982 49774 29034
rect 49774 28982 49776 29034
rect 49720 28980 49776 28982
rect 49756 28082 49812 28084
rect 49756 28030 49758 28082
rect 49758 28030 49810 28082
rect 49810 28030 49812 28082
rect 49756 28028 49812 28030
rect 49512 27466 49568 27468
rect 49512 27414 49514 27466
rect 49514 27414 49566 27466
rect 49566 27414 49568 27466
rect 49512 27412 49568 27414
rect 49616 27466 49672 27468
rect 49616 27414 49618 27466
rect 49618 27414 49670 27466
rect 49670 27414 49672 27466
rect 49616 27412 49672 27414
rect 49720 27466 49776 27468
rect 49720 27414 49722 27466
rect 49722 27414 49774 27466
rect 49774 27414 49776 27466
rect 49720 27412 49776 27414
rect 49980 28754 50036 28756
rect 49980 28702 49982 28754
rect 49982 28702 50034 28754
rect 50034 28702 50036 28754
rect 49980 28700 50036 28702
rect 49980 28082 50036 28084
rect 49980 28030 49982 28082
rect 49982 28030 50034 28082
rect 50034 28030 50036 28082
rect 49980 28028 50036 28030
rect 49196 26796 49252 26852
rect 49532 26684 49588 26740
rect 49084 26124 49140 26180
rect 47740 25228 47796 25284
rect 48636 24892 48692 24948
rect 47516 23548 47572 23604
rect 47516 23378 47572 23380
rect 47516 23326 47518 23378
rect 47518 23326 47570 23378
rect 47570 23326 47572 23378
rect 47516 23324 47572 23326
rect 47180 23212 47236 23268
rect 45948 22988 46004 23044
rect 46172 22652 46228 22708
rect 46620 22482 46676 22484
rect 46620 22430 46622 22482
rect 46622 22430 46674 22482
rect 46674 22430 46676 22482
rect 46620 22428 46676 22430
rect 44940 22146 44996 22148
rect 44940 22094 44942 22146
rect 44942 22094 44994 22146
rect 44994 22094 44996 22146
rect 44940 22092 44996 22094
rect 44828 21532 44884 21588
rect 44940 21084 44996 21140
rect 47068 22764 47124 22820
rect 46732 22092 46788 22148
rect 45612 21586 45668 21588
rect 45612 21534 45614 21586
rect 45614 21534 45666 21586
rect 45666 21534 45668 21586
rect 45612 21532 45668 21534
rect 45500 21474 45556 21476
rect 45500 21422 45502 21474
rect 45502 21422 45554 21474
rect 45554 21422 45556 21474
rect 45500 21420 45556 21422
rect 45388 21308 45444 21364
rect 45948 21362 46004 21364
rect 45948 21310 45950 21362
rect 45950 21310 46002 21362
rect 46002 21310 46004 21362
rect 45948 21308 46004 21310
rect 45500 21084 45556 21140
rect 45164 20524 45220 20580
rect 44940 19122 44996 19124
rect 44940 19070 44942 19122
rect 44942 19070 44994 19122
rect 44994 19070 44996 19122
rect 44940 19068 44996 19070
rect 44716 18450 44772 18452
rect 44716 18398 44718 18450
rect 44718 18398 44770 18450
rect 44770 18398 44772 18450
rect 44716 18396 44772 18398
rect 45052 17612 45108 17668
rect 45948 20578 46004 20580
rect 45948 20526 45950 20578
rect 45950 20526 46002 20578
rect 46002 20526 46004 20578
rect 45948 20524 46004 20526
rect 47964 23212 48020 23268
rect 47516 21586 47572 21588
rect 47516 21534 47518 21586
rect 47518 21534 47570 21586
rect 47570 21534 47572 21586
rect 47516 21532 47572 21534
rect 47180 21474 47236 21476
rect 47180 21422 47182 21474
rect 47182 21422 47234 21474
rect 47234 21422 47236 21474
rect 47180 21420 47236 21422
rect 47068 19852 47124 19908
rect 46732 19404 46788 19460
rect 44828 16716 44884 16772
rect 44716 15820 44772 15876
rect 44604 13356 44660 13412
rect 44492 12236 44548 12292
rect 44604 11788 44660 11844
rect 44604 11004 44660 11060
rect 44044 8204 44100 8260
rect 43932 7756 43988 7812
rect 44604 7756 44660 7812
rect 44044 7532 44100 7588
rect 43932 6972 43988 7028
rect 43372 6860 43428 6916
rect 43932 6636 43988 6692
rect 42812 6188 42868 6244
rect 42700 5122 42756 5124
rect 42700 5070 42702 5122
rect 42702 5070 42754 5122
rect 42754 5070 42756 5122
rect 42700 5068 42756 5070
rect 43036 5906 43092 5908
rect 43036 5854 43038 5906
rect 43038 5854 43090 5906
rect 43090 5854 43092 5906
rect 43036 5852 43092 5854
rect 42924 4898 42980 4900
rect 42924 4846 42926 4898
rect 42926 4846 42978 4898
rect 42978 4846 42980 4898
rect 42924 4844 42980 4846
rect 44268 6300 44324 6356
rect 44380 4844 44436 4900
rect 42812 4284 42868 4340
rect 42476 3724 42532 3780
rect 44828 13244 44884 13300
rect 44940 13132 44996 13188
rect 44940 11394 44996 11396
rect 44940 11342 44942 11394
rect 44942 11342 44994 11394
rect 44994 11342 44996 11394
rect 44940 11340 44996 11342
rect 44828 5292 44884 5348
rect 44940 5122 44996 5124
rect 44940 5070 44942 5122
rect 44942 5070 44994 5122
rect 44994 5070 44996 5122
rect 44940 5068 44996 5070
rect 45500 17052 45556 17108
rect 46060 17164 46116 17220
rect 46396 17666 46452 17668
rect 46396 17614 46398 17666
rect 46398 17614 46450 17666
rect 46450 17614 46452 17666
rect 46396 17612 46452 17614
rect 49308 26124 49364 26180
rect 50652 31948 50708 32004
rect 51212 31948 51268 32004
rect 51772 34524 51828 34580
rect 51660 33346 51716 33348
rect 51660 33294 51662 33346
rect 51662 33294 51714 33346
rect 51714 33294 51716 33346
rect 51660 33292 51716 33294
rect 50540 31276 50596 31332
rect 50876 31500 50932 31556
rect 50988 31388 51044 31444
rect 50428 29596 50484 29652
rect 51436 31666 51492 31668
rect 51436 31614 51438 31666
rect 51438 31614 51490 31666
rect 51490 31614 51492 31666
rect 51436 31612 51492 31614
rect 51324 30994 51380 30996
rect 51324 30942 51326 30994
rect 51326 30942 51378 30994
rect 51378 30942 51380 30994
rect 51324 30940 51380 30942
rect 52220 35084 52276 35140
rect 52332 35756 52388 35812
rect 51996 33964 52052 34020
rect 51548 31388 51604 31444
rect 50316 28530 50372 28532
rect 50316 28478 50318 28530
rect 50318 28478 50370 28530
rect 50370 28478 50372 28530
rect 50316 28476 50372 28478
rect 50652 26908 50708 26964
rect 49512 25898 49568 25900
rect 49512 25846 49514 25898
rect 49514 25846 49566 25898
rect 49566 25846 49568 25898
rect 49512 25844 49568 25846
rect 49616 25898 49672 25900
rect 49616 25846 49618 25898
rect 49618 25846 49670 25898
rect 49670 25846 49672 25898
rect 49616 25844 49672 25846
rect 49720 25898 49776 25900
rect 49720 25846 49722 25898
rect 49722 25846 49774 25898
rect 49774 25846 49776 25898
rect 49720 25844 49776 25846
rect 49512 24330 49568 24332
rect 49512 24278 49514 24330
rect 49514 24278 49566 24330
rect 49566 24278 49568 24330
rect 49512 24276 49568 24278
rect 49616 24330 49672 24332
rect 49616 24278 49618 24330
rect 49618 24278 49670 24330
rect 49670 24278 49672 24330
rect 49616 24276 49672 24278
rect 49720 24330 49776 24332
rect 49720 24278 49722 24330
rect 49722 24278 49774 24330
rect 49774 24278 49776 24330
rect 49720 24276 49776 24278
rect 49420 24050 49476 24052
rect 49420 23998 49422 24050
rect 49422 23998 49474 24050
rect 49474 23998 49476 24050
rect 49420 23996 49476 23998
rect 49420 23042 49476 23044
rect 49420 22990 49422 23042
rect 49422 22990 49474 23042
rect 49474 22990 49476 23042
rect 49420 22988 49476 22990
rect 47852 20748 47908 20804
rect 47516 18956 47572 19012
rect 48188 20412 48244 20468
rect 48636 21420 48692 21476
rect 48860 21586 48916 21588
rect 48860 21534 48862 21586
rect 48862 21534 48914 21586
rect 48914 21534 48916 21586
rect 48860 21532 48916 21534
rect 48748 20802 48804 20804
rect 48748 20750 48750 20802
rect 48750 20750 48802 20802
rect 48802 20750 48804 20802
rect 48748 20748 48804 20750
rect 48636 20636 48692 20692
rect 48860 20188 48916 20244
rect 47628 18172 47684 18228
rect 47404 17724 47460 17780
rect 47068 17612 47124 17668
rect 46172 17052 46228 17108
rect 46620 17164 46676 17220
rect 45276 13356 45332 13412
rect 45276 12908 45332 12964
rect 45612 14364 45668 14420
rect 45612 14140 45668 14196
rect 46396 15874 46452 15876
rect 46396 15822 46398 15874
rect 46398 15822 46450 15874
rect 46450 15822 46452 15874
rect 46396 15820 46452 15822
rect 46060 15538 46116 15540
rect 46060 15486 46062 15538
rect 46062 15486 46114 15538
rect 46114 15486 46116 15538
rect 46060 15484 46116 15486
rect 46060 14364 46116 14420
rect 45724 13468 45780 13524
rect 45612 12684 45668 12740
rect 45500 12236 45556 12292
rect 45276 10050 45332 10052
rect 45276 9998 45278 10050
rect 45278 9998 45330 10050
rect 45330 9998 45332 10050
rect 45276 9996 45332 9998
rect 45500 11116 45556 11172
rect 45500 10444 45556 10500
rect 45276 5346 45332 5348
rect 45276 5294 45278 5346
rect 45278 5294 45330 5346
rect 45330 5294 45332 5346
rect 45276 5292 45332 5294
rect 45052 4732 45108 4788
rect 44716 3500 44772 3556
rect 39852 3162 39908 3164
rect 39852 3110 39854 3162
rect 39854 3110 39906 3162
rect 39906 3110 39908 3162
rect 39852 3108 39908 3110
rect 39956 3162 40012 3164
rect 39956 3110 39958 3162
rect 39958 3110 40010 3162
rect 40010 3110 40012 3162
rect 39956 3108 40012 3110
rect 40060 3162 40116 3164
rect 40060 3110 40062 3162
rect 40062 3110 40114 3162
rect 40114 3110 40116 3162
rect 40060 3108 40116 3110
rect 44492 3442 44548 3444
rect 44492 3390 44494 3442
rect 44494 3390 44546 3442
rect 44546 3390 44548 3442
rect 44492 3388 44548 3390
rect 45612 7084 45668 7140
rect 45724 6524 45780 6580
rect 45724 5180 45780 5236
rect 45948 13634 46004 13636
rect 45948 13582 45950 13634
rect 45950 13582 46002 13634
rect 46002 13582 46004 13634
rect 45948 13580 46004 13582
rect 46844 17052 46900 17108
rect 46956 17388 47012 17444
rect 46956 16882 47012 16884
rect 46956 16830 46958 16882
rect 46958 16830 47010 16882
rect 47010 16830 47012 16882
rect 46956 16828 47012 16830
rect 46396 13970 46452 13972
rect 46396 13918 46398 13970
rect 46398 13918 46450 13970
rect 46450 13918 46452 13970
rect 46396 13916 46452 13918
rect 46396 13132 46452 13188
rect 45948 11116 46004 11172
rect 46396 12796 46452 12852
rect 46732 13468 46788 13524
rect 47628 16828 47684 16884
rect 49512 22762 49568 22764
rect 49512 22710 49514 22762
rect 49514 22710 49566 22762
rect 49566 22710 49568 22762
rect 49512 22708 49568 22710
rect 49616 22762 49672 22764
rect 49616 22710 49618 22762
rect 49618 22710 49670 22762
rect 49670 22710 49672 22762
rect 49616 22708 49672 22710
rect 49720 22762 49776 22764
rect 49720 22710 49722 22762
rect 49722 22710 49774 22762
rect 49774 22710 49776 22762
rect 49720 22708 49776 22710
rect 49756 21756 49812 21812
rect 49868 21586 49924 21588
rect 49868 21534 49870 21586
rect 49870 21534 49922 21586
rect 49922 21534 49924 21586
rect 49868 21532 49924 21534
rect 49512 21194 49568 21196
rect 49512 21142 49514 21194
rect 49514 21142 49566 21194
rect 49566 21142 49568 21194
rect 49512 21140 49568 21142
rect 49616 21194 49672 21196
rect 49616 21142 49618 21194
rect 49618 21142 49670 21194
rect 49670 21142 49672 21194
rect 49616 21140 49672 21142
rect 49720 21194 49776 21196
rect 49720 21142 49722 21194
rect 49722 21142 49774 21194
rect 49774 21142 49776 21194
rect 49720 21140 49776 21142
rect 49084 20860 49140 20916
rect 48972 18562 49028 18564
rect 48972 18510 48974 18562
rect 48974 18510 49026 18562
rect 49026 18510 49028 18562
rect 48972 18508 49028 18510
rect 49196 18956 49252 19012
rect 48636 18284 48692 18340
rect 48748 17724 48804 17780
rect 49420 20188 49476 20244
rect 50204 26290 50260 26292
rect 50204 26238 50206 26290
rect 50206 26238 50258 26290
rect 50258 26238 50260 26290
rect 50204 26236 50260 26238
rect 50540 26796 50596 26852
rect 50876 27916 50932 27972
rect 50988 27692 51044 27748
rect 50428 26236 50484 26292
rect 50652 25788 50708 25844
rect 50316 24220 50372 24276
rect 50092 23378 50148 23380
rect 50092 23326 50094 23378
rect 50094 23326 50146 23378
rect 50146 23326 50148 23378
rect 50092 23324 50148 23326
rect 49980 20748 50036 20804
rect 50092 22316 50148 22372
rect 49868 19964 49924 20020
rect 50204 22204 50260 22260
rect 50316 21810 50372 21812
rect 50316 21758 50318 21810
rect 50318 21758 50370 21810
rect 50370 21758 50372 21810
rect 50316 21756 50372 21758
rect 50764 25394 50820 25396
rect 50764 25342 50766 25394
rect 50766 25342 50818 25394
rect 50818 25342 50820 25394
rect 50764 25340 50820 25342
rect 50764 25004 50820 25060
rect 50764 24444 50820 24500
rect 51100 26908 51156 26964
rect 51436 29148 51492 29204
rect 51436 28364 51492 28420
rect 51212 25788 51268 25844
rect 51100 24444 51156 24500
rect 50876 23996 50932 24052
rect 50652 23436 50708 23492
rect 51100 23324 51156 23380
rect 50988 22988 51044 23044
rect 50652 22316 50708 22372
rect 50876 21810 50932 21812
rect 50876 21758 50878 21810
rect 50878 21758 50930 21810
rect 50930 21758 50932 21810
rect 50876 21756 50932 21758
rect 51324 23660 51380 23716
rect 51324 23100 51380 23156
rect 51324 21980 51380 22036
rect 51436 21756 51492 21812
rect 51324 21644 51380 21700
rect 50316 20748 50372 20804
rect 50204 20690 50260 20692
rect 50204 20638 50206 20690
rect 50206 20638 50258 20690
rect 50258 20638 50260 20690
rect 50204 20636 50260 20638
rect 50988 20636 51044 20692
rect 50316 19906 50372 19908
rect 50316 19854 50318 19906
rect 50318 19854 50370 19906
rect 50370 19854 50372 19906
rect 50316 19852 50372 19854
rect 49512 19626 49568 19628
rect 49512 19574 49514 19626
rect 49514 19574 49566 19626
rect 49566 19574 49568 19626
rect 49512 19572 49568 19574
rect 49616 19626 49672 19628
rect 49616 19574 49618 19626
rect 49618 19574 49670 19626
rect 49670 19574 49672 19626
rect 49616 19572 49672 19574
rect 49720 19626 49776 19628
rect 49720 19574 49722 19626
rect 49722 19574 49774 19626
rect 49774 19574 49776 19626
rect 49720 19572 49776 19574
rect 49420 18844 49476 18900
rect 49308 18172 49364 18228
rect 49512 18058 49568 18060
rect 49512 18006 49514 18058
rect 49514 18006 49566 18058
rect 49566 18006 49568 18058
rect 49512 18004 49568 18006
rect 49616 18058 49672 18060
rect 49616 18006 49618 18058
rect 49618 18006 49670 18058
rect 49670 18006 49672 18058
rect 49616 18004 49672 18006
rect 49720 18058 49776 18060
rect 49720 18006 49722 18058
rect 49722 18006 49774 18058
rect 49774 18006 49776 18058
rect 49720 18004 49776 18006
rect 49308 17778 49364 17780
rect 49308 17726 49310 17778
rect 49310 17726 49362 17778
rect 49362 17726 49364 17778
rect 49308 17724 49364 17726
rect 48636 17052 48692 17108
rect 47404 15484 47460 15540
rect 47292 15036 47348 15092
rect 46844 13132 46900 13188
rect 46732 12684 46788 12740
rect 46620 12236 46676 12292
rect 45948 9100 46004 9156
rect 46172 9660 46228 9716
rect 45836 5740 45892 5796
rect 45948 7196 46004 7252
rect 47068 12962 47124 12964
rect 47068 12910 47070 12962
rect 47070 12910 47122 12962
rect 47122 12910 47124 12962
rect 47068 12908 47124 12910
rect 46956 12796 47012 12852
rect 47516 14418 47572 14420
rect 47516 14366 47518 14418
rect 47518 14366 47570 14418
rect 47570 14366 47572 14418
rect 47516 14364 47572 14366
rect 47292 13916 47348 13972
rect 47964 15708 48020 15764
rect 47964 14252 48020 14308
rect 47852 13804 47908 13860
rect 47292 13356 47348 13412
rect 47628 12124 47684 12180
rect 47740 13132 47796 13188
rect 47180 11676 47236 11732
rect 47068 9714 47124 9716
rect 47068 9662 47070 9714
rect 47070 9662 47122 9714
rect 47122 9662 47124 9714
rect 47068 9660 47124 9662
rect 47852 12796 47908 12852
rect 47740 9436 47796 9492
rect 48188 16604 48244 16660
rect 48412 15148 48468 15204
rect 48300 14530 48356 14532
rect 48300 14478 48302 14530
rect 48302 14478 48354 14530
rect 48354 14478 48356 14530
rect 48300 14476 48356 14478
rect 48188 14364 48244 14420
rect 48188 13692 48244 13748
rect 48300 13580 48356 13636
rect 48188 11228 48244 11284
rect 48972 16882 49028 16884
rect 48972 16830 48974 16882
rect 48974 16830 49026 16882
rect 49026 16830 49028 16882
rect 48972 16828 49028 16830
rect 48636 15708 48692 15764
rect 48636 12684 48692 12740
rect 48972 15036 49028 15092
rect 48860 14588 48916 14644
rect 48860 14140 48916 14196
rect 49512 16490 49568 16492
rect 49512 16438 49514 16490
rect 49514 16438 49566 16490
rect 49566 16438 49568 16490
rect 49512 16436 49568 16438
rect 49616 16490 49672 16492
rect 49616 16438 49618 16490
rect 49618 16438 49670 16490
rect 49670 16438 49672 16490
rect 49616 16436 49672 16438
rect 49720 16490 49776 16492
rect 49720 16438 49722 16490
rect 49722 16438 49774 16490
rect 49774 16438 49776 16490
rect 49720 16436 49776 16438
rect 49644 16156 49700 16212
rect 49512 14922 49568 14924
rect 49512 14870 49514 14922
rect 49514 14870 49566 14922
rect 49566 14870 49568 14922
rect 49512 14868 49568 14870
rect 49616 14922 49672 14924
rect 49616 14870 49618 14922
rect 49618 14870 49670 14922
rect 49670 14870 49672 14922
rect 49616 14868 49672 14870
rect 49720 14922 49776 14924
rect 49720 14870 49722 14922
rect 49722 14870 49774 14922
rect 49774 14870 49776 14922
rect 49720 14868 49776 14870
rect 49308 14476 49364 14532
rect 50428 19852 50484 19908
rect 50316 19292 50372 19348
rect 50204 18620 50260 18676
rect 49980 18284 50036 18340
rect 48860 13244 48916 13300
rect 49512 13354 49568 13356
rect 49512 13302 49514 13354
rect 49514 13302 49566 13354
rect 49566 13302 49568 13354
rect 49512 13300 49568 13302
rect 49616 13354 49672 13356
rect 49616 13302 49618 13354
rect 49618 13302 49670 13354
rect 49670 13302 49672 13354
rect 49616 13300 49672 13302
rect 49720 13354 49776 13356
rect 49720 13302 49722 13354
rect 49722 13302 49774 13354
rect 49774 13302 49776 13354
rect 49720 13300 49776 13302
rect 48972 12962 49028 12964
rect 48972 12910 48974 12962
rect 48974 12910 49026 12962
rect 49026 12910 49028 12962
rect 48972 12908 49028 12910
rect 48972 12348 49028 12404
rect 48748 11900 48804 11956
rect 49512 11786 49568 11788
rect 49512 11734 49514 11786
rect 49514 11734 49566 11786
rect 49566 11734 49568 11786
rect 49512 11732 49568 11734
rect 49616 11786 49672 11788
rect 49616 11734 49618 11786
rect 49618 11734 49670 11786
rect 49670 11734 49672 11786
rect 49616 11732 49672 11734
rect 49720 11786 49776 11788
rect 49720 11734 49722 11786
rect 49722 11734 49774 11786
rect 49774 11734 49776 11786
rect 49720 11732 49776 11734
rect 48524 11452 48580 11508
rect 50092 16882 50148 16884
rect 50092 16830 50094 16882
rect 50094 16830 50146 16882
rect 50146 16830 50148 16882
rect 50092 16828 50148 16830
rect 51100 18284 51156 18340
rect 50204 16268 50260 16324
rect 50988 16156 51044 16212
rect 50988 15538 51044 15540
rect 50988 15486 50990 15538
rect 50990 15486 51042 15538
rect 51042 15486 51044 15538
rect 50988 15484 51044 15486
rect 50764 15372 50820 15428
rect 50876 14924 50932 14980
rect 50316 14530 50372 14532
rect 50316 14478 50318 14530
rect 50318 14478 50370 14530
rect 50370 14478 50372 14530
rect 50316 14476 50372 14478
rect 50764 14140 50820 14196
rect 50428 13858 50484 13860
rect 50428 13806 50430 13858
rect 50430 13806 50482 13858
rect 50482 13806 50484 13858
rect 50428 13804 50484 13806
rect 50092 13692 50148 13748
rect 51100 14588 51156 14644
rect 51100 12908 51156 12964
rect 49980 11340 50036 11396
rect 50092 12066 50148 12068
rect 50092 12014 50094 12066
rect 50094 12014 50146 12066
rect 50146 12014 50148 12066
rect 50092 12012 50148 12014
rect 48748 11004 48804 11060
rect 48748 9772 48804 9828
rect 48076 9212 48132 9268
rect 47180 9154 47236 9156
rect 47180 9102 47182 9154
rect 47182 9102 47234 9154
rect 47234 9102 47236 9154
rect 47180 9100 47236 9102
rect 47740 9042 47796 9044
rect 47740 8990 47742 9042
rect 47742 8990 47794 9042
rect 47794 8990 47796 9042
rect 47740 8988 47796 8990
rect 48076 9042 48132 9044
rect 48076 8990 48078 9042
rect 48078 8990 48130 9042
rect 48130 8990 48132 9042
rect 48076 8988 48132 8990
rect 47292 8370 47348 8372
rect 47292 8318 47294 8370
rect 47294 8318 47346 8370
rect 47346 8318 47348 8370
rect 47292 8316 47348 8318
rect 50204 11506 50260 11508
rect 50204 11454 50206 11506
rect 50206 11454 50258 11506
rect 50258 11454 50260 11506
rect 50204 11452 50260 11454
rect 50092 10892 50148 10948
rect 50428 11228 50484 11284
rect 49512 10218 49568 10220
rect 49512 10166 49514 10218
rect 49514 10166 49566 10218
rect 49566 10166 49568 10218
rect 49512 10164 49568 10166
rect 49616 10218 49672 10220
rect 49616 10166 49618 10218
rect 49618 10166 49670 10218
rect 49670 10166 49672 10218
rect 49616 10164 49672 10166
rect 49720 10218 49776 10220
rect 49720 10166 49722 10218
rect 49722 10166 49774 10218
rect 49774 10166 49776 10218
rect 49720 10164 49776 10166
rect 48860 9100 48916 9156
rect 49308 9884 49364 9940
rect 48972 9042 49028 9044
rect 48972 8990 48974 9042
rect 48974 8990 49026 9042
rect 49026 8990 49028 9042
rect 48972 8988 49028 8990
rect 50652 10556 50708 10612
rect 49644 9266 49700 9268
rect 49644 9214 49646 9266
rect 49646 9214 49698 9266
rect 49698 9214 49700 9266
rect 49644 9212 49700 9214
rect 49308 8876 49364 8932
rect 48748 8316 48804 8372
rect 48860 8428 48916 8484
rect 46844 7532 46900 7588
rect 47404 7756 47460 7812
rect 46620 6636 46676 6692
rect 46508 5292 46564 5348
rect 46060 5010 46116 5012
rect 46060 4958 46062 5010
rect 46062 4958 46114 5010
rect 46114 4958 46116 5010
rect 46060 4956 46116 4958
rect 47068 5292 47124 5348
rect 46620 5234 46676 5236
rect 46620 5182 46622 5234
rect 46622 5182 46674 5234
rect 46674 5182 46676 5234
rect 46620 5180 46676 5182
rect 50540 8876 50596 8932
rect 49512 8650 49568 8652
rect 49512 8598 49514 8650
rect 49514 8598 49566 8650
rect 49566 8598 49568 8650
rect 49512 8596 49568 8598
rect 49616 8650 49672 8652
rect 49616 8598 49618 8650
rect 49618 8598 49670 8650
rect 49670 8598 49672 8650
rect 49616 8596 49672 8598
rect 49720 8650 49776 8652
rect 49720 8598 49722 8650
rect 49722 8598 49774 8650
rect 49774 8598 49776 8650
rect 49720 8596 49776 8598
rect 48860 7644 48916 7700
rect 48748 7196 48804 7252
rect 47852 5852 47908 5908
rect 49512 7082 49568 7084
rect 49512 7030 49514 7082
rect 49514 7030 49566 7082
rect 49566 7030 49568 7082
rect 49512 7028 49568 7030
rect 49616 7082 49672 7084
rect 49616 7030 49618 7082
rect 49618 7030 49670 7082
rect 49670 7030 49672 7082
rect 49616 7028 49672 7030
rect 49720 7082 49776 7084
rect 49720 7030 49722 7082
rect 49722 7030 49774 7082
rect 49774 7030 49776 7082
rect 49720 7028 49776 7030
rect 48972 6914 49028 6916
rect 48972 6862 48974 6914
rect 48974 6862 49026 6914
rect 49026 6862 49028 6914
rect 48972 6860 49028 6862
rect 49196 6412 49252 6468
rect 48748 6076 48804 6132
rect 48188 6018 48244 6020
rect 48188 5966 48190 6018
rect 48190 5966 48242 6018
rect 48242 5966 48244 6018
rect 48188 5964 48244 5966
rect 49532 6018 49588 6020
rect 49532 5966 49534 6018
rect 49534 5966 49586 6018
rect 49586 5966 49588 6018
rect 49532 5964 49588 5966
rect 48860 5906 48916 5908
rect 48860 5854 48862 5906
rect 48862 5854 48914 5906
rect 48914 5854 48916 5906
rect 48860 5852 48916 5854
rect 49512 5514 49568 5516
rect 49512 5462 49514 5514
rect 49514 5462 49566 5514
rect 49566 5462 49568 5514
rect 49512 5460 49568 5462
rect 49616 5514 49672 5516
rect 49616 5462 49618 5514
rect 49618 5462 49670 5514
rect 49670 5462 49672 5514
rect 49616 5460 49672 5462
rect 49720 5514 49776 5516
rect 49720 5462 49722 5514
rect 49722 5462 49774 5514
rect 49774 5462 49776 5514
rect 49720 5460 49776 5462
rect 50428 6578 50484 6580
rect 50428 6526 50430 6578
rect 50430 6526 50482 6578
rect 50482 6526 50484 6578
rect 50428 6524 50484 6526
rect 49868 4956 49924 5012
rect 49196 4844 49252 4900
rect 47964 4338 48020 4340
rect 47964 4286 47966 4338
rect 47966 4286 48018 4338
rect 48018 4286 48020 4338
rect 47964 4284 48020 4286
rect 48860 4338 48916 4340
rect 48860 4286 48862 4338
rect 48862 4286 48914 4338
rect 48914 4286 48916 4338
rect 48860 4284 48916 4286
rect 49420 4732 49476 4788
rect 49420 4450 49476 4452
rect 49420 4398 49422 4450
rect 49422 4398 49474 4450
rect 49474 4398 49476 4450
rect 49420 4396 49476 4398
rect 50988 9772 51044 9828
rect 50988 9436 51044 9492
rect 51100 8876 51156 8932
rect 50876 6412 50932 6468
rect 50652 4844 50708 4900
rect 50652 4620 50708 4676
rect 49512 3946 49568 3948
rect 49512 3894 49514 3946
rect 49514 3894 49566 3946
rect 49566 3894 49568 3946
rect 49512 3892 49568 3894
rect 49616 3946 49672 3948
rect 49616 3894 49618 3946
rect 49618 3894 49670 3946
rect 49670 3894 49672 3946
rect 49616 3892 49672 3894
rect 49720 3946 49776 3948
rect 49720 3894 49722 3946
rect 49722 3894 49774 3946
rect 49774 3894 49776 3946
rect 49720 3892 49776 3894
rect 47404 3388 47460 3444
rect 45388 2940 45444 2996
rect 45948 2716 46004 2772
rect 48524 3442 48580 3444
rect 48524 3390 48526 3442
rect 48526 3390 48578 3442
rect 48578 3390 48580 3442
rect 48524 3388 48580 3390
rect 51772 29650 51828 29652
rect 51772 29598 51774 29650
rect 51774 29598 51826 29650
rect 51826 29598 51828 29650
rect 51772 29596 51828 29598
rect 52220 29932 52276 29988
rect 51772 28924 51828 28980
rect 52108 28364 52164 28420
rect 52220 28252 52276 28308
rect 51884 27746 51940 27748
rect 51884 27694 51886 27746
rect 51886 27694 51938 27746
rect 51938 27694 51940 27746
rect 51884 27692 51940 27694
rect 51660 26796 51716 26852
rect 51772 25228 51828 25284
rect 51660 24780 51716 24836
rect 51660 23772 51716 23828
rect 51660 23378 51716 23380
rect 51660 23326 51662 23378
rect 51662 23326 51714 23378
rect 51714 23326 51716 23378
rect 51660 23324 51716 23326
rect 51660 23100 51716 23156
rect 51660 21868 51716 21924
rect 52108 26236 52164 26292
rect 51996 23772 52052 23828
rect 51996 21980 52052 22036
rect 51772 21698 51828 21700
rect 51772 21646 51774 21698
rect 51774 21646 51826 21698
rect 51826 21646 51828 21698
rect 51772 21644 51828 21646
rect 51548 21532 51604 21588
rect 51884 21532 51940 21588
rect 51772 20690 51828 20692
rect 51772 20638 51774 20690
rect 51774 20638 51826 20690
rect 51826 20638 51828 20690
rect 51772 20636 51828 20638
rect 53340 36652 53396 36708
rect 53116 35084 53172 35140
rect 53116 34860 53172 34916
rect 53564 34748 53620 34804
rect 53228 33852 53284 33908
rect 52892 29932 52948 29988
rect 52780 29820 52836 29876
rect 52556 27356 52612 27412
rect 52668 28252 52724 28308
rect 52556 26908 52612 26964
rect 53116 29596 53172 29652
rect 54908 35698 54964 35700
rect 54908 35646 54910 35698
rect 54910 35646 54962 35698
rect 54962 35646 54964 35698
rect 54908 35644 54964 35646
rect 54348 34972 54404 35028
rect 55132 34802 55188 34804
rect 55132 34750 55134 34802
rect 55134 34750 55186 34802
rect 55186 34750 55188 34802
rect 55132 34748 55188 34750
rect 53676 34412 53732 34468
rect 54460 34300 54516 34356
rect 53676 33292 53732 33348
rect 53564 30940 53620 30996
rect 54124 33964 54180 34020
rect 54348 33292 54404 33348
rect 54908 33346 54964 33348
rect 54908 33294 54910 33346
rect 54910 33294 54962 33346
rect 54962 33294 54964 33346
rect 54908 33292 54964 33294
rect 53900 31778 53956 31780
rect 53900 31726 53902 31778
rect 53902 31726 53954 31778
rect 53954 31726 53956 31778
rect 53900 31724 53956 31726
rect 53788 30434 53844 30436
rect 53788 30382 53790 30434
rect 53790 30382 53842 30434
rect 53842 30382 53844 30434
rect 53788 30380 53844 30382
rect 53452 29820 53508 29876
rect 52780 28588 52836 28644
rect 52892 28418 52948 28420
rect 52892 28366 52894 28418
rect 52894 28366 52946 28418
rect 52946 28366 52948 28418
rect 52892 28364 52948 28366
rect 53004 28252 53060 28308
rect 52892 28140 52948 28196
rect 53116 27692 53172 27748
rect 53340 28140 53396 28196
rect 53564 28364 53620 28420
rect 53788 28530 53844 28532
rect 53788 28478 53790 28530
rect 53790 28478 53842 28530
rect 53842 28478 53844 28530
rect 53788 28476 53844 28478
rect 53676 28252 53732 28308
rect 54684 29650 54740 29652
rect 54684 29598 54686 29650
rect 54686 29598 54738 29650
rect 54738 29598 54740 29650
rect 54684 29596 54740 29598
rect 54124 29148 54180 29204
rect 54460 29036 54516 29092
rect 53564 27356 53620 27412
rect 53116 26796 53172 26852
rect 53564 26796 53620 26852
rect 52668 26290 52724 26292
rect 52668 26238 52670 26290
rect 52670 26238 52722 26290
rect 52722 26238 52724 26290
rect 52668 26236 52724 26238
rect 52892 25788 52948 25844
rect 53228 25506 53284 25508
rect 53228 25454 53230 25506
rect 53230 25454 53282 25506
rect 53282 25454 53284 25506
rect 53228 25452 53284 25454
rect 53676 25506 53732 25508
rect 53676 25454 53678 25506
rect 53678 25454 53730 25506
rect 53730 25454 53732 25506
rect 53676 25452 53732 25454
rect 53788 25900 53844 25956
rect 52892 25228 52948 25284
rect 52780 24668 52836 24724
rect 54124 25228 54180 25284
rect 53788 24780 53844 24836
rect 53900 25004 53956 25060
rect 53900 24722 53956 24724
rect 53900 24670 53902 24722
rect 53902 24670 53954 24722
rect 53954 24670 53956 24722
rect 53900 24668 53956 24670
rect 53228 23938 53284 23940
rect 53228 23886 53230 23938
rect 53230 23886 53282 23938
rect 53282 23886 53284 23938
rect 53228 23884 53284 23886
rect 54796 29372 54852 29428
rect 54908 30380 54964 30436
rect 54572 28476 54628 28532
rect 54908 28530 54964 28532
rect 54908 28478 54910 28530
rect 54910 28478 54962 28530
rect 54962 28478 54964 28530
rect 54908 28476 54964 28478
rect 56028 36706 56084 36708
rect 56028 36654 56030 36706
rect 56030 36654 56082 36706
rect 56082 36654 56084 36706
rect 56028 36652 56084 36654
rect 55804 35196 55860 35252
rect 57148 35644 57204 35700
rect 58044 35420 58100 35476
rect 57148 35084 57204 35140
rect 58268 35084 58324 35140
rect 57260 34860 57316 34916
rect 55580 34354 55636 34356
rect 55580 34302 55582 34354
rect 55582 34302 55634 34354
rect 55634 34302 55636 34354
rect 55580 34300 55636 34302
rect 55356 34018 55412 34020
rect 55356 33966 55358 34018
rect 55358 33966 55410 34018
rect 55410 33966 55412 34018
rect 55356 33964 55412 33966
rect 55804 33346 55860 33348
rect 55804 33294 55806 33346
rect 55806 33294 55858 33346
rect 55858 33294 55860 33346
rect 55804 33292 55860 33294
rect 56364 33346 56420 33348
rect 56364 33294 56366 33346
rect 56366 33294 56418 33346
rect 56418 33294 56420 33346
rect 56364 33292 56420 33294
rect 56700 30828 56756 30884
rect 55468 30604 55524 30660
rect 55020 27804 55076 27860
rect 55244 27746 55300 27748
rect 55244 27694 55246 27746
rect 55246 27694 55298 27746
rect 55298 27694 55300 27746
rect 55244 27692 55300 27694
rect 54572 25506 54628 25508
rect 54572 25454 54574 25506
rect 54574 25454 54626 25506
rect 54626 25454 54628 25506
rect 54572 25452 54628 25454
rect 54796 24668 54852 24724
rect 55132 25228 55188 25284
rect 54460 24220 54516 24276
rect 53564 23100 53620 23156
rect 53900 22988 53956 23044
rect 53564 22876 53620 22932
rect 52892 21868 52948 21924
rect 52332 21810 52388 21812
rect 52332 21758 52334 21810
rect 52334 21758 52386 21810
rect 52386 21758 52388 21810
rect 52332 21756 52388 21758
rect 52108 20578 52164 20580
rect 52108 20526 52110 20578
rect 52110 20526 52162 20578
rect 52162 20526 52164 20578
rect 52108 20524 52164 20526
rect 51324 17554 51380 17556
rect 51324 17502 51326 17554
rect 51326 17502 51378 17554
rect 51378 17502 51380 17554
rect 51324 17500 51380 17502
rect 51548 16210 51604 16212
rect 51548 16158 51550 16210
rect 51550 16158 51602 16210
rect 51602 16158 51604 16210
rect 51548 16156 51604 16158
rect 51436 15932 51492 15988
rect 51436 15484 51492 15540
rect 51660 15036 51716 15092
rect 51660 13746 51716 13748
rect 51660 13694 51662 13746
rect 51662 13694 51714 13746
rect 51714 13694 51716 13746
rect 51660 13692 51716 13694
rect 51660 13020 51716 13076
rect 51772 13580 51828 13636
rect 51324 9996 51380 10052
rect 51996 18172 52052 18228
rect 52220 16492 52276 16548
rect 52220 15986 52276 15988
rect 52220 15934 52222 15986
rect 52222 15934 52274 15986
rect 52274 15934 52276 15986
rect 52220 15932 52276 15934
rect 52780 20578 52836 20580
rect 52780 20526 52782 20578
rect 52782 20526 52834 20578
rect 52834 20526 52836 20578
rect 52780 20524 52836 20526
rect 52668 20300 52724 20356
rect 52780 19852 52836 19908
rect 53228 19852 53284 19908
rect 53004 19068 53060 19124
rect 53452 18172 53508 18228
rect 52780 17554 52836 17556
rect 52780 17502 52782 17554
rect 52782 17502 52834 17554
rect 52834 17502 52836 17554
rect 52780 17500 52836 17502
rect 52892 16770 52948 16772
rect 52892 16718 52894 16770
rect 52894 16718 52946 16770
rect 52946 16718 52948 16770
rect 52892 16716 52948 16718
rect 52780 16492 52836 16548
rect 52556 16044 52612 16100
rect 51996 13468 52052 13524
rect 52108 14530 52164 14532
rect 52108 14478 52110 14530
rect 52110 14478 52162 14530
rect 52162 14478 52164 14530
rect 52108 14476 52164 14478
rect 52108 13356 52164 13412
rect 52108 11676 52164 11732
rect 51548 11340 51604 11396
rect 52108 11282 52164 11284
rect 52108 11230 52110 11282
rect 52110 11230 52162 11282
rect 52162 11230 52164 11282
rect 52108 11228 52164 11230
rect 51436 9884 51492 9940
rect 51996 9602 52052 9604
rect 51996 9550 51998 9602
rect 51998 9550 52050 9602
rect 52050 9550 52052 9602
rect 51996 9548 52052 9550
rect 51772 8316 51828 8372
rect 52780 14812 52836 14868
rect 52892 14924 52948 14980
rect 52780 14364 52836 14420
rect 53004 14140 53060 14196
rect 52556 13692 52612 13748
rect 52444 12908 52500 12964
rect 52892 12348 52948 12404
rect 52332 12178 52388 12180
rect 52332 12126 52334 12178
rect 52334 12126 52386 12178
rect 52386 12126 52388 12178
rect 52332 12124 52388 12126
rect 53340 16940 53396 16996
rect 53340 16492 53396 16548
rect 53228 14588 53284 14644
rect 52780 11282 52836 11284
rect 52780 11230 52782 11282
rect 52782 11230 52834 11282
rect 52834 11230 52836 11282
rect 52780 11228 52836 11230
rect 53116 11394 53172 11396
rect 53116 11342 53118 11394
rect 53118 11342 53170 11394
rect 53170 11342 53172 11394
rect 53116 11340 53172 11342
rect 52220 7756 52276 7812
rect 51772 6860 51828 6916
rect 52668 5852 52724 5908
rect 51212 3388 51268 3444
rect 53340 13746 53396 13748
rect 53340 13694 53342 13746
rect 53342 13694 53394 13746
rect 53394 13694 53396 13746
rect 53340 13692 53396 13694
rect 54124 24050 54180 24052
rect 54124 23998 54126 24050
rect 54126 23998 54178 24050
rect 54178 23998 54180 24050
rect 54124 23996 54180 23998
rect 54460 23938 54516 23940
rect 54460 23886 54462 23938
rect 54462 23886 54514 23938
rect 54514 23886 54516 23938
rect 54460 23884 54516 23886
rect 54236 23154 54292 23156
rect 54236 23102 54238 23154
rect 54238 23102 54290 23154
rect 54290 23102 54292 23154
rect 54236 23100 54292 23102
rect 54460 23436 54516 23492
rect 54572 22876 54628 22932
rect 54460 22428 54516 22484
rect 54684 22428 54740 22484
rect 54796 24332 54852 24388
rect 54348 20018 54404 20020
rect 54348 19966 54350 20018
rect 54350 19966 54402 20018
rect 54402 19966 54404 20018
rect 54348 19964 54404 19966
rect 54124 19068 54180 19124
rect 54236 18508 54292 18564
rect 54012 18060 54068 18116
rect 53676 17724 53732 17780
rect 53676 17276 53732 17332
rect 53900 16716 53956 16772
rect 54012 15932 54068 15988
rect 55132 25004 55188 25060
rect 54796 20188 54852 20244
rect 55020 19516 55076 19572
rect 54684 18172 54740 18228
rect 54460 17778 54516 17780
rect 54460 17726 54462 17778
rect 54462 17726 54514 17778
rect 54514 17726 54516 17778
rect 54460 17724 54516 17726
rect 54348 16882 54404 16884
rect 54348 16830 54350 16882
rect 54350 16830 54402 16882
rect 54402 16830 54404 16882
rect 54348 16828 54404 16830
rect 54348 16098 54404 16100
rect 54348 16046 54350 16098
rect 54350 16046 54402 16098
rect 54402 16046 54404 16098
rect 54348 16044 54404 16046
rect 54684 17106 54740 17108
rect 54684 17054 54686 17106
rect 54686 17054 54738 17106
rect 54738 17054 54740 17106
rect 54684 17052 54740 17054
rect 54684 16716 54740 16772
rect 54460 15932 54516 15988
rect 54908 18562 54964 18564
rect 54908 18510 54910 18562
rect 54910 18510 54962 18562
rect 54962 18510 54964 18562
rect 54908 18508 54964 18510
rect 54460 15484 54516 15540
rect 55132 18620 55188 18676
rect 55020 17836 55076 17892
rect 55020 16940 55076 16996
rect 54908 15708 54964 15764
rect 54348 14642 54404 14644
rect 54348 14590 54350 14642
rect 54350 14590 54402 14642
rect 54402 14590 54404 14642
rect 54348 14588 54404 14590
rect 53788 13804 53844 13860
rect 53564 13132 53620 13188
rect 53452 12908 53508 12964
rect 54796 15538 54852 15540
rect 54796 15486 54798 15538
rect 54798 15486 54850 15538
rect 54850 15486 54852 15538
rect 54796 15484 54852 15486
rect 56700 30268 56756 30324
rect 55580 29426 55636 29428
rect 55580 29374 55582 29426
rect 55582 29374 55634 29426
rect 55634 29374 55636 29426
rect 55580 29372 55636 29374
rect 55916 28476 55972 28532
rect 55692 27804 55748 27860
rect 56252 27804 56308 27860
rect 56700 26908 56756 26964
rect 56700 26460 56756 26516
rect 55468 26348 55524 26404
rect 55580 26236 55636 26292
rect 57932 34802 57988 34804
rect 57932 34750 57934 34802
rect 57934 34750 57986 34802
rect 57986 34750 57988 34802
rect 57932 34748 57988 34750
rect 59172 36090 59228 36092
rect 59172 36038 59174 36090
rect 59174 36038 59226 36090
rect 59226 36038 59228 36090
rect 59172 36036 59228 36038
rect 59276 36090 59332 36092
rect 59276 36038 59278 36090
rect 59278 36038 59330 36090
rect 59330 36038 59332 36090
rect 59276 36036 59332 36038
rect 59380 36090 59436 36092
rect 59380 36038 59382 36090
rect 59382 36038 59434 36090
rect 59434 36038 59436 36090
rect 59380 36036 59436 36038
rect 60620 35196 60676 35252
rect 60284 34748 60340 34804
rect 60620 34914 60676 34916
rect 60620 34862 60622 34914
rect 60622 34862 60674 34914
rect 60674 34862 60676 34914
rect 60620 34860 60676 34862
rect 58940 34524 58996 34580
rect 59172 34522 59228 34524
rect 58828 34412 58884 34468
rect 59172 34470 59174 34522
rect 59174 34470 59226 34522
rect 59226 34470 59228 34522
rect 59172 34468 59228 34470
rect 59276 34522 59332 34524
rect 59276 34470 59278 34522
rect 59278 34470 59330 34522
rect 59330 34470 59332 34522
rect 59276 34468 59332 34470
rect 59380 34522 59436 34524
rect 59380 34470 59382 34522
rect 59382 34470 59434 34522
rect 59434 34470 59436 34522
rect 59380 34468 59436 34470
rect 57596 33404 57652 33460
rect 57148 33234 57204 33236
rect 57148 33182 57150 33234
rect 57150 33182 57202 33234
rect 57202 33182 57204 33234
rect 57148 33180 57204 33182
rect 57372 32786 57428 32788
rect 57372 32734 57374 32786
rect 57374 32734 57426 32786
rect 57426 32734 57428 32786
rect 57372 32732 57428 32734
rect 57596 32396 57652 32452
rect 58044 34130 58100 34132
rect 58044 34078 58046 34130
rect 58046 34078 58098 34130
rect 58098 34078 58100 34130
rect 58044 34076 58100 34078
rect 58044 33346 58100 33348
rect 58044 33294 58046 33346
rect 58046 33294 58098 33346
rect 58098 33294 58100 33346
rect 58044 33292 58100 33294
rect 60060 34242 60116 34244
rect 60060 34190 60062 34242
rect 60062 34190 60114 34242
rect 60114 34190 60116 34242
rect 60060 34188 60116 34190
rect 62636 36482 62692 36484
rect 62636 36430 62638 36482
rect 62638 36430 62690 36482
rect 62690 36430 62692 36482
rect 62636 36428 62692 36430
rect 63196 35868 63252 35924
rect 63868 35810 63924 35812
rect 63868 35758 63870 35810
rect 63870 35758 63922 35810
rect 63922 35758 63924 35810
rect 63868 35756 63924 35758
rect 60956 34860 61012 34916
rect 61068 35420 61124 35476
rect 60732 34188 60788 34244
rect 58828 33964 58884 34020
rect 58828 33516 58884 33572
rect 59052 33346 59108 33348
rect 59052 33294 59054 33346
rect 59054 33294 59106 33346
rect 59106 33294 59108 33346
rect 59052 33292 59108 33294
rect 59276 33516 59332 33572
rect 59172 32954 59228 32956
rect 59172 32902 59174 32954
rect 59174 32902 59226 32954
rect 59226 32902 59228 32954
rect 59172 32900 59228 32902
rect 59276 32954 59332 32956
rect 59276 32902 59278 32954
rect 59278 32902 59330 32954
rect 59330 32902 59332 32954
rect 59276 32900 59332 32902
rect 59380 32954 59436 32956
rect 59380 32902 59382 32954
rect 59382 32902 59434 32954
rect 59434 32902 59436 32954
rect 59380 32900 59436 32902
rect 58156 32732 58212 32788
rect 59500 32732 59556 32788
rect 58492 32450 58548 32452
rect 58492 32398 58494 32450
rect 58494 32398 58546 32450
rect 58546 32398 58548 32450
rect 58492 32396 58548 32398
rect 57372 30156 57428 30212
rect 57148 29708 57204 29764
rect 57148 28924 57204 28980
rect 57036 27916 57092 27972
rect 57148 26908 57204 26964
rect 57148 26684 57204 26740
rect 57820 29708 57876 29764
rect 57484 29148 57540 29204
rect 57596 28364 57652 28420
rect 57484 27916 57540 27972
rect 56924 25788 56980 25844
rect 56252 24780 56308 24836
rect 57372 25228 57428 25284
rect 55356 24668 55412 24724
rect 56588 24722 56644 24724
rect 56588 24670 56590 24722
rect 56590 24670 56642 24722
rect 56642 24670 56644 24722
rect 56588 24668 56644 24670
rect 56364 24332 56420 24388
rect 56252 24050 56308 24052
rect 56252 23998 56254 24050
rect 56254 23998 56306 24050
rect 56306 23998 56308 24050
rect 56252 23996 56308 23998
rect 55468 23884 55524 23940
rect 56028 22988 56084 23044
rect 56140 22482 56196 22484
rect 56140 22430 56142 22482
rect 56142 22430 56194 22482
rect 56194 22430 56196 22482
rect 56140 22428 56196 22430
rect 57260 24668 57316 24724
rect 57036 23996 57092 24052
rect 58156 30268 58212 30324
rect 58156 29372 58212 29428
rect 59172 31386 59228 31388
rect 59172 31334 59174 31386
rect 59174 31334 59226 31386
rect 59226 31334 59228 31386
rect 59172 31332 59228 31334
rect 59276 31386 59332 31388
rect 59276 31334 59278 31386
rect 59278 31334 59330 31386
rect 59330 31334 59332 31386
rect 59276 31332 59332 31334
rect 59380 31386 59436 31388
rect 59380 31334 59382 31386
rect 59382 31334 59434 31386
rect 59434 31334 59436 31386
rect 59380 31332 59436 31334
rect 58716 30940 58772 30996
rect 58604 30604 58660 30660
rect 58716 30268 58772 30324
rect 58940 30210 58996 30212
rect 58940 30158 58942 30210
rect 58942 30158 58994 30210
rect 58994 30158 58996 30210
rect 58940 30156 58996 30158
rect 58828 30098 58884 30100
rect 58828 30046 58830 30098
rect 58830 30046 58882 30098
rect 58882 30046 58884 30098
rect 58828 30044 58884 30046
rect 59836 32786 59892 32788
rect 59836 32734 59838 32786
rect 59838 32734 59890 32786
rect 59890 32734 59892 32786
rect 59836 32732 59892 32734
rect 59612 32060 59668 32116
rect 59500 30380 59556 30436
rect 59500 30210 59556 30212
rect 59500 30158 59502 30210
rect 59502 30158 59554 30210
rect 59554 30158 59556 30210
rect 59500 30156 59556 30158
rect 57932 28642 57988 28644
rect 57932 28590 57934 28642
rect 57934 28590 57986 28642
rect 57986 28590 57988 28642
rect 57932 28588 57988 28590
rect 59172 29818 59228 29820
rect 59172 29766 59174 29818
rect 59174 29766 59226 29818
rect 59226 29766 59228 29818
rect 59172 29764 59228 29766
rect 59276 29818 59332 29820
rect 59276 29766 59278 29818
rect 59278 29766 59330 29818
rect 59330 29766 59332 29818
rect 59276 29764 59332 29766
rect 59380 29818 59436 29820
rect 59380 29766 59382 29818
rect 59382 29766 59434 29818
rect 59434 29766 59436 29818
rect 59380 29764 59436 29766
rect 59052 28812 59108 28868
rect 59276 29484 59332 29540
rect 58492 28700 58548 28756
rect 58716 28642 58772 28644
rect 58716 28590 58718 28642
rect 58718 28590 58770 28642
rect 58770 28590 58772 28642
rect 58716 28588 58772 28590
rect 58268 28476 58324 28532
rect 59276 28588 59332 28644
rect 58940 28364 58996 28420
rect 59052 28530 59108 28532
rect 59052 28478 59054 28530
rect 59054 28478 59106 28530
rect 59106 28478 59108 28530
rect 59052 28476 59108 28478
rect 59948 31724 60004 31780
rect 60060 31612 60116 31668
rect 59948 30994 60004 30996
rect 59948 30942 59950 30994
rect 59950 30942 60002 30994
rect 60002 30942 60004 30994
rect 59948 30940 60004 30942
rect 59724 30604 59780 30660
rect 59836 30380 59892 30436
rect 59724 30044 59780 30100
rect 59388 28364 59444 28420
rect 59172 28250 59228 28252
rect 59172 28198 59174 28250
rect 59174 28198 59226 28250
rect 59226 28198 59228 28250
rect 59172 28196 59228 28198
rect 59276 28250 59332 28252
rect 59276 28198 59278 28250
rect 59278 28198 59330 28250
rect 59330 28198 59332 28250
rect 59276 28196 59332 28198
rect 59380 28250 59436 28252
rect 59380 28198 59382 28250
rect 59382 28198 59434 28250
rect 59434 28198 59436 28250
rect 59380 28196 59436 28198
rect 58940 26684 58996 26740
rect 59052 27356 59108 27412
rect 58604 26514 58660 26516
rect 58604 26462 58606 26514
rect 58606 26462 58658 26514
rect 58658 26462 58660 26514
rect 58604 26460 58660 26462
rect 58940 26236 58996 26292
rect 57820 25228 57876 25284
rect 57932 24834 57988 24836
rect 57932 24782 57934 24834
rect 57934 24782 57986 24834
rect 57986 24782 57988 24834
rect 57932 24780 57988 24782
rect 57820 24556 57876 24612
rect 57820 24220 57876 24276
rect 57372 23826 57428 23828
rect 57372 23774 57374 23826
rect 57374 23774 57426 23826
rect 57426 23774 57428 23826
rect 57372 23772 57428 23774
rect 57708 23100 57764 23156
rect 58044 23996 58100 24052
rect 57036 22652 57092 22708
rect 56812 22428 56868 22484
rect 56588 21980 56644 22036
rect 56812 21532 56868 21588
rect 56812 20636 56868 20692
rect 56700 20242 56756 20244
rect 56700 20190 56702 20242
rect 56702 20190 56754 20242
rect 56754 20190 56756 20242
rect 56700 20188 56756 20190
rect 56028 19906 56084 19908
rect 56028 19854 56030 19906
rect 56030 19854 56082 19906
rect 56082 19854 56084 19906
rect 56028 19852 56084 19854
rect 55468 19516 55524 19572
rect 55468 18508 55524 18564
rect 55692 18450 55748 18452
rect 55692 18398 55694 18450
rect 55694 18398 55746 18450
rect 55746 18398 55748 18450
rect 55692 18396 55748 18398
rect 55804 18284 55860 18340
rect 55916 17836 55972 17892
rect 55468 16882 55524 16884
rect 55468 16830 55470 16882
rect 55470 16830 55522 16882
rect 55522 16830 55524 16882
rect 55468 16828 55524 16830
rect 55356 16716 55412 16772
rect 55468 16492 55524 16548
rect 55468 15426 55524 15428
rect 55468 15374 55470 15426
rect 55470 15374 55522 15426
rect 55522 15374 55524 15426
rect 55468 15372 55524 15374
rect 54684 14588 54740 14644
rect 56028 16828 56084 16884
rect 56476 18060 56532 18116
rect 57036 18620 57092 18676
rect 56700 18284 56756 18340
rect 56588 16882 56644 16884
rect 56588 16830 56590 16882
rect 56590 16830 56642 16882
rect 56642 16830 56644 16882
rect 56588 16828 56644 16830
rect 54460 13858 54516 13860
rect 54460 13806 54462 13858
rect 54462 13806 54514 13858
rect 54514 13806 54516 13858
rect 54460 13804 54516 13806
rect 54908 13746 54964 13748
rect 54908 13694 54910 13746
rect 54910 13694 54962 13746
rect 54962 13694 54964 13746
rect 54908 13692 54964 13694
rect 54348 13468 54404 13524
rect 53788 11900 53844 11956
rect 54236 11788 54292 11844
rect 53676 10444 53732 10500
rect 53452 9938 53508 9940
rect 53452 9886 53454 9938
rect 53454 9886 53506 9938
rect 53506 9886 53508 9938
rect 53452 9884 53508 9886
rect 53228 9772 53284 9828
rect 52892 9548 52948 9604
rect 53228 9042 53284 9044
rect 53228 8990 53230 9042
rect 53230 8990 53282 9042
rect 53282 8990 53284 9042
rect 53228 8988 53284 8990
rect 53900 11116 53956 11172
rect 54012 8988 54068 9044
rect 53676 8540 53732 8596
rect 55244 14140 55300 14196
rect 55468 14028 55524 14084
rect 55244 13132 55300 13188
rect 55580 13970 55636 13972
rect 55580 13918 55582 13970
rect 55582 13918 55634 13970
rect 55634 13918 55636 13970
rect 55580 13916 55636 13918
rect 55356 12962 55412 12964
rect 55356 12910 55358 12962
rect 55358 12910 55410 12962
rect 55410 12910 55412 12962
rect 55356 12908 55412 12910
rect 54572 11900 54628 11956
rect 54460 11170 54516 11172
rect 54460 11118 54462 11170
rect 54462 11118 54514 11170
rect 54514 11118 54516 11170
rect 54460 11116 54516 11118
rect 54348 10220 54404 10276
rect 54236 8316 54292 8372
rect 53676 6578 53732 6580
rect 53676 6526 53678 6578
rect 53678 6526 53730 6578
rect 53730 6526 53732 6578
rect 53676 6524 53732 6526
rect 54348 6578 54404 6580
rect 54348 6526 54350 6578
rect 54350 6526 54402 6578
rect 54402 6526 54404 6578
rect 54348 6524 54404 6526
rect 54908 11788 54964 11844
rect 55132 11788 55188 11844
rect 55132 10220 55188 10276
rect 56028 15314 56084 15316
rect 56028 15262 56030 15314
rect 56030 15262 56082 15314
rect 56082 15262 56084 15314
rect 56028 15260 56084 15262
rect 56140 14924 56196 14980
rect 56588 15708 56644 15764
rect 55916 14140 55972 14196
rect 56924 16380 56980 16436
rect 57260 18450 57316 18452
rect 57260 18398 57262 18450
rect 57262 18398 57314 18450
rect 57314 18398 57316 18450
rect 57260 18396 57316 18398
rect 57260 17948 57316 18004
rect 57260 16380 57316 16436
rect 57260 15820 57316 15876
rect 56924 15538 56980 15540
rect 56924 15486 56926 15538
rect 56926 15486 56978 15538
rect 56978 15486 56980 15538
rect 56924 15484 56980 15486
rect 56812 15260 56868 15316
rect 55916 13804 55972 13860
rect 55804 13132 55860 13188
rect 57596 21756 57652 21812
rect 57932 23714 57988 23716
rect 57932 23662 57934 23714
rect 57934 23662 57986 23714
rect 57986 23662 57988 23714
rect 57932 23660 57988 23662
rect 59612 29202 59668 29204
rect 59612 29150 59614 29202
rect 59614 29150 59666 29202
rect 59666 29150 59668 29202
rect 59612 29148 59668 29150
rect 59612 28924 59668 28980
rect 59612 28588 59668 28644
rect 60844 33516 60900 33572
rect 65436 35922 65492 35924
rect 65436 35870 65438 35922
rect 65438 35870 65490 35922
rect 65490 35870 65492 35922
rect 65436 35868 65492 35870
rect 64428 35756 64484 35812
rect 65884 36428 65940 36484
rect 66556 36482 66612 36484
rect 66556 36430 66558 36482
rect 66558 36430 66610 36482
rect 66610 36430 66612 36482
rect 66556 36428 66612 36430
rect 65884 35644 65940 35700
rect 65660 35196 65716 35252
rect 64092 35084 64148 35140
rect 63532 34300 63588 34356
rect 66444 34242 66500 34244
rect 66444 34190 66446 34242
rect 66446 34190 66498 34242
rect 66498 34190 66500 34242
rect 66444 34188 66500 34190
rect 67452 35308 67508 35364
rect 67340 34188 67396 34244
rect 64764 34076 64820 34132
rect 61292 32732 61348 32788
rect 60396 31836 60452 31892
rect 63644 34018 63700 34020
rect 63644 33966 63646 34018
rect 63646 33966 63698 34018
rect 63698 33966 63700 34018
rect 63644 33964 63700 33966
rect 61964 33570 62020 33572
rect 61964 33518 61966 33570
rect 61966 33518 62018 33570
rect 62018 33518 62020 33570
rect 61964 33516 62020 33518
rect 63644 32060 63700 32116
rect 64428 32396 64484 32452
rect 60844 31724 60900 31780
rect 60620 31666 60676 31668
rect 60620 31614 60622 31666
rect 60622 31614 60674 31666
rect 60674 31614 60676 31666
rect 60620 31612 60676 31614
rect 61516 31724 61572 31780
rect 60396 30994 60452 30996
rect 60396 30942 60398 30994
rect 60398 30942 60450 30994
rect 60450 30942 60452 30994
rect 60396 30940 60452 30942
rect 60172 30044 60228 30100
rect 59948 29426 60004 29428
rect 59948 29374 59950 29426
rect 59950 29374 60002 29426
rect 60002 29374 60004 29426
rect 59948 29372 60004 29374
rect 60284 30492 60340 30548
rect 61068 30604 61124 30660
rect 60508 30210 60564 30212
rect 60508 30158 60510 30210
rect 60510 30158 60562 30210
rect 60562 30158 60564 30210
rect 60508 30156 60564 30158
rect 60956 30210 61012 30212
rect 60956 30158 60958 30210
rect 60958 30158 61010 30210
rect 61010 30158 61012 30210
rect 60956 30156 61012 30158
rect 60396 29932 60452 29988
rect 60284 29820 60340 29876
rect 60172 28924 60228 28980
rect 59948 28866 60004 28868
rect 59948 28814 59950 28866
rect 59950 28814 60002 28866
rect 60002 28814 60004 28866
rect 59948 28812 60004 28814
rect 59172 26682 59228 26684
rect 59172 26630 59174 26682
rect 59174 26630 59226 26682
rect 59226 26630 59228 26682
rect 59172 26628 59228 26630
rect 59276 26682 59332 26684
rect 59276 26630 59278 26682
rect 59278 26630 59330 26682
rect 59330 26630 59332 26682
rect 59276 26628 59332 26630
rect 59380 26682 59436 26684
rect 59380 26630 59382 26682
rect 59382 26630 59434 26682
rect 59434 26630 59436 26682
rect 59380 26628 59436 26630
rect 60284 28364 60340 28420
rect 60172 27132 60228 27188
rect 60508 28364 60564 28420
rect 60844 29538 60900 29540
rect 60844 29486 60846 29538
rect 60846 29486 60898 29538
rect 60898 29486 60900 29538
rect 60844 29484 60900 29486
rect 60956 28812 61012 28868
rect 60284 27020 60340 27076
rect 60844 28252 60900 28308
rect 59948 26514 60004 26516
rect 59948 26462 59950 26514
rect 59950 26462 60002 26514
rect 60002 26462 60004 26514
rect 59948 26460 60004 26462
rect 59724 26290 59780 26292
rect 59724 26238 59726 26290
rect 59726 26238 59778 26290
rect 59778 26238 59780 26290
rect 59724 26236 59780 26238
rect 59388 25228 59444 25284
rect 58716 24668 58772 24724
rect 58380 23996 58436 24052
rect 58492 23714 58548 23716
rect 58492 23662 58494 23714
rect 58494 23662 58546 23714
rect 58546 23662 58548 23714
rect 58492 23660 58548 23662
rect 58828 24220 58884 24276
rect 59172 25114 59228 25116
rect 59172 25062 59174 25114
rect 59174 25062 59226 25114
rect 59226 25062 59228 25114
rect 59172 25060 59228 25062
rect 59276 25114 59332 25116
rect 59276 25062 59278 25114
rect 59278 25062 59330 25114
rect 59330 25062 59332 25114
rect 59276 25060 59332 25062
rect 59380 25114 59436 25116
rect 59380 25062 59382 25114
rect 59382 25062 59434 25114
rect 59434 25062 59436 25114
rect 59380 25060 59436 25062
rect 59612 25004 59668 25060
rect 59052 23826 59108 23828
rect 59052 23774 59054 23826
rect 59054 23774 59106 23826
rect 59106 23774 59108 23826
rect 59052 23772 59108 23774
rect 58156 22988 58212 23044
rect 58268 21980 58324 22036
rect 57484 17052 57540 17108
rect 57596 17612 57652 17668
rect 57484 16882 57540 16884
rect 57484 16830 57486 16882
rect 57486 16830 57538 16882
rect 57538 16830 57540 16882
rect 57484 16828 57540 16830
rect 57484 16156 57540 16212
rect 57372 15372 57428 15428
rect 57148 15148 57204 15204
rect 56812 15036 56868 15092
rect 56700 14530 56756 14532
rect 56700 14478 56702 14530
rect 56702 14478 56754 14530
rect 56754 14478 56756 14530
rect 56700 14476 56756 14478
rect 56364 14140 56420 14196
rect 56028 13244 56084 13300
rect 57036 14588 57092 14644
rect 56924 14418 56980 14420
rect 56924 14366 56926 14418
rect 56926 14366 56978 14418
rect 56978 14366 56980 14418
rect 56924 14364 56980 14366
rect 56812 13916 56868 13972
rect 56364 12124 56420 12180
rect 56476 13692 56532 13748
rect 56924 13580 56980 13636
rect 57036 13074 57092 13076
rect 57036 13022 57038 13074
rect 57038 13022 57090 13074
rect 57090 13022 57092 13074
rect 57036 13020 57092 13022
rect 56924 12908 56980 12964
rect 57260 14812 57316 14868
rect 57596 15148 57652 15204
rect 57372 14700 57428 14756
rect 57596 14418 57652 14420
rect 57596 14366 57598 14418
rect 57598 14366 57650 14418
rect 57650 14366 57652 14418
rect 57596 14364 57652 14366
rect 57372 13020 57428 13076
rect 57036 12850 57092 12852
rect 57036 12798 57038 12850
rect 57038 12798 57090 12850
rect 57090 12798 57092 12850
rect 57036 12796 57092 12798
rect 56700 11900 56756 11956
rect 56924 12012 56980 12068
rect 57372 12402 57428 12404
rect 57372 12350 57374 12402
rect 57374 12350 57426 12402
rect 57426 12350 57428 12402
rect 57372 12348 57428 12350
rect 57036 11788 57092 11844
rect 57260 12236 57316 12292
rect 58380 21586 58436 21588
rect 58380 21534 58382 21586
rect 58382 21534 58434 21586
rect 58434 21534 58436 21586
rect 58380 21532 58436 21534
rect 58044 19852 58100 19908
rect 57820 19234 57876 19236
rect 57820 19182 57822 19234
rect 57822 19182 57874 19234
rect 57874 19182 57876 19234
rect 57820 19180 57876 19182
rect 58268 20076 58324 20132
rect 58044 18450 58100 18452
rect 58044 18398 58046 18450
rect 58046 18398 58098 18450
rect 58098 18398 58100 18450
rect 58044 18396 58100 18398
rect 57820 18284 57876 18340
rect 58156 17836 58212 17892
rect 57820 15148 57876 15204
rect 57932 17052 57988 17108
rect 57932 16156 57988 16212
rect 58044 15708 58100 15764
rect 57820 13356 57876 13412
rect 58156 15036 58212 15092
rect 58380 17554 58436 17556
rect 58380 17502 58382 17554
rect 58382 17502 58434 17554
rect 58434 17502 58436 17554
rect 58380 17500 58436 17502
rect 58380 17276 58436 17332
rect 59612 24780 59668 24836
rect 59388 23660 59444 23716
rect 59172 23546 59228 23548
rect 59172 23494 59174 23546
rect 59174 23494 59226 23546
rect 59226 23494 59228 23546
rect 59172 23492 59228 23494
rect 59276 23546 59332 23548
rect 59276 23494 59278 23546
rect 59278 23494 59330 23546
rect 59330 23494 59332 23546
rect 59276 23492 59332 23494
rect 59380 23546 59436 23548
rect 59380 23494 59382 23546
rect 59382 23494 59434 23546
rect 59434 23494 59436 23546
rect 59380 23492 59436 23494
rect 59724 24722 59780 24724
rect 59724 24670 59726 24722
rect 59726 24670 59778 24722
rect 59778 24670 59780 24722
rect 59724 24668 59780 24670
rect 59836 24556 59892 24612
rect 59500 23154 59556 23156
rect 59500 23102 59502 23154
rect 59502 23102 59554 23154
rect 59554 23102 59556 23154
rect 59500 23100 59556 23102
rect 59948 25004 60004 25060
rect 59948 24332 60004 24388
rect 60396 24780 60452 24836
rect 59948 23884 60004 23940
rect 59500 22316 59556 22372
rect 59172 21978 59228 21980
rect 59172 21926 59174 21978
rect 59174 21926 59226 21978
rect 59226 21926 59228 21978
rect 59172 21924 59228 21926
rect 59276 21978 59332 21980
rect 59276 21926 59278 21978
rect 59278 21926 59330 21978
rect 59330 21926 59332 21978
rect 59276 21924 59332 21926
rect 59380 21978 59436 21980
rect 59380 21926 59382 21978
rect 59382 21926 59434 21978
rect 59434 21926 59436 21978
rect 59380 21924 59436 21926
rect 59052 21756 59108 21812
rect 59612 22204 59668 22260
rect 59948 22652 60004 22708
rect 60060 23548 60116 23604
rect 60396 23996 60452 24052
rect 60620 27186 60676 27188
rect 60620 27134 60622 27186
rect 60622 27134 60674 27186
rect 60674 27134 60676 27186
rect 60620 27132 60676 27134
rect 60732 26460 60788 26516
rect 60620 23714 60676 23716
rect 60620 23662 60622 23714
rect 60622 23662 60674 23714
rect 60674 23662 60676 23714
rect 60620 23660 60676 23662
rect 60620 23378 60676 23380
rect 60620 23326 60622 23378
rect 60622 23326 60674 23378
rect 60674 23326 60676 23378
rect 60620 23324 60676 23326
rect 62636 30156 62692 30212
rect 61740 30098 61796 30100
rect 61740 30046 61742 30098
rect 61742 30046 61794 30098
rect 61794 30046 61796 30098
rect 61740 30044 61796 30046
rect 61404 29932 61460 29988
rect 61180 29820 61236 29876
rect 61180 29426 61236 29428
rect 61180 29374 61182 29426
rect 61182 29374 61234 29426
rect 61234 29374 61236 29426
rect 61180 29372 61236 29374
rect 61404 28588 61460 28644
rect 61292 28476 61348 28532
rect 61628 28364 61684 28420
rect 61516 28252 61572 28308
rect 62748 29484 62804 29540
rect 62076 29372 62132 29428
rect 62076 28642 62132 28644
rect 62076 28590 62078 28642
rect 62078 28590 62130 28642
rect 62130 28590 62132 28642
rect 62076 28588 62132 28590
rect 62412 29426 62468 29428
rect 62412 29374 62414 29426
rect 62414 29374 62466 29426
rect 62466 29374 62468 29426
rect 62412 29372 62468 29374
rect 62524 28418 62580 28420
rect 62524 28366 62526 28418
rect 62526 28366 62578 28418
rect 62578 28366 62580 28418
rect 62524 28364 62580 28366
rect 62076 28252 62132 28308
rect 61180 27858 61236 27860
rect 61180 27806 61182 27858
rect 61182 27806 61234 27858
rect 61234 27806 61236 27858
rect 61180 27804 61236 27806
rect 61404 27356 61460 27412
rect 62972 28476 63028 28532
rect 62636 28252 62692 28308
rect 62300 27244 62356 27300
rect 63420 27244 63476 27300
rect 63532 27580 63588 27636
rect 61628 27074 61684 27076
rect 61628 27022 61630 27074
rect 61630 27022 61682 27074
rect 61682 27022 61684 27074
rect 61628 27020 61684 27022
rect 61292 26962 61348 26964
rect 61292 26910 61294 26962
rect 61294 26910 61346 26962
rect 61346 26910 61348 26962
rect 61292 26908 61348 26910
rect 62412 27132 62468 27188
rect 61628 26796 61684 26852
rect 61292 26460 61348 26516
rect 62188 26236 62244 26292
rect 61852 24556 61908 24612
rect 61628 24332 61684 24388
rect 61404 24162 61460 24164
rect 61404 24110 61406 24162
rect 61406 24110 61458 24162
rect 61458 24110 61460 24162
rect 61404 24108 61460 24110
rect 61292 23884 61348 23940
rect 61740 23378 61796 23380
rect 61740 23326 61742 23378
rect 61742 23326 61794 23378
rect 61794 23326 61796 23378
rect 61740 23324 61796 23326
rect 61180 23266 61236 23268
rect 61180 23214 61182 23266
rect 61182 23214 61234 23266
rect 61234 23214 61236 23266
rect 61180 23212 61236 23214
rect 60732 23154 60788 23156
rect 60732 23102 60734 23154
rect 60734 23102 60786 23154
rect 60786 23102 60788 23154
rect 60732 23100 60788 23102
rect 60172 23042 60228 23044
rect 60172 22990 60174 23042
rect 60174 22990 60226 23042
rect 60226 22990 60228 23042
rect 60172 22988 60228 22990
rect 60060 22204 60116 22260
rect 59836 21810 59892 21812
rect 59836 21758 59838 21810
rect 59838 21758 59890 21810
rect 59890 21758 59892 21810
rect 59836 21756 59892 21758
rect 59948 21420 60004 21476
rect 59724 20972 59780 21028
rect 58604 20300 58660 20356
rect 59172 20410 59228 20412
rect 59172 20358 59174 20410
rect 59174 20358 59226 20410
rect 59226 20358 59228 20410
rect 59172 20356 59228 20358
rect 59276 20410 59332 20412
rect 59276 20358 59278 20410
rect 59278 20358 59330 20410
rect 59330 20358 59332 20410
rect 59276 20356 59332 20358
rect 59380 20410 59436 20412
rect 59380 20358 59382 20410
rect 59382 20358 59434 20410
rect 59434 20358 59436 20410
rect 59380 20356 59436 20358
rect 59724 20300 59780 20356
rect 59164 20130 59220 20132
rect 59164 20078 59166 20130
rect 59166 20078 59218 20130
rect 59218 20078 59220 20130
rect 59164 20076 59220 20078
rect 59388 19964 59444 20020
rect 59276 19234 59332 19236
rect 59276 19182 59278 19234
rect 59278 19182 59330 19234
rect 59330 19182 59332 19234
rect 59276 19180 59332 19182
rect 59388 19122 59444 19124
rect 59388 19070 59390 19122
rect 59390 19070 59442 19122
rect 59442 19070 59444 19122
rect 59388 19068 59444 19070
rect 59172 18842 59228 18844
rect 59172 18790 59174 18842
rect 59174 18790 59226 18842
rect 59226 18790 59228 18842
rect 59172 18788 59228 18790
rect 59276 18842 59332 18844
rect 59276 18790 59278 18842
rect 59278 18790 59330 18842
rect 59330 18790 59332 18842
rect 59276 18788 59332 18790
rect 59380 18842 59436 18844
rect 59380 18790 59382 18842
rect 59382 18790 59434 18842
rect 59434 18790 59436 18842
rect 59380 18788 59436 18790
rect 58604 18620 58660 18676
rect 58940 18620 58996 18676
rect 58828 18396 58884 18452
rect 58716 17948 58772 18004
rect 59388 17666 59444 17668
rect 59388 17614 59390 17666
rect 59390 17614 59442 17666
rect 59442 17614 59444 17666
rect 59388 17612 59444 17614
rect 58604 17276 58660 17332
rect 58772 17276 58828 17332
rect 58492 16882 58548 16884
rect 58492 16830 58494 16882
rect 58494 16830 58546 16882
rect 58546 16830 58548 16882
rect 58492 16828 58548 16830
rect 58380 16380 58436 16436
rect 59172 17274 59228 17276
rect 59172 17222 59174 17274
rect 59174 17222 59226 17274
rect 59226 17222 59228 17274
rect 59172 17220 59228 17222
rect 59276 17274 59332 17276
rect 59276 17222 59278 17274
rect 59278 17222 59330 17274
rect 59330 17222 59332 17274
rect 59276 17220 59332 17222
rect 59380 17274 59436 17276
rect 59380 17222 59382 17274
rect 59382 17222 59434 17274
rect 59434 17222 59436 17274
rect 59380 17220 59436 17222
rect 58940 15820 58996 15876
rect 59052 16828 59108 16884
rect 59388 16210 59444 16212
rect 59388 16158 59390 16210
rect 59390 16158 59442 16210
rect 59442 16158 59444 16210
rect 59388 16156 59444 16158
rect 59172 15706 59228 15708
rect 59172 15654 59174 15706
rect 59174 15654 59226 15706
rect 59226 15654 59228 15706
rect 59172 15652 59228 15654
rect 59276 15706 59332 15708
rect 59276 15654 59278 15706
rect 59278 15654 59330 15706
rect 59330 15654 59332 15706
rect 59276 15652 59332 15654
rect 59380 15706 59436 15708
rect 59380 15654 59382 15706
rect 59382 15654 59434 15706
rect 59434 15654 59436 15706
rect 59380 15652 59436 15654
rect 58380 14252 58436 14308
rect 58492 15372 58548 15428
rect 58268 14028 58324 14084
rect 58044 13746 58100 13748
rect 58044 13694 58046 13746
rect 58046 13694 58098 13746
rect 58098 13694 58100 13746
rect 58044 13692 58100 13694
rect 57932 12850 57988 12852
rect 57932 12798 57934 12850
rect 57934 12798 57986 12850
rect 57986 12798 57988 12850
rect 57932 12796 57988 12798
rect 58380 13580 58436 13636
rect 58156 12572 58212 12628
rect 58380 13244 58436 13300
rect 58828 14700 58884 14756
rect 58604 14476 58660 14532
rect 58380 12908 58436 12964
rect 57932 12236 57988 12292
rect 58044 12178 58100 12180
rect 58044 12126 58046 12178
rect 58046 12126 58098 12178
rect 58098 12126 58100 12178
rect 58044 12124 58100 12126
rect 58268 12178 58324 12180
rect 58268 12126 58270 12178
rect 58270 12126 58322 12178
rect 58322 12126 58324 12178
rect 58268 12124 58324 12126
rect 58044 11900 58100 11956
rect 56812 11004 56868 11060
rect 55916 10722 55972 10724
rect 55916 10670 55918 10722
rect 55918 10670 55970 10722
rect 55970 10670 55972 10722
rect 55916 10668 55972 10670
rect 56812 10220 56868 10276
rect 56924 10668 56980 10724
rect 55804 9884 55860 9940
rect 55132 8092 55188 8148
rect 55244 6578 55300 6580
rect 55244 6526 55246 6578
rect 55246 6526 55298 6578
rect 55298 6526 55300 6578
rect 55244 6524 55300 6526
rect 53004 5180 53060 5236
rect 53564 5122 53620 5124
rect 53564 5070 53566 5122
rect 53566 5070 53618 5122
rect 53618 5070 53620 5122
rect 53564 5068 53620 5070
rect 54236 5122 54292 5124
rect 54236 5070 54238 5122
rect 54238 5070 54290 5122
rect 54290 5070 54292 5122
rect 54236 5068 54292 5070
rect 55804 8092 55860 8148
rect 55468 6690 55524 6692
rect 55468 6638 55470 6690
rect 55470 6638 55522 6690
rect 55522 6638 55524 6690
rect 55468 6636 55524 6638
rect 56028 7420 56084 7476
rect 56028 6690 56084 6692
rect 56028 6638 56030 6690
rect 56030 6638 56082 6690
rect 56082 6638 56084 6690
rect 56028 6636 56084 6638
rect 55580 6524 55636 6580
rect 55356 6130 55412 6132
rect 55356 6078 55358 6130
rect 55358 6078 55410 6130
rect 55410 6078 55412 6130
rect 55356 6076 55412 6078
rect 55692 6300 55748 6356
rect 55356 5292 55412 5348
rect 56028 6076 56084 6132
rect 56700 8258 56756 8260
rect 56700 8206 56702 8258
rect 56702 8206 56754 8258
rect 56754 8206 56756 8258
rect 56700 8204 56756 8206
rect 56588 6130 56644 6132
rect 56588 6078 56590 6130
rect 56590 6078 56642 6130
rect 56642 6078 56644 6130
rect 56588 6076 56644 6078
rect 55692 5068 55748 5124
rect 55356 4620 55412 4676
rect 56028 5180 56084 5236
rect 55916 5122 55972 5124
rect 55916 5070 55918 5122
rect 55918 5070 55970 5122
rect 55970 5070 55972 5122
rect 55916 5068 55972 5070
rect 56924 4396 56980 4452
rect 59500 15484 59556 15540
rect 59276 15426 59332 15428
rect 59276 15374 59278 15426
rect 59278 15374 59330 15426
rect 59330 15374 59332 15426
rect 59276 15372 59332 15374
rect 59276 14700 59332 14756
rect 61292 23154 61348 23156
rect 61292 23102 61294 23154
rect 61294 23102 61346 23154
rect 61346 23102 61348 23154
rect 61292 23100 61348 23102
rect 63308 26236 63364 26292
rect 62412 25564 62468 25620
rect 63084 25676 63140 25732
rect 62300 24556 62356 24612
rect 62748 24610 62804 24612
rect 62748 24558 62750 24610
rect 62750 24558 62802 24610
rect 62802 24558 62804 24610
rect 62748 24556 62804 24558
rect 62300 23212 62356 23268
rect 61964 23100 62020 23156
rect 63644 24722 63700 24724
rect 63644 24670 63646 24722
rect 63646 24670 63698 24722
rect 63698 24670 63700 24722
rect 63644 24668 63700 24670
rect 63196 23266 63252 23268
rect 63196 23214 63198 23266
rect 63198 23214 63250 23266
rect 63250 23214 63252 23266
rect 63196 23212 63252 23214
rect 62636 23154 62692 23156
rect 62636 23102 62638 23154
rect 62638 23102 62690 23154
rect 62690 23102 62692 23154
rect 62636 23100 62692 23102
rect 63308 23154 63364 23156
rect 63308 23102 63310 23154
rect 63310 23102 63362 23154
rect 63362 23102 63364 23154
rect 63308 23100 63364 23102
rect 60508 21756 60564 21812
rect 60620 21474 60676 21476
rect 60620 21422 60622 21474
rect 60622 21422 60674 21474
rect 60674 21422 60676 21474
rect 60620 21420 60676 21422
rect 60508 21308 60564 21364
rect 60508 20412 60564 20468
rect 62300 22092 62356 22148
rect 61068 20860 61124 20916
rect 62412 20802 62468 20804
rect 62412 20750 62414 20802
rect 62414 20750 62466 20802
rect 62466 20750 62468 20802
rect 62412 20748 62468 20750
rect 62860 20802 62916 20804
rect 62860 20750 62862 20802
rect 62862 20750 62914 20802
rect 62914 20750 62916 20802
rect 62860 20748 62916 20750
rect 60732 20636 60788 20692
rect 60956 20578 61012 20580
rect 60956 20526 60958 20578
rect 60958 20526 61010 20578
rect 61010 20526 61012 20578
rect 60956 20524 61012 20526
rect 61628 20578 61684 20580
rect 61628 20526 61630 20578
rect 61630 20526 61682 20578
rect 61682 20526 61684 20578
rect 61628 20524 61684 20526
rect 62076 20412 62132 20468
rect 60620 20188 60676 20244
rect 61628 20188 61684 20244
rect 61180 20130 61236 20132
rect 61180 20078 61182 20130
rect 61182 20078 61234 20130
rect 61234 20078 61236 20130
rect 61180 20076 61236 20078
rect 60844 20018 60900 20020
rect 60844 19966 60846 20018
rect 60846 19966 60898 20018
rect 60898 19966 60900 20018
rect 60844 19964 60900 19966
rect 61068 19740 61124 19796
rect 60172 19180 60228 19236
rect 59948 18060 60004 18116
rect 60060 18172 60116 18228
rect 60620 18060 60676 18116
rect 61404 18396 61460 18452
rect 60956 17612 61012 17668
rect 60060 17052 60116 17108
rect 59612 14530 59668 14532
rect 59612 14478 59614 14530
rect 59614 14478 59666 14530
rect 59666 14478 59668 14530
rect 59612 14476 59668 14478
rect 59276 14306 59332 14308
rect 59276 14254 59278 14306
rect 59278 14254 59330 14306
rect 59330 14254 59332 14306
rect 59276 14252 59332 14254
rect 58828 12236 58884 12292
rect 59172 14138 59228 14140
rect 59172 14086 59174 14138
rect 59174 14086 59226 14138
rect 59226 14086 59228 14138
rect 59172 14084 59228 14086
rect 59276 14138 59332 14140
rect 59276 14086 59278 14138
rect 59278 14086 59330 14138
rect 59330 14086 59332 14138
rect 59276 14084 59332 14086
rect 59380 14138 59436 14140
rect 59380 14086 59382 14138
rect 59382 14086 59434 14138
rect 59434 14086 59436 14138
rect 59380 14084 59436 14086
rect 60844 16828 60900 16884
rect 60396 15596 60452 15652
rect 59172 12570 59228 12572
rect 59172 12518 59174 12570
rect 59174 12518 59226 12570
rect 59226 12518 59228 12570
rect 59172 12516 59228 12518
rect 59276 12570 59332 12572
rect 59276 12518 59278 12570
rect 59278 12518 59330 12570
rect 59330 12518 59332 12570
rect 59276 12516 59332 12518
rect 59380 12570 59436 12572
rect 59380 12518 59382 12570
rect 59382 12518 59434 12570
rect 59434 12518 59436 12570
rect 59380 12516 59436 12518
rect 59724 13356 59780 13412
rect 59724 12796 59780 12852
rect 59052 12348 59108 12404
rect 59388 12290 59444 12292
rect 59388 12238 59390 12290
rect 59390 12238 59442 12290
rect 59442 12238 59444 12290
rect 59388 12236 59444 12238
rect 59052 11452 59108 11508
rect 58716 11004 58772 11060
rect 59500 11282 59556 11284
rect 59500 11230 59502 11282
rect 59502 11230 59554 11282
rect 59554 11230 59556 11282
rect 59500 11228 59556 11230
rect 59388 11116 59444 11172
rect 57932 9884 57988 9940
rect 57148 8146 57204 8148
rect 57148 8094 57150 8146
rect 57150 8094 57202 8146
rect 57202 8094 57204 8146
rect 57148 8092 57204 8094
rect 58380 8876 58436 8932
rect 58156 8370 58212 8372
rect 58156 8318 58158 8370
rect 58158 8318 58210 8370
rect 58210 8318 58212 8370
rect 58156 8316 58212 8318
rect 58380 8204 58436 8260
rect 57260 6690 57316 6692
rect 57260 6638 57262 6690
rect 57262 6638 57314 6690
rect 57314 6638 57316 6690
rect 57260 6636 57316 6638
rect 57372 6524 57428 6580
rect 57148 6412 57204 6468
rect 57148 5180 57204 5236
rect 58044 6578 58100 6580
rect 58044 6526 58046 6578
rect 58046 6526 58098 6578
rect 58098 6526 58100 6578
rect 58044 6524 58100 6526
rect 58268 6412 58324 6468
rect 58268 6188 58324 6244
rect 57484 5906 57540 5908
rect 57484 5854 57486 5906
rect 57486 5854 57538 5906
rect 57538 5854 57540 5906
rect 57484 5852 57540 5854
rect 57820 5122 57876 5124
rect 57820 5070 57822 5122
rect 57822 5070 57874 5122
rect 57874 5070 57876 5122
rect 57820 5068 57876 5070
rect 58156 5122 58212 5124
rect 58156 5070 58158 5122
rect 58158 5070 58210 5122
rect 58210 5070 58212 5122
rect 58156 5068 58212 5070
rect 58716 8146 58772 8148
rect 58716 8094 58718 8146
rect 58718 8094 58770 8146
rect 58770 8094 58772 8146
rect 58716 8092 58772 8094
rect 59172 11002 59228 11004
rect 59172 10950 59174 11002
rect 59174 10950 59226 11002
rect 59226 10950 59228 11002
rect 59172 10948 59228 10950
rect 59276 11002 59332 11004
rect 59276 10950 59278 11002
rect 59278 10950 59330 11002
rect 59330 10950 59332 11002
rect 59276 10948 59332 10950
rect 59380 11002 59436 11004
rect 59380 10950 59382 11002
rect 59382 10950 59434 11002
rect 59434 10950 59436 11002
rect 59380 10948 59436 10950
rect 59172 9434 59228 9436
rect 59172 9382 59174 9434
rect 59174 9382 59226 9434
rect 59226 9382 59228 9434
rect 59172 9380 59228 9382
rect 59276 9434 59332 9436
rect 59276 9382 59278 9434
rect 59278 9382 59330 9434
rect 59330 9382 59332 9434
rect 59276 9380 59332 9382
rect 59380 9434 59436 9436
rect 59380 9382 59382 9434
rect 59382 9382 59434 9434
rect 59434 9382 59436 9434
rect 59380 9380 59436 9382
rect 59836 12236 59892 12292
rect 59724 8316 59780 8372
rect 59836 8540 59892 8596
rect 59172 7866 59228 7868
rect 59172 7814 59174 7866
rect 59174 7814 59226 7866
rect 59226 7814 59228 7866
rect 59172 7812 59228 7814
rect 59276 7866 59332 7868
rect 59276 7814 59278 7866
rect 59278 7814 59330 7866
rect 59330 7814 59332 7866
rect 59276 7812 59332 7814
rect 59380 7866 59436 7868
rect 59380 7814 59382 7866
rect 59382 7814 59434 7866
rect 59434 7814 59436 7866
rect 59380 7812 59436 7814
rect 59164 6690 59220 6692
rect 59164 6638 59166 6690
rect 59166 6638 59218 6690
rect 59218 6638 59220 6690
rect 59164 6636 59220 6638
rect 59724 6466 59780 6468
rect 59724 6414 59726 6466
rect 59726 6414 59778 6466
rect 59778 6414 59780 6466
rect 59724 6412 59780 6414
rect 59172 6298 59228 6300
rect 59172 6246 59174 6298
rect 59174 6246 59226 6298
rect 59226 6246 59228 6298
rect 59172 6244 59228 6246
rect 59276 6298 59332 6300
rect 59276 6246 59278 6298
rect 59278 6246 59330 6298
rect 59330 6246 59332 6298
rect 59276 6244 59332 6246
rect 59380 6298 59436 6300
rect 59380 6246 59382 6298
rect 59382 6246 59434 6298
rect 59434 6246 59436 6298
rect 59380 6244 59436 6246
rect 60396 15260 60452 15316
rect 60732 14812 60788 14868
rect 60732 13858 60788 13860
rect 60732 13806 60734 13858
rect 60734 13806 60786 13858
rect 60786 13806 60788 13858
rect 60732 13804 60788 13806
rect 60396 12402 60452 12404
rect 60396 12350 60398 12402
rect 60398 12350 60450 12402
rect 60450 12350 60452 12402
rect 60396 12348 60452 12350
rect 61516 17500 61572 17556
rect 61852 19740 61908 19796
rect 61852 19404 61908 19460
rect 61964 18172 62020 18228
rect 60396 12178 60452 12180
rect 60396 12126 60398 12178
rect 60398 12126 60450 12178
rect 60450 12126 60452 12178
rect 60396 12124 60452 12126
rect 60732 11506 60788 11508
rect 60732 11454 60734 11506
rect 60734 11454 60786 11506
rect 60786 11454 60788 11506
rect 60732 11452 60788 11454
rect 60396 11228 60452 11284
rect 60620 8540 60676 8596
rect 59948 5964 60004 6020
rect 60508 5852 60564 5908
rect 59836 5404 59892 5460
rect 59388 5234 59444 5236
rect 59388 5182 59390 5234
rect 59390 5182 59442 5234
rect 59442 5182 59444 5234
rect 59388 5180 59444 5182
rect 58828 5122 58884 5124
rect 58828 5070 58830 5122
rect 58830 5070 58882 5122
rect 58882 5070 58884 5122
rect 58828 5068 58884 5070
rect 58716 4956 58772 5012
rect 59500 4956 59556 5012
rect 59172 4730 59228 4732
rect 59172 4678 59174 4730
rect 59174 4678 59226 4730
rect 59226 4678 59228 4730
rect 59172 4676 59228 4678
rect 59276 4730 59332 4732
rect 59276 4678 59278 4730
rect 59278 4678 59330 4730
rect 59330 4678 59332 4730
rect 59276 4676 59332 4678
rect 59380 4730 59436 4732
rect 59380 4678 59382 4730
rect 59382 4678 59434 4730
rect 59434 4678 59436 4730
rect 59380 4676 59436 4678
rect 55804 3612 55860 3668
rect 60620 5740 60676 5796
rect 60844 8930 60900 8932
rect 60844 8878 60846 8930
rect 60846 8878 60898 8930
rect 60898 8878 60900 8930
rect 60844 8876 60900 8878
rect 60844 5740 60900 5796
rect 60732 5180 60788 5236
rect 57036 3666 57092 3668
rect 57036 3614 57038 3666
rect 57038 3614 57090 3666
rect 57090 3614 57092 3666
rect 57036 3612 57092 3614
rect 59172 3162 59228 3164
rect 59172 3110 59174 3162
rect 59174 3110 59226 3162
rect 59226 3110 59228 3162
rect 59172 3108 59228 3110
rect 59276 3162 59332 3164
rect 59276 3110 59278 3162
rect 59278 3110 59330 3162
rect 59330 3110 59332 3162
rect 59276 3108 59332 3110
rect 59380 3162 59436 3164
rect 59380 3110 59382 3162
rect 59382 3110 59434 3162
rect 59434 3110 59436 3162
rect 59380 3108 59436 3110
rect 61292 14364 61348 14420
rect 61068 12402 61124 12404
rect 61068 12350 61070 12402
rect 61070 12350 61122 12402
rect 61122 12350 61124 12402
rect 61068 12348 61124 12350
rect 61740 12402 61796 12404
rect 61740 12350 61742 12402
rect 61742 12350 61794 12402
rect 61794 12350 61796 12402
rect 61740 12348 61796 12350
rect 62188 19964 62244 20020
rect 62300 19740 62356 19796
rect 62300 19516 62356 19572
rect 62188 12348 62244 12404
rect 61068 11170 61124 11172
rect 61068 11118 61070 11170
rect 61070 11118 61122 11170
rect 61122 11118 61124 11170
rect 61068 11116 61124 11118
rect 61068 9884 61124 9940
rect 61292 9266 61348 9268
rect 61292 9214 61294 9266
rect 61294 9214 61346 9266
rect 61346 9214 61348 9266
rect 61292 9212 61348 9214
rect 62412 18396 62468 18452
rect 62860 18450 62916 18452
rect 62860 18398 62862 18450
rect 62862 18398 62914 18450
rect 62914 18398 62916 18450
rect 62860 18396 62916 18398
rect 62412 17724 62468 17780
rect 62860 15820 62916 15876
rect 62412 12012 62468 12068
rect 62748 14364 62804 14420
rect 62300 9042 62356 9044
rect 62300 8990 62302 9042
rect 62302 8990 62354 9042
rect 62354 8990 62356 9042
rect 62300 8988 62356 8990
rect 61964 6860 62020 6916
rect 61740 6188 61796 6244
rect 61180 5122 61236 5124
rect 61180 5070 61182 5122
rect 61182 5070 61234 5122
rect 61234 5070 61236 5122
rect 61180 5068 61236 5070
rect 61404 5292 61460 5348
rect 61404 5068 61460 5124
rect 61628 5404 61684 5460
rect 62524 9154 62580 9156
rect 62524 9102 62526 9154
rect 62526 9102 62578 9154
rect 62578 9102 62580 9154
rect 62524 9100 62580 9102
rect 64204 23548 64260 23604
rect 63756 22988 63812 23044
rect 63084 22370 63140 22372
rect 63084 22318 63086 22370
rect 63086 22318 63138 22370
rect 63138 22318 63140 22370
rect 63084 22316 63140 22318
rect 64652 31836 64708 31892
rect 65660 34130 65716 34132
rect 65660 34078 65662 34130
rect 65662 34078 65714 34130
rect 65714 34078 65716 34130
rect 65660 34076 65716 34078
rect 65100 33516 65156 33572
rect 66444 33570 66500 33572
rect 66444 33518 66446 33570
rect 66446 33518 66498 33570
rect 66498 33518 66500 33570
rect 66444 33516 66500 33518
rect 66780 33346 66836 33348
rect 66780 33294 66782 33346
rect 66782 33294 66834 33346
rect 66834 33294 66836 33346
rect 66780 33292 66836 33294
rect 65996 33122 66052 33124
rect 65996 33070 65998 33122
rect 65998 33070 66050 33122
rect 66050 33070 66052 33122
rect 65996 33068 66052 33070
rect 66220 32450 66276 32452
rect 66220 32398 66222 32450
rect 66222 32398 66274 32450
rect 66274 32398 66276 32450
rect 66220 32396 66276 32398
rect 66668 32396 66724 32452
rect 64876 31836 64932 31892
rect 65212 31500 65268 31556
rect 64988 29596 65044 29652
rect 64540 25900 64596 25956
rect 64764 25116 64820 25172
rect 64876 24722 64932 24724
rect 64876 24670 64878 24722
rect 64878 24670 64930 24722
rect 64930 24670 64932 24722
rect 64876 24668 64932 24670
rect 64764 24050 64820 24052
rect 64764 23998 64766 24050
rect 64766 23998 64818 24050
rect 64818 23998 64820 24050
rect 64764 23996 64820 23998
rect 64876 22540 64932 22596
rect 63084 20524 63140 20580
rect 63196 19740 63252 19796
rect 63308 20300 63364 20356
rect 64316 20636 64372 20692
rect 63756 20076 63812 20132
rect 64540 20130 64596 20132
rect 64540 20078 64542 20130
rect 64542 20078 64594 20130
rect 64594 20078 64596 20130
rect 64540 20076 64596 20078
rect 63868 19628 63924 19684
rect 63868 18396 63924 18452
rect 63532 18338 63588 18340
rect 63532 18286 63534 18338
rect 63534 18286 63586 18338
rect 63586 18286 63588 18338
rect 63532 18284 63588 18286
rect 63420 17500 63476 17556
rect 63308 17388 63364 17444
rect 66332 31554 66388 31556
rect 66332 31502 66334 31554
rect 66334 31502 66386 31554
rect 66386 31502 66388 31554
rect 66332 31500 66388 31502
rect 66668 30156 66724 30212
rect 65772 29596 65828 29652
rect 65212 29148 65268 29204
rect 66556 29932 66612 29988
rect 66556 29202 66612 29204
rect 66556 29150 66558 29202
rect 66558 29150 66610 29202
rect 66610 29150 66612 29202
rect 66556 29148 66612 29150
rect 65884 28642 65940 28644
rect 65884 28590 65886 28642
rect 65886 28590 65938 28642
rect 65938 28590 65940 28642
rect 65884 28588 65940 28590
rect 65324 26908 65380 26964
rect 66220 27298 66276 27300
rect 66220 27246 66222 27298
rect 66222 27246 66274 27298
rect 66274 27246 66276 27298
rect 66220 27244 66276 27246
rect 66556 26962 66612 26964
rect 66556 26910 66558 26962
rect 66558 26910 66610 26962
rect 66610 26910 66612 26962
rect 66556 26908 66612 26910
rect 65436 26402 65492 26404
rect 65436 26350 65438 26402
rect 65438 26350 65490 26402
rect 65490 26350 65492 26402
rect 65436 26348 65492 26350
rect 65212 25452 65268 25508
rect 67676 33292 67732 33348
rect 67004 33068 67060 33124
rect 68832 36874 68888 36876
rect 68832 36822 68834 36874
rect 68834 36822 68886 36874
rect 68886 36822 68888 36874
rect 68832 36820 68888 36822
rect 68936 36874 68992 36876
rect 68936 36822 68938 36874
rect 68938 36822 68990 36874
rect 68990 36822 68992 36874
rect 68936 36820 68992 36822
rect 69040 36874 69096 36876
rect 69040 36822 69042 36874
rect 69042 36822 69094 36874
rect 69094 36822 69096 36874
rect 69040 36820 69096 36822
rect 68348 36652 68404 36708
rect 73948 38332 74004 38388
rect 73052 36652 73108 36708
rect 73724 36876 73780 36932
rect 70476 36258 70532 36260
rect 70476 36206 70478 36258
rect 70478 36206 70530 36258
rect 70530 36206 70532 36258
rect 70476 36204 70532 36206
rect 70812 36204 70868 36260
rect 72380 36316 72436 36372
rect 68124 35084 68180 35140
rect 68832 35306 68888 35308
rect 68832 35254 68834 35306
rect 68834 35254 68886 35306
rect 68886 35254 68888 35306
rect 68832 35252 68888 35254
rect 68936 35306 68992 35308
rect 68936 35254 68938 35306
rect 68938 35254 68990 35306
rect 68990 35254 68992 35306
rect 68936 35252 68992 35254
rect 69040 35306 69096 35308
rect 69040 35254 69042 35306
rect 69042 35254 69094 35306
rect 69094 35254 69096 35306
rect 69040 35252 69096 35254
rect 69356 35084 69412 35140
rect 70028 34242 70084 34244
rect 70028 34190 70030 34242
rect 70030 34190 70082 34242
rect 70082 34190 70084 34242
rect 70028 34188 70084 34190
rect 69692 34130 69748 34132
rect 69692 34078 69694 34130
rect 69694 34078 69746 34130
rect 69746 34078 69748 34130
rect 69692 34076 69748 34078
rect 69356 34018 69412 34020
rect 69356 33966 69358 34018
rect 69358 33966 69410 34018
rect 69410 33966 69412 34018
rect 69356 33964 69412 33966
rect 68832 33738 68888 33740
rect 68832 33686 68834 33738
rect 68834 33686 68886 33738
rect 68886 33686 68888 33738
rect 68832 33684 68888 33686
rect 68936 33738 68992 33740
rect 68936 33686 68938 33738
rect 68938 33686 68990 33738
rect 68990 33686 68992 33738
rect 68936 33684 68992 33686
rect 69040 33738 69096 33740
rect 69040 33686 69042 33738
rect 69042 33686 69094 33738
rect 69094 33686 69096 33738
rect 69040 33684 69096 33686
rect 70476 34130 70532 34132
rect 70476 34078 70478 34130
rect 70478 34078 70530 34130
rect 70530 34078 70532 34130
rect 70476 34076 70532 34078
rect 70924 34412 70980 34468
rect 70812 34130 70868 34132
rect 70812 34078 70814 34130
rect 70814 34078 70866 34130
rect 70866 34078 70868 34130
rect 70812 34076 70868 34078
rect 71036 33964 71092 34020
rect 69356 33068 69412 33124
rect 69692 33068 69748 33124
rect 67564 30156 67620 30212
rect 67564 29986 67620 29988
rect 67564 29934 67566 29986
rect 67566 29934 67618 29986
rect 67618 29934 67620 29986
rect 67564 29932 67620 29934
rect 67228 29820 67284 29876
rect 66892 29260 66948 29316
rect 67116 28642 67172 28644
rect 67116 28590 67118 28642
rect 67118 28590 67170 28642
rect 67170 28590 67172 28642
rect 67116 28588 67172 28590
rect 67004 27692 67060 27748
rect 66220 25452 66276 25508
rect 65996 25340 66052 25396
rect 65996 25116 66052 25172
rect 65436 23548 65492 23604
rect 65660 23378 65716 23380
rect 65660 23326 65662 23378
rect 65662 23326 65714 23378
rect 65714 23326 65716 23378
rect 65660 23324 65716 23326
rect 65548 23212 65604 23268
rect 65100 20690 65156 20692
rect 65100 20638 65102 20690
rect 65102 20638 65154 20690
rect 65154 20638 65156 20690
rect 65100 20636 65156 20638
rect 64876 20018 64932 20020
rect 64876 19966 64878 20018
rect 64878 19966 64930 20018
rect 64930 19966 64932 20018
rect 64876 19964 64932 19966
rect 64988 19628 65044 19684
rect 65660 22876 65716 22932
rect 65772 22482 65828 22484
rect 65772 22430 65774 22482
rect 65774 22430 65826 22482
rect 65826 22430 65828 22482
rect 65772 22428 65828 22430
rect 65324 21586 65380 21588
rect 65324 21534 65326 21586
rect 65326 21534 65378 21586
rect 65378 21534 65380 21586
rect 65324 21532 65380 21534
rect 65212 18956 65268 19012
rect 65436 19740 65492 19796
rect 64652 18284 64708 18340
rect 64204 17666 64260 17668
rect 64204 17614 64206 17666
rect 64206 17614 64258 17666
rect 64258 17614 64260 17666
rect 64204 17612 64260 17614
rect 63532 16604 63588 16660
rect 63644 17388 63700 17444
rect 62972 15372 63028 15428
rect 63308 15708 63364 15764
rect 63308 15148 63364 15204
rect 63532 14812 63588 14868
rect 63532 14140 63588 14196
rect 63868 16882 63924 16884
rect 63868 16830 63870 16882
rect 63870 16830 63922 16882
rect 63922 16830 63924 16882
rect 63868 16828 63924 16830
rect 65324 18172 65380 18228
rect 65660 18508 65716 18564
rect 66220 23548 66276 23604
rect 65996 22988 66052 23044
rect 65884 18284 65940 18340
rect 66220 21756 66276 21812
rect 64876 16716 64932 16772
rect 65100 17052 65156 17108
rect 64988 15874 65044 15876
rect 64988 15822 64990 15874
rect 64990 15822 65042 15874
rect 65042 15822 65044 15874
rect 64988 15820 65044 15822
rect 63868 15596 63924 15652
rect 64652 15426 64708 15428
rect 64652 15374 64654 15426
rect 64654 15374 64706 15426
rect 64706 15374 64708 15426
rect 64652 15372 64708 15374
rect 65548 16882 65604 16884
rect 65548 16830 65550 16882
rect 65550 16830 65602 16882
rect 65602 16830 65604 16882
rect 65548 16828 65604 16830
rect 64092 15036 64148 15092
rect 63644 14476 63700 14532
rect 63532 13970 63588 13972
rect 63532 13918 63534 13970
rect 63534 13918 63586 13970
rect 63586 13918 63588 13970
rect 63532 13916 63588 13918
rect 64540 14588 64596 14644
rect 63980 14364 64036 14420
rect 63868 14028 63924 14084
rect 62860 13858 62916 13860
rect 62860 13806 62862 13858
rect 62862 13806 62914 13858
rect 62914 13806 62916 13858
rect 62860 13804 62916 13806
rect 63420 13746 63476 13748
rect 63420 13694 63422 13746
rect 63422 13694 63474 13746
rect 63474 13694 63476 13746
rect 63420 13692 63476 13694
rect 65324 14700 65380 14756
rect 64876 14252 64932 14308
rect 64204 13580 64260 13636
rect 62860 13020 62916 13076
rect 63756 13074 63812 13076
rect 63756 13022 63758 13074
rect 63758 13022 63810 13074
rect 63810 13022 63812 13074
rect 63756 13020 63812 13022
rect 63980 12684 64036 12740
rect 63868 12572 63924 12628
rect 63868 12178 63924 12180
rect 63868 12126 63870 12178
rect 63870 12126 63922 12178
rect 63922 12126 63924 12178
rect 63868 12124 63924 12126
rect 63308 12012 63364 12068
rect 63868 10498 63924 10500
rect 63868 10446 63870 10498
rect 63870 10446 63922 10498
rect 63922 10446 63924 10498
rect 63868 10444 63924 10446
rect 63084 9154 63140 9156
rect 63084 9102 63086 9154
rect 63086 9102 63138 9154
rect 63138 9102 63140 9154
rect 63084 9100 63140 9102
rect 63196 8316 63252 8372
rect 62972 6636 63028 6692
rect 63084 6860 63140 6916
rect 63756 9100 63812 9156
rect 63980 8988 64036 9044
rect 64540 13356 64596 13412
rect 65996 17778 66052 17780
rect 65996 17726 65998 17778
rect 65998 17726 66050 17778
rect 66050 17726 66052 17778
rect 65996 17724 66052 17726
rect 65884 15708 65940 15764
rect 65436 14140 65492 14196
rect 65660 14588 65716 14644
rect 66780 25340 66836 25396
rect 66892 23436 66948 23492
rect 67340 25506 67396 25508
rect 67340 25454 67342 25506
rect 67342 25454 67394 25506
rect 67394 25454 67396 25506
rect 67340 25452 67396 25454
rect 69244 32450 69300 32452
rect 69244 32398 69246 32450
rect 69246 32398 69298 32450
rect 69298 32398 69300 32450
rect 69244 32396 69300 32398
rect 68832 32170 68888 32172
rect 68832 32118 68834 32170
rect 68834 32118 68886 32170
rect 68886 32118 68888 32170
rect 68832 32116 68888 32118
rect 68936 32170 68992 32172
rect 68936 32118 68938 32170
rect 68938 32118 68990 32170
rect 68990 32118 68992 32170
rect 68936 32116 68992 32118
rect 69040 32170 69096 32172
rect 69040 32118 69042 32170
rect 69042 32118 69094 32170
rect 69094 32118 69096 32170
rect 69040 32116 69096 32118
rect 69132 31500 69188 31556
rect 68832 30602 68888 30604
rect 68832 30550 68834 30602
rect 68834 30550 68886 30602
rect 68886 30550 68888 30602
rect 68832 30548 68888 30550
rect 68936 30602 68992 30604
rect 68936 30550 68938 30602
rect 68938 30550 68990 30602
rect 68990 30550 68992 30602
rect 68936 30548 68992 30550
rect 69040 30602 69096 30604
rect 69040 30550 69042 30602
rect 69042 30550 69094 30602
rect 69094 30550 69096 30602
rect 69040 30548 69096 30550
rect 69132 30380 69188 30436
rect 68572 30268 68628 30324
rect 68348 29820 68404 29876
rect 67900 29314 67956 29316
rect 67900 29262 67902 29314
rect 67902 29262 67954 29314
rect 67954 29262 67956 29314
rect 67900 29260 67956 29262
rect 68832 29034 68888 29036
rect 68832 28982 68834 29034
rect 68834 28982 68886 29034
rect 68886 28982 68888 29034
rect 68832 28980 68888 28982
rect 68936 29034 68992 29036
rect 68936 28982 68938 29034
rect 68938 28982 68990 29034
rect 68990 28982 68992 29034
rect 68936 28980 68992 28982
rect 69040 29034 69096 29036
rect 69040 28982 69042 29034
rect 69042 28982 69094 29034
rect 69094 28982 69096 29034
rect 69040 28980 69096 28982
rect 68572 27858 68628 27860
rect 68572 27806 68574 27858
rect 68574 27806 68626 27858
rect 68626 27806 68628 27858
rect 68572 27804 68628 27806
rect 68796 27746 68852 27748
rect 68796 27694 68798 27746
rect 68798 27694 68850 27746
rect 68850 27694 68852 27746
rect 68796 27692 68852 27694
rect 69020 27692 69076 27748
rect 68832 27466 68888 27468
rect 68832 27414 68834 27466
rect 68834 27414 68886 27466
rect 68886 27414 68888 27466
rect 68832 27412 68888 27414
rect 68936 27466 68992 27468
rect 68936 27414 68938 27466
rect 68938 27414 68990 27466
rect 68990 27414 68992 27466
rect 68936 27412 68992 27414
rect 69040 27466 69096 27468
rect 69040 27414 69042 27466
rect 69042 27414 69094 27466
rect 69094 27414 69096 27466
rect 69040 27412 69096 27414
rect 68684 26908 68740 26964
rect 68124 26012 68180 26068
rect 67116 23772 67172 23828
rect 67452 23212 67508 23268
rect 67340 22988 67396 23044
rect 67004 22428 67060 22484
rect 66892 21810 66948 21812
rect 66892 21758 66894 21810
rect 66894 21758 66946 21810
rect 66946 21758 66948 21810
rect 66892 21756 66948 21758
rect 66668 21420 66724 21476
rect 67116 21698 67172 21700
rect 67116 21646 67118 21698
rect 67118 21646 67170 21698
rect 67170 21646 67172 21698
rect 67116 21644 67172 21646
rect 67228 21420 67284 21476
rect 67004 20748 67060 20804
rect 67116 20076 67172 20132
rect 66444 19180 66500 19236
rect 66332 16940 66388 16996
rect 66220 16716 66276 16772
rect 67004 18844 67060 18900
rect 66780 18508 66836 18564
rect 66556 17442 66612 17444
rect 66556 17390 66558 17442
rect 66558 17390 66610 17442
rect 66610 17390 66612 17442
rect 66556 17388 66612 17390
rect 66668 17052 66724 17108
rect 66556 16828 66612 16884
rect 67228 19964 67284 20020
rect 69916 31500 69972 31556
rect 73052 34076 73108 34132
rect 72940 33458 72996 33460
rect 72940 33406 72942 33458
rect 72942 33406 72994 33458
rect 72994 33406 72996 33458
rect 72940 33404 72996 33406
rect 73164 33180 73220 33236
rect 70476 32396 70532 32452
rect 69916 31052 69972 31108
rect 69916 30380 69972 30436
rect 69692 29314 69748 29316
rect 69692 29262 69694 29314
rect 69694 29262 69746 29314
rect 69746 29262 69748 29314
rect 69692 29260 69748 29262
rect 71260 32338 71316 32340
rect 71260 32286 71262 32338
rect 71262 32286 71314 32338
rect 71314 32286 71316 32338
rect 71260 32284 71316 32286
rect 71372 30156 71428 30212
rect 71484 29932 71540 29988
rect 71036 29538 71092 29540
rect 71036 29486 71038 29538
rect 71038 29486 71090 29538
rect 71090 29486 71092 29538
rect 71036 29484 71092 29486
rect 70700 29260 70756 29316
rect 70476 29036 70532 29092
rect 69692 28588 69748 28644
rect 69356 27186 69412 27188
rect 69356 27134 69358 27186
rect 69358 27134 69410 27186
rect 69410 27134 69412 27186
rect 69356 27132 69412 27134
rect 69468 27804 69524 27860
rect 69132 26236 69188 26292
rect 68832 25898 68888 25900
rect 68832 25846 68834 25898
rect 68834 25846 68886 25898
rect 68886 25846 68888 25898
rect 68832 25844 68888 25846
rect 68936 25898 68992 25900
rect 68936 25846 68938 25898
rect 68938 25846 68990 25898
rect 68990 25846 68992 25898
rect 68936 25844 68992 25846
rect 69040 25898 69096 25900
rect 69040 25846 69042 25898
rect 69042 25846 69094 25898
rect 69094 25846 69096 25898
rect 69040 25844 69096 25846
rect 69356 26908 69412 26964
rect 70028 27634 70084 27636
rect 70028 27582 70030 27634
rect 70030 27582 70082 27634
rect 70082 27582 70084 27634
rect 70028 27580 70084 27582
rect 69468 26124 69524 26180
rect 69580 26290 69636 26292
rect 69580 26238 69582 26290
rect 69582 26238 69634 26290
rect 69634 26238 69636 26290
rect 69580 26236 69636 26238
rect 68572 25676 68628 25732
rect 68348 25506 68404 25508
rect 68348 25454 68350 25506
rect 68350 25454 68402 25506
rect 68402 25454 68404 25506
rect 68348 25452 68404 25454
rect 68236 25228 68292 25284
rect 68572 25282 68628 25284
rect 68572 25230 68574 25282
rect 68574 25230 68626 25282
rect 68626 25230 68628 25282
rect 68572 25228 68628 25230
rect 69356 25564 69412 25620
rect 69356 25394 69412 25396
rect 69356 25342 69358 25394
rect 69358 25342 69410 25394
rect 69410 25342 69412 25394
rect 69356 25340 69412 25342
rect 69020 24780 69076 24836
rect 70028 26572 70084 26628
rect 69916 26124 69972 26180
rect 69804 25788 69860 25844
rect 69580 25340 69636 25396
rect 68832 24330 68888 24332
rect 68832 24278 68834 24330
rect 68834 24278 68886 24330
rect 68886 24278 68888 24330
rect 68832 24276 68888 24278
rect 68936 24330 68992 24332
rect 68936 24278 68938 24330
rect 68938 24278 68990 24330
rect 68990 24278 68992 24330
rect 68936 24276 68992 24278
rect 69040 24330 69096 24332
rect 69040 24278 69042 24330
rect 69042 24278 69094 24330
rect 69094 24278 69096 24330
rect 69040 24276 69096 24278
rect 68908 23436 68964 23492
rect 68348 23100 68404 23156
rect 69244 23100 69300 23156
rect 68460 22876 68516 22932
rect 68832 22762 68888 22764
rect 68832 22710 68834 22762
rect 68834 22710 68886 22762
rect 68886 22710 68888 22762
rect 68832 22708 68888 22710
rect 68936 22762 68992 22764
rect 68936 22710 68938 22762
rect 68938 22710 68990 22762
rect 68990 22710 68992 22762
rect 68936 22708 68992 22710
rect 69040 22762 69096 22764
rect 69040 22710 69042 22762
rect 69042 22710 69094 22762
rect 69094 22710 69096 22762
rect 69040 22708 69096 22710
rect 71372 27970 71428 27972
rect 71372 27918 71374 27970
rect 71374 27918 71426 27970
rect 71426 27918 71428 27970
rect 71372 27916 71428 27918
rect 70364 27858 70420 27860
rect 70364 27806 70366 27858
rect 70366 27806 70418 27858
rect 70418 27806 70420 27858
rect 70364 27804 70420 27806
rect 70140 25228 70196 25284
rect 70252 27692 70308 27748
rect 70364 26572 70420 26628
rect 69468 22428 69524 22484
rect 69580 23826 69636 23828
rect 69580 23774 69582 23826
rect 69582 23774 69634 23826
rect 69634 23774 69636 23826
rect 69580 23772 69636 23774
rect 69356 22258 69412 22260
rect 69356 22206 69358 22258
rect 69358 22206 69410 22258
rect 69410 22206 69412 22258
rect 69356 22204 69412 22206
rect 68684 21756 68740 21812
rect 67564 18844 67620 18900
rect 67676 21698 67732 21700
rect 67676 21646 67678 21698
rect 67678 21646 67730 21698
rect 67730 21646 67732 21698
rect 67676 21644 67732 21646
rect 67340 16716 67396 16772
rect 66556 15820 66612 15876
rect 66108 15036 66164 15092
rect 66220 14700 66276 14756
rect 65548 13916 65604 13972
rect 65772 13916 65828 13972
rect 65436 13858 65492 13860
rect 65436 13806 65438 13858
rect 65438 13806 65490 13858
rect 65490 13806 65492 13858
rect 65436 13804 65492 13806
rect 65548 12962 65604 12964
rect 65548 12910 65550 12962
rect 65550 12910 65602 12962
rect 65602 12910 65604 12962
rect 65548 12908 65604 12910
rect 64652 12738 64708 12740
rect 64652 12686 64654 12738
rect 64654 12686 64706 12738
rect 64706 12686 64708 12738
rect 64652 12684 64708 12686
rect 65548 12684 65604 12740
rect 65100 12460 65156 12516
rect 65660 12460 65716 12516
rect 66220 13580 66276 13636
rect 66556 13692 66612 13748
rect 66444 13132 66500 13188
rect 64540 11900 64596 11956
rect 66780 13916 66836 13972
rect 66668 13356 66724 13412
rect 65212 11676 65268 11732
rect 65212 11452 65268 11508
rect 65436 11676 65492 11732
rect 64988 10722 65044 10724
rect 64988 10670 64990 10722
rect 64990 10670 65042 10722
rect 65042 10670 65044 10722
rect 64988 10668 65044 10670
rect 64988 9714 65044 9716
rect 64988 9662 64990 9714
rect 64990 9662 65042 9714
rect 65042 9662 65044 9714
rect 64988 9660 65044 9662
rect 65436 11116 65492 11172
rect 64316 8316 64372 8372
rect 63532 8092 63588 8148
rect 64092 6690 64148 6692
rect 64092 6638 64094 6690
rect 64094 6638 64146 6690
rect 64146 6638 64148 6690
rect 64092 6636 64148 6638
rect 66892 13020 66948 13076
rect 67116 13468 67172 13524
rect 66892 12178 66948 12180
rect 66892 12126 66894 12178
rect 66894 12126 66946 12178
rect 66946 12126 66948 12178
rect 66892 12124 66948 12126
rect 66780 11676 66836 11732
rect 65996 10610 66052 10612
rect 65996 10558 65998 10610
rect 65998 10558 66050 10610
rect 66050 10558 66052 10610
rect 65996 10556 66052 10558
rect 66780 10610 66836 10612
rect 66780 10558 66782 10610
rect 66782 10558 66834 10610
rect 66834 10558 66836 10610
rect 66780 10556 66836 10558
rect 65660 10498 65716 10500
rect 65660 10446 65662 10498
rect 65662 10446 65714 10498
rect 65714 10446 65716 10498
rect 65660 10444 65716 10446
rect 65884 9714 65940 9716
rect 65884 9662 65886 9714
rect 65886 9662 65938 9714
rect 65938 9662 65940 9714
rect 65884 9660 65940 9662
rect 65660 8316 65716 8372
rect 65548 8146 65604 8148
rect 65548 8094 65550 8146
rect 65550 8094 65602 8146
rect 65602 8094 65604 8146
rect 65548 8092 65604 8094
rect 63196 6018 63252 6020
rect 63196 5966 63198 6018
rect 63198 5966 63250 6018
rect 63250 5966 63252 6018
rect 63196 5964 63252 5966
rect 62972 5122 63028 5124
rect 62972 5070 62974 5122
rect 62974 5070 63026 5122
rect 63026 5070 63028 5122
rect 62972 5068 63028 5070
rect 63868 5122 63924 5124
rect 63868 5070 63870 5122
rect 63870 5070 63922 5122
rect 63922 5070 63924 5122
rect 63868 5068 63924 5070
rect 63308 5010 63364 5012
rect 63308 4958 63310 5010
rect 63310 4958 63362 5010
rect 63362 4958 63364 5010
rect 63308 4956 63364 4958
rect 65324 7532 65380 7588
rect 65660 7420 65716 7476
rect 65324 6690 65380 6692
rect 65324 6638 65326 6690
rect 65326 6638 65378 6690
rect 65378 6638 65380 6690
rect 65324 6636 65380 6638
rect 65660 6578 65716 6580
rect 65660 6526 65662 6578
rect 65662 6526 65714 6578
rect 65714 6526 65716 6578
rect 65660 6524 65716 6526
rect 65436 5906 65492 5908
rect 65436 5854 65438 5906
rect 65438 5854 65490 5906
rect 65490 5854 65492 5906
rect 65436 5852 65492 5854
rect 64988 5180 65044 5236
rect 65660 5180 65716 5236
rect 66332 8876 66388 8932
rect 66220 6690 66276 6692
rect 66220 6638 66222 6690
rect 66222 6638 66274 6690
rect 66274 6638 66276 6690
rect 66220 6636 66276 6638
rect 67228 13132 67284 13188
rect 68832 21194 68888 21196
rect 68832 21142 68834 21194
rect 68834 21142 68886 21194
rect 68886 21142 68888 21194
rect 68832 21140 68888 21142
rect 68936 21194 68992 21196
rect 68936 21142 68938 21194
rect 68938 21142 68990 21194
rect 68990 21142 68992 21194
rect 68936 21140 68992 21142
rect 69040 21194 69096 21196
rect 69040 21142 69042 21194
rect 69042 21142 69094 21194
rect 69094 21142 69096 21194
rect 69040 21140 69096 21142
rect 68460 20300 68516 20356
rect 67676 17612 67732 17668
rect 67564 17500 67620 17556
rect 67676 17388 67732 17444
rect 67564 15596 67620 15652
rect 68124 18450 68180 18452
rect 68124 18398 68126 18450
rect 68126 18398 68178 18450
rect 68178 18398 68180 18450
rect 68124 18396 68180 18398
rect 69020 20300 69076 20356
rect 68684 19852 68740 19908
rect 68460 17164 68516 17220
rect 67900 16940 67956 16996
rect 67900 15820 67956 15876
rect 69020 19740 69076 19796
rect 68832 19626 68888 19628
rect 68832 19574 68834 19626
rect 68834 19574 68886 19626
rect 68886 19574 68888 19626
rect 68832 19572 68888 19574
rect 68936 19626 68992 19628
rect 68936 19574 68938 19626
rect 68938 19574 68990 19626
rect 68990 19574 68992 19626
rect 68936 19572 68992 19574
rect 69040 19626 69096 19628
rect 69040 19574 69042 19626
rect 69042 19574 69094 19626
rect 69094 19574 69096 19626
rect 69040 19572 69096 19574
rect 69468 22146 69524 22148
rect 69468 22094 69470 22146
rect 69470 22094 69522 22146
rect 69522 22094 69524 22146
rect 69468 22092 69524 22094
rect 69692 23324 69748 23380
rect 69580 21420 69636 21476
rect 69692 21532 69748 21588
rect 69356 20076 69412 20132
rect 69580 20018 69636 20020
rect 69580 19966 69582 20018
rect 69582 19966 69634 20018
rect 69634 19966 69636 20018
rect 69580 19964 69636 19966
rect 70252 23884 70308 23940
rect 69916 22876 69972 22932
rect 69916 22092 69972 22148
rect 70028 20914 70084 20916
rect 70028 20862 70030 20914
rect 70030 20862 70082 20914
rect 70082 20862 70084 20914
rect 70028 20860 70084 20862
rect 70476 26124 70532 26180
rect 70700 25452 70756 25508
rect 71260 27858 71316 27860
rect 71260 27806 71262 27858
rect 71262 27806 71314 27858
rect 71314 27806 71316 27858
rect 71260 27804 71316 27806
rect 71148 27692 71204 27748
rect 70812 26348 70868 26404
rect 70476 25116 70532 25172
rect 71036 26402 71092 26404
rect 71036 26350 71038 26402
rect 71038 26350 71090 26402
rect 71090 26350 71092 26402
rect 71036 26348 71092 26350
rect 72268 29538 72324 29540
rect 72268 29486 72270 29538
rect 72270 29486 72322 29538
rect 72322 29486 72324 29538
rect 72268 29484 72324 29486
rect 72716 29484 72772 29540
rect 72044 29036 72100 29092
rect 71932 28642 71988 28644
rect 71932 28590 71934 28642
rect 71934 28590 71986 28642
rect 71986 28590 71988 28642
rect 71932 28588 71988 28590
rect 71596 27858 71652 27860
rect 71596 27806 71598 27858
rect 71598 27806 71650 27858
rect 71650 27806 71652 27858
rect 71596 27804 71652 27806
rect 72492 28588 72548 28644
rect 72716 29260 72772 29316
rect 72828 29148 72884 29204
rect 71148 25564 71204 25620
rect 70364 22988 70420 23044
rect 70588 23154 70644 23156
rect 70588 23102 70590 23154
rect 70590 23102 70642 23154
rect 70642 23102 70644 23154
rect 70588 23100 70644 23102
rect 70476 22428 70532 22484
rect 70364 22092 70420 22148
rect 69692 19292 69748 19348
rect 68908 19068 68964 19124
rect 69244 18396 69300 18452
rect 69804 19068 69860 19124
rect 69916 19010 69972 19012
rect 69916 18958 69918 19010
rect 69918 18958 69970 19010
rect 69970 18958 69972 19010
rect 69916 18956 69972 18958
rect 68832 18058 68888 18060
rect 68832 18006 68834 18058
rect 68834 18006 68886 18058
rect 68886 18006 68888 18058
rect 68832 18004 68888 18006
rect 68936 18058 68992 18060
rect 68936 18006 68938 18058
rect 68938 18006 68990 18058
rect 68990 18006 68992 18058
rect 68936 18004 68992 18006
rect 69040 18058 69096 18060
rect 69040 18006 69042 18058
rect 69042 18006 69094 18058
rect 69094 18006 69096 18058
rect 69040 18004 69096 18006
rect 68796 17836 68852 17892
rect 69356 17724 69412 17780
rect 69916 18450 69972 18452
rect 69916 18398 69918 18450
rect 69918 18398 69970 18450
rect 69970 18398 69972 18450
rect 69916 18396 69972 18398
rect 70028 18284 70084 18340
rect 70700 22204 70756 22260
rect 71036 23938 71092 23940
rect 71036 23886 71038 23938
rect 71038 23886 71090 23938
rect 71090 23886 71092 23938
rect 71036 23884 71092 23886
rect 70812 22988 70868 23044
rect 70588 21308 70644 21364
rect 70700 21868 70756 21924
rect 70700 21084 70756 21140
rect 70588 20860 70644 20916
rect 70812 20860 70868 20916
rect 70476 19852 70532 19908
rect 68908 17276 68964 17332
rect 69468 17164 69524 17220
rect 68832 16490 68888 16492
rect 68832 16438 68834 16490
rect 68834 16438 68886 16490
rect 68886 16438 68888 16490
rect 68832 16436 68888 16438
rect 68936 16490 68992 16492
rect 68936 16438 68938 16490
rect 68938 16438 68990 16490
rect 68990 16438 68992 16490
rect 68936 16436 68992 16438
rect 69040 16490 69096 16492
rect 69040 16438 69042 16490
rect 69042 16438 69094 16490
rect 69094 16438 69096 16490
rect 69040 16436 69096 16438
rect 69132 16322 69188 16324
rect 69132 16270 69134 16322
rect 69134 16270 69186 16322
rect 69186 16270 69188 16322
rect 69132 16268 69188 16270
rect 68348 15596 68404 15652
rect 68236 14364 68292 14420
rect 68832 14922 68888 14924
rect 68832 14870 68834 14922
rect 68834 14870 68886 14922
rect 68886 14870 68888 14922
rect 68832 14868 68888 14870
rect 68936 14922 68992 14924
rect 68936 14870 68938 14922
rect 68938 14870 68990 14922
rect 68990 14870 68992 14922
rect 68936 14868 68992 14870
rect 69040 14922 69096 14924
rect 69040 14870 69042 14922
rect 69042 14870 69094 14922
rect 69094 14870 69096 14922
rect 69040 14868 69096 14870
rect 68908 14364 68964 14420
rect 68684 13804 68740 13860
rect 68460 13692 68516 13748
rect 67900 13356 67956 13412
rect 67452 12908 67508 12964
rect 67228 11676 67284 11732
rect 67788 10668 67844 10724
rect 68124 11452 68180 11508
rect 68124 10668 68180 10724
rect 67900 8930 67956 8932
rect 67900 8878 67902 8930
rect 67902 8878 67954 8930
rect 67954 8878 67956 8930
rect 67900 8876 67956 8878
rect 68832 13354 68888 13356
rect 68832 13302 68834 13354
rect 68834 13302 68886 13354
rect 68886 13302 68888 13354
rect 68832 13300 68888 13302
rect 68936 13354 68992 13356
rect 68936 13302 68938 13354
rect 68938 13302 68990 13354
rect 68990 13302 68992 13354
rect 68936 13300 68992 13302
rect 69040 13354 69096 13356
rect 69040 13302 69042 13354
rect 69042 13302 69094 13354
rect 69094 13302 69096 13354
rect 69040 13300 69096 13302
rect 69244 12124 69300 12180
rect 68832 11786 68888 11788
rect 68832 11734 68834 11786
rect 68834 11734 68886 11786
rect 68886 11734 68888 11786
rect 68832 11732 68888 11734
rect 68936 11786 68992 11788
rect 68936 11734 68938 11786
rect 68938 11734 68990 11786
rect 68990 11734 68992 11786
rect 68936 11732 68992 11734
rect 69040 11786 69096 11788
rect 69040 11734 69042 11786
rect 69042 11734 69094 11786
rect 69094 11734 69096 11786
rect 69040 11732 69096 11734
rect 69356 10722 69412 10724
rect 69356 10670 69358 10722
rect 69358 10670 69410 10722
rect 69410 10670 69412 10722
rect 69356 10668 69412 10670
rect 68572 10498 68628 10500
rect 68572 10446 68574 10498
rect 68574 10446 68626 10498
rect 68626 10446 68628 10498
rect 68572 10444 68628 10446
rect 69132 10444 69188 10500
rect 68832 10218 68888 10220
rect 68832 10166 68834 10218
rect 68834 10166 68886 10218
rect 68886 10166 68888 10218
rect 68832 10164 68888 10166
rect 68936 10218 68992 10220
rect 68936 10166 68938 10218
rect 68938 10166 68990 10218
rect 68990 10166 68992 10218
rect 68936 10164 68992 10166
rect 69040 10218 69096 10220
rect 69040 10166 69042 10218
rect 69042 10166 69094 10218
rect 69094 10166 69096 10218
rect 69040 10164 69096 10166
rect 68908 9996 68964 10052
rect 68572 9826 68628 9828
rect 68572 9774 68574 9826
rect 68574 9774 68626 9826
rect 68626 9774 68628 9826
rect 68572 9772 68628 9774
rect 69580 16828 69636 16884
rect 69804 17666 69860 17668
rect 69804 17614 69806 17666
rect 69806 17614 69858 17666
rect 69858 17614 69860 17666
rect 69804 17612 69860 17614
rect 69804 16994 69860 16996
rect 69804 16942 69806 16994
rect 69806 16942 69858 16994
rect 69858 16942 69860 16994
rect 69804 16940 69860 16942
rect 69580 13468 69636 13524
rect 69692 14476 69748 14532
rect 70028 14588 70084 14644
rect 70252 19346 70308 19348
rect 70252 19294 70254 19346
rect 70254 19294 70306 19346
rect 70306 19294 70308 19346
rect 70252 19292 70308 19294
rect 70252 19010 70308 19012
rect 70252 18958 70254 19010
rect 70254 18958 70306 19010
rect 70306 18958 70308 19010
rect 70252 18956 70308 18958
rect 70812 19740 70868 19796
rect 71260 24780 71316 24836
rect 71036 22764 71092 22820
rect 71036 21868 71092 21924
rect 72156 27074 72212 27076
rect 72156 27022 72158 27074
rect 72158 27022 72210 27074
rect 72210 27022 72212 27074
rect 72156 27020 72212 27022
rect 71932 26012 71988 26068
rect 73276 33404 73332 33460
rect 73276 32284 73332 32340
rect 72828 27858 72884 27860
rect 72828 27806 72830 27858
rect 72830 27806 72882 27858
rect 72882 27806 72884 27858
rect 72828 27804 72884 27806
rect 72604 27020 72660 27076
rect 72492 26124 72548 26180
rect 72380 25900 72436 25956
rect 72156 25676 72212 25732
rect 71596 24668 71652 24724
rect 71708 24108 71764 24164
rect 71820 24220 71876 24276
rect 71484 23212 71540 23268
rect 71372 21644 71428 21700
rect 70588 18844 70644 18900
rect 70588 18508 70644 18564
rect 70476 17276 70532 17332
rect 70364 14364 70420 14420
rect 70812 18620 70868 18676
rect 70812 18284 70868 18340
rect 71148 21308 71204 21364
rect 71820 23548 71876 23604
rect 71596 22876 71652 22932
rect 71484 20636 71540 20692
rect 71596 22204 71652 22260
rect 72156 25228 72212 25284
rect 72268 25116 72324 25172
rect 72380 25452 72436 25508
rect 72268 24220 72324 24276
rect 72716 25452 72772 25508
rect 72604 24722 72660 24724
rect 72604 24670 72606 24722
rect 72606 24670 72658 24722
rect 72658 24670 72660 24722
rect 72604 24668 72660 24670
rect 72604 23884 72660 23940
rect 72044 23772 72100 23828
rect 72268 23826 72324 23828
rect 72268 23774 72270 23826
rect 72270 23774 72322 23826
rect 72322 23774 72324 23826
rect 72268 23772 72324 23774
rect 72156 23548 72212 23604
rect 72828 23772 72884 23828
rect 72268 23436 72324 23492
rect 72380 23548 72436 23604
rect 72156 23324 72212 23380
rect 72268 22876 72324 22932
rect 72268 22652 72324 22708
rect 71932 22204 71988 22260
rect 73164 25564 73220 25620
rect 73052 24780 73108 24836
rect 73276 25228 73332 25284
rect 73052 24108 73108 24164
rect 72716 23212 72772 23268
rect 72492 23100 72548 23156
rect 71708 21532 71764 21588
rect 72604 21810 72660 21812
rect 72604 21758 72606 21810
rect 72606 21758 72658 21810
rect 72658 21758 72660 21810
rect 72604 21756 72660 21758
rect 72828 23154 72884 23156
rect 72828 23102 72830 23154
rect 72830 23102 72882 23154
rect 72882 23102 72884 23154
rect 72828 23100 72884 23102
rect 73500 27692 73556 27748
rect 73724 30210 73780 30212
rect 73724 30158 73726 30210
rect 73726 30158 73778 30210
rect 73778 30158 73780 30210
rect 73724 30156 73780 30158
rect 74060 36876 74116 36932
rect 75068 36706 75124 36708
rect 75068 36654 75070 36706
rect 75070 36654 75122 36706
rect 75122 36654 75124 36706
rect 75068 36652 75124 36654
rect 75516 35868 75572 35924
rect 76636 35922 76692 35924
rect 76636 35870 76638 35922
rect 76638 35870 76690 35922
rect 76690 35870 76692 35922
rect 76636 35868 76692 35870
rect 75068 35756 75124 35812
rect 76300 34524 76356 34580
rect 75068 34076 75124 34132
rect 73948 31164 74004 31220
rect 73836 29314 73892 29316
rect 73836 29262 73838 29314
rect 73838 29262 73890 29314
rect 73890 29262 73892 29314
rect 73836 29260 73892 29262
rect 74172 31106 74228 31108
rect 74172 31054 74174 31106
rect 74174 31054 74226 31106
rect 74226 31054 74228 31106
rect 74172 31052 74228 31054
rect 74508 30156 74564 30212
rect 74732 29260 74788 29316
rect 73948 29036 74004 29092
rect 73836 28588 73892 28644
rect 73724 28140 73780 28196
rect 73500 25506 73556 25508
rect 73500 25454 73502 25506
rect 73502 25454 73554 25506
rect 73554 25454 73556 25506
rect 73500 25452 73556 25454
rect 73724 24892 73780 24948
rect 78492 36090 78548 36092
rect 78492 36038 78494 36090
rect 78494 36038 78546 36090
rect 78546 36038 78548 36090
rect 78492 36036 78548 36038
rect 78596 36090 78652 36092
rect 78596 36038 78598 36090
rect 78598 36038 78650 36090
rect 78650 36038 78652 36090
rect 78596 36036 78652 36038
rect 78700 36090 78756 36092
rect 78700 36038 78702 36090
rect 78702 36038 78754 36090
rect 78754 36038 78756 36090
rect 78700 36036 78756 36038
rect 78492 34522 78548 34524
rect 78492 34470 78494 34522
rect 78494 34470 78546 34522
rect 78546 34470 78548 34522
rect 78492 34468 78548 34470
rect 78596 34522 78652 34524
rect 78596 34470 78598 34522
rect 78598 34470 78650 34522
rect 78650 34470 78652 34522
rect 78596 34468 78652 34470
rect 78700 34522 78756 34524
rect 78700 34470 78702 34522
rect 78702 34470 78754 34522
rect 78754 34470 78756 34522
rect 78700 34468 78756 34470
rect 77980 34076 78036 34132
rect 77980 33404 78036 33460
rect 76300 33234 76356 33236
rect 76300 33182 76302 33234
rect 76302 33182 76354 33234
rect 76354 33182 76356 33234
rect 76300 33180 76356 33182
rect 75404 33122 75460 33124
rect 75404 33070 75406 33122
rect 75406 33070 75458 33122
rect 75458 33070 75460 33122
rect 75404 33068 75460 33070
rect 78492 32954 78548 32956
rect 78492 32902 78494 32954
rect 78494 32902 78546 32954
rect 78546 32902 78548 32954
rect 78492 32900 78548 32902
rect 78596 32954 78652 32956
rect 78596 32902 78598 32954
rect 78598 32902 78650 32954
rect 78650 32902 78652 32954
rect 78596 32900 78652 32902
rect 78700 32954 78756 32956
rect 78700 32902 78702 32954
rect 78702 32902 78754 32954
rect 78754 32902 78756 32954
rect 78700 32900 78756 32902
rect 75180 28140 75236 28196
rect 75292 30828 75348 30884
rect 73948 26348 74004 26404
rect 75404 30044 75460 30100
rect 75628 30156 75684 30212
rect 75516 29932 75572 29988
rect 78492 31386 78548 31388
rect 78492 31334 78494 31386
rect 78494 31334 78546 31386
rect 78546 31334 78548 31386
rect 78492 31332 78548 31334
rect 78596 31386 78652 31388
rect 78596 31334 78598 31386
rect 78598 31334 78650 31386
rect 78650 31334 78652 31386
rect 78596 31332 78652 31334
rect 78700 31386 78756 31388
rect 78700 31334 78702 31386
rect 78702 31334 78754 31386
rect 78754 31334 78756 31386
rect 78700 31332 78756 31334
rect 77980 30940 78036 30996
rect 77756 30882 77812 30884
rect 77756 30830 77758 30882
rect 77758 30830 77810 30882
rect 77810 30830 77812 30882
rect 77756 30828 77812 30830
rect 76636 30322 76692 30324
rect 76636 30270 76638 30322
rect 76638 30270 76690 30322
rect 76690 30270 76692 30322
rect 76636 30268 76692 30270
rect 77308 30268 77364 30324
rect 76300 30098 76356 30100
rect 76300 30046 76302 30098
rect 76302 30046 76354 30098
rect 76354 30046 76356 30098
rect 76300 30044 76356 30046
rect 76972 29932 77028 29988
rect 76524 29036 76580 29092
rect 75404 28476 75460 28532
rect 75292 27804 75348 27860
rect 75180 27692 75236 27748
rect 73836 24780 73892 24836
rect 73612 23436 73668 23492
rect 73724 23212 73780 23268
rect 73164 22540 73220 22596
rect 73052 22316 73108 22372
rect 72492 21420 72548 21476
rect 71372 18620 71428 18676
rect 71596 19964 71652 20020
rect 71036 17836 71092 17892
rect 71148 17388 71204 17444
rect 71484 17500 71540 17556
rect 71372 17388 71428 17444
rect 71372 17106 71428 17108
rect 71372 17054 71374 17106
rect 71374 17054 71426 17106
rect 71426 17054 71428 17106
rect 71372 17052 71428 17054
rect 70700 16940 70756 16996
rect 71596 16940 71652 16996
rect 71484 16716 71540 16772
rect 71820 19180 71876 19236
rect 71932 20860 71988 20916
rect 71260 16492 71316 16548
rect 71036 14642 71092 14644
rect 71036 14590 71038 14642
rect 71038 14590 71090 14642
rect 71090 14590 71092 14642
rect 71036 14588 71092 14590
rect 71148 13858 71204 13860
rect 71148 13806 71150 13858
rect 71150 13806 71202 13858
rect 71202 13806 71204 13858
rect 71148 13804 71204 13806
rect 70588 13692 70644 13748
rect 69468 9996 69524 10052
rect 70812 12290 70868 12292
rect 70812 12238 70814 12290
rect 70814 12238 70866 12290
rect 70866 12238 70868 12290
rect 70812 12236 70868 12238
rect 70252 11228 70308 11284
rect 71820 18620 71876 18676
rect 71820 16492 71876 16548
rect 71932 16044 71988 16100
rect 71260 10892 71316 10948
rect 70140 10668 70196 10724
rect 70476 10668 70532 10724
rect 69916 10444 69972 10500
rect 69804 9884 69860 9940
rect 69244 8988 69300 9044
rect 69916 9042 69972 9044
rect 69916 8990 69918 9042
rect 69918 8990 69970 9042
rect 69970 8990 69972 9042
rect 69916 8988 69972 8990
rect 70364 9042 70420 9044
rect 70364 8990 70366 9042
rect 70366 8990 70418 9042
rect 70418 8990 70420 9042
rect 70364 8988 70420 8990
rect 68460 8540 68516 8596
rect 68832 8650 68888 8652
rect 68832 8598 68834 8650
rect 68834 8598 68886 8650
rect 68886 8598 68888 8650
rect 68832 8596 68888 8598
rect 68936 8650 68992 8652
rect 68936 8598 68938 8650
rect 68938 8598 68990 8650
rect 68990 8598 68992 8650
rect 68936 8596 68992 8598
rect 69040 8650 69096 8652
rect 69040 8598 69042 8650
rect 69042 8598 69094 8650
rect 69094 8598 69096 8650
rect 69040 8596 69096 8598
rect 69244 8428 69300 8484
rect 67116 8370 67172 8372
rect 67116 8318 67118 8370
rect 67118 8318 67170 8370
rect 67170 8318 67172 8370
rect 67116 8316 67172 8318
rect 68908 7196 68964 7252
rect 68832 7082 68888 7084
rect 68832 7030 68834 7082
rect 68834 7030 68886 7082
rect 68886 7030 68888 7082
rect 68832 7028 68888 7030
rect 68936 7082 68992 7084
rect 68936 7030 68938 7082
rect 68938 7030 68990 7082
rect 68990 7030 68992 7082
rect 68936 7028 68992 7030
rect 69040 7082 69096 7084
rect 69040 7030 69042 7082
rect 69042 7030 69094 7082
rect 69094 7030 69096 7082
rect 69040 7028 69096 7030
rect 69020 6578 69076 6580
rect 69020 6526 69022 6578
rect 69022 6526 69074 6578
rect 69074 6526 69076 6578
rect 69020 6524 69076 6526
rect 65884 5906 65940 5908
rect 65884 5854 65886 5906
rect 65886 5854 65938 5906
rect 65938 5854 65940 5906
rect 65884 5852 65940 5854
rect 65772 5122 65828 5124
rect 65772 5070 65774 5122
rect 65774 5070 65826 5122
rect 65826 5070 65828 5122
rect 65772 5068 65828 5070
rect 65548 5010 65604 5012
rect 65548 4958 65550 5010
rect 65550 4958 65602 5010
rect 65602 4958 65604 5010
rect 65548 4956 65604 4958
rect 65996 4956 66052 5012
rect 66332 4956 66388 5012
rect 66332 4172 66388 4228
rect 68684 6412 68740 6468
rect 69916 7644 69972 7700
rect 69580 6636 69636 6692
rect 69692 7196 69748 7252
rect 69692 6748 69748 6804
rect 69356 6466 69412 6468
rect 69356 6414 69358 6466
rect 69358 6414 69410 6466
rect 69410 6414 69412 6466
rect 69356 6412 69412 6414
rect 69916 7308 69972 7364
rect 71820 15036 71876 15092
rect 71820 14530 71876 14532
rect 71820 14478 71822 14530
rect 71822 14478 71874 14530
rect 71874 14478 71876 14530
rect 71820 14476 71876 14478
rect 71708 13746 71764 13748
rect 71708 13694 71710 13746
rect 71710 13694 71762 13746
rect 71762 13694 71764 13746
rect 71708 13692 71764 13694
rect 71372 9938 71428 9940
rect 71372 9886 71374 9938
rect 71374 9886 71426 9938
rect 71426 9886 71428 9938
rect 71372 9884 71428 9886
rect 71708 10556 71764 10612
rect 70700 9772 70756 9828
rect 70476 6524 70532 6580
rect 69804 6412 69860 6468
rect 68684 5852 68740 5908
rect 69580 6188 69636 6244
rect 68460 5740 68516 5796
rect 67228 5122 67284 5124
rect 67228 5070 67230 5122
rect 67230 5070 67282 5122
rect 67282 5070 67284 5122
rect 67228 5068 67284 5070
rect 67900 5122 67956 5124
rect 67900 5070 67902 5122
rect 67902 5070 67954 5122
rect 67954 5070 67956 5122
rect 67900 5068 67956 5070
rect 67116 4956 67172 5012
rect 62412 3612 62468 3668
rect 64764 3666 64820 3668
rect 64764 3614 64766 3666
rect 64766 3614 64818 3666
rect 64818 3614 64820 3666
rect 64764 3612 64820 3614
rect 67676 5010 67732 5012
rect 67676 4958 67678 5010
rect 67678 4958 67730 5010
rect 67730 4958 67732 5010
rect 67676 4956 67732 4958
rect 69356 5794 69412 5796
rect 69356 5742 69358 5794
rect 69358 5742 69410 5794
rect 69410 5742 69412 5794
rect 69356 5740 69412 5742
rect 68832 5514 68888 5516
rect 68832 5462 68834 5514
rect 68834 5462 68886 5514
rect 68886 5462 68888 5514
rect 68832 5460 68888 5462
rect 68936 5514 68992 5516
rect 68936 5462 68938 5514
rect 68938 5462 68990 5514
rect 68990 5462 68992 5514
rect 68936 5460 68992 5462
rect 69040 5514 69096 5516
rect 69040 5462 69042 5514
rect 69042 5462 69094 5514
rect 69094 5462 69096 5514
rect 69040 5460 69096 5462
rect 69020 5122 69076 5124
rect 69020 5070 69022 5122
rect 69022 5070 69074 5122
rect 69074 5070 69076 5122
rect 69020 5068 69076 5070
rect 68572 5010 68628 5012
rect 68572 4958 68574 5010
rect 68574 4958 68626 5010
rect 68626 4958 68628 5010
rect 68572 4956 68628 4958
rect 68124 4226 68180 4228
rect 68124 4174 68126 4226
rect 68126 4174 68178 4226
rect 68178 4174 68180 4226
rect 68124 4172 68180 4174
rect 68236 4060 68292 4116
rect 67900 2828 67956 2884
rect 69692 4396 69748 4452
rect 70028 6188 70084 6244
rect 69916 5740 69972 5796
rect 69468 4114 69524 4116
rect 69468 4062 69470 4114
rect 69470 4062 69522 4114
rect 69522 4062 69524 4114
rect 69468 4060 69524 4062
rect 68832 3946 68888 3948
rect 68832 3894 68834 3946
rect 68834 3894 68886 3946
rect 68886 3894 68888 3946
rect 68832 3892 68888 3894
rect 68936 3946 68992 3948
rect 68936 3894 68938 3946
rect 68938 3894 68990 3946
rect 68990 3894 68992 3946
rect 68936 3892 68992 3894
rect 69040 3946 69096 3948
rect 69040 3894 69042 3946
rect 69042 3894 69094 3946
rect 69094 3894 69096 3946
rect 69040 3892 69096 3894
rect 68684 3724 68740 3780
rect 70252 6300 70308 6356
rect 71036 9324 71092 9380
rect 70700 6690 70756 6692
rect 70700 6638 70702 6690
rect 70702 6638 70754 6690
rect 70754 6638 70756 6690
rect 70700 6636 70756 6638
rect 70588 6188 70644 6244
rect 70700 6076 70756 6132
rect 70588 5628 70644 5684
rect 70924 6412 70980 6468
rect 70924 5794 70980 5796
rect 70924 5742 70926 5794
rect 70926 5742 70978 5794
rect 70978 5742 70980 5794
rect 70924 5740 70980 5742
rect 70812 5404 70868 5460
rect 70364 4956 70420 5012
rect 71260 8316 71316 8372
rect 71148 7644 71204 7700
rect 71484 8146 71540 8148
rect 71484 8094 71486 8146
rect 71486 8094 71538 8146
rect 71538 8094 71540 8146
rect 71484 8092 71540 8094
rect 71260 6748 71316 6804
rect 71484 7362 71540 7364
rect 71484 7310 71486 7362
rect 71486 7310 71538 7362
rect 71538 7310 71540 7362
rect 71484 7308 71540 7310
rect 71372 6188 71428 6244
rect 71036 4508 71092 4564
rect 69916 2604 69972 2660
rect 72044 9772 72100 9828
rect 72716 21084 72772 21140
rect 72828 21980 72884 22036
rect 72940 21586 72996 21588
rect 72940 21534 72942 21586
rect 72942 21534 72994 21586
rect 72994 21534 72996 21586
rect 72940 21532 72996 21534
rect 72268 18396 72324 18452
rect 72828 20690 72884 20692
rect 72828 20638 72830 20690
rect 72830 20638 72882 20690
rect 72882 20638 72884 20690
rect 72828 20636 72884 20638
rect 73500 22540 73556 22596
rect 73500 21810 73556 21812
rect 73500 21758 73502 21810
rect 73502 21758 73554 21810
rect 73554 21758 73556 21810
rect 73500 21756 73556 21758
rect 74060 23436 74116 23492
rect 72492 18732 72548 18788
rect 72604 19068 72660 19124
rect 72268 17666 72324 17668
rect 72268 17614 72270 17666
rect 72270 17614 72322 17666
rect 72322 17614 72324 17666
rect 72268 17612 72324 17614
rect 72268 16994 72324 16996
rect 72268 16942 72270 16994
rect 72270 16942 72322 16994
rect 72322 16942 72324 16994
rect 72268 16940 72324 16942
rect 73276 19122 73332 19124
rect 73276 19070 73278 19122
rect 73278 19070 73330 19122
rect 73330 19070 73332 19122
rect 73276 19068 73332 19070
rect 73836 22092 73892 22148
rect 73724 21698 73780 21700
rect 73724 21646 73726 21698
rect 73726 21646 73778 21698
rect 73778 21646 73780 21698
rect 73724 21644 73780 21646
rect 73724 20802 73780 20804
rect 73724 20750 73726 20802
rect 73726 20750 73778 20802
rect 73778 20750 73780 20802
rect 73724 20748 73780 20750
rect 74620 24946 74676 24948
rect 74620 24894 74622 24946
rect 74622 24894 74674 24946
rect 74674 24894 74676 24946
rect 74620 24892 74676 24894
rect 74284 23548 74340 23604
rect 75292 26124 75348 26180
rect 75292 25452 75348 25508
rect 75628 26460 75684 26516
rect 75516 25452 75572 25508
rect 76636 25730 76692 25732
rect 76636 25678 76638 25730
rect 76638 25678 76690 25730
rect 76690 25678 76692 25730
rect 76636 25676 76692 25678
rect 77084 26178 77140 26180
rect 77084 26126 77086 26178
rect 77086 26126 77138 26178
rect 77138 26126 77140 26178
rect 77084 26124 77140 26126
rect 77980 30268 78036 30324
rect 78492 29818 78548 29820
rect 78492 29766 78494 29818
rect 78494 29766 78546 29818
rect 78546 29766 78548 29818
rect 78492 29764 78548 29766
rect 78596 29818 78652 29820
rect 78596 29766 78598 29818
rect 78598 29766 78650 29818
rect 78650 29766 78652 29818
rect 78596 29764 78652 29766
rect 78700 29818 78756 29820
rect 78700 29766 78702 29818
rect 78702 29766 78754 29818
rect 78754 29766 78756 29818
rect 78700 29764 78756 29766
rect 78492 28250 78548 28252
rect 78492 28198 78494 28250
rect 78494 28198 78546 28250
rect 78546 28198 78548 28250
rect 78492 28196 78548 28198
rect 78596 28250 78652 28252
rect 78596 28198 78598 28250
rect 78598 28198 78650 28250
rect 78650 28198 78652 28250
rect 78596 28196 78652 28198
rect 78700 28250 78756 28252
rect 78700 28198 78702 28250
rect 78702 28198 78754 28250
rect 78754 28198 78756 28250
rect 78700 28196 78756 28198
rect 77756 26908 77812 26964
rect 78492 26682 78548 26684
rect 78492 26630 78494 26682
rect 78494 26630 78546 26682
rect 78546 26630 78548 26682
rect 78492 26628 78548 26630
rect 78596 26682 78652 26684
rect 78596 26630 78598 26682
rect 78598 26630 78650 26682
rect 78650 26630 78652 26682
rect 78596 26628 78652 26630
rect 78700 26682 78756 26684
rect 78700 26630 78702 26682
rect 78702 26630 78754 26682
rect 78754 26630 78756 26682
rect 78700 26628 78756 26630
rect 77980 26012 78036 26068
rect 77308 25676 77364 25732
rect 77980 25676 78036 25732
rect 75404 23660 75460 23716
rect 74844 23436 74900 23492
rect 76860 25452 76916 25508
rect 74172 22092 74228 22148
rect 74060 21868 74116 21924
rect 76412 23042 76468 23044
rect 76412 22990 76414 23042
rect 76414 22990 76466 23042
rect 76466 22990 76468 23042
rect 76412 22988 76468 22990
rect 75628 22764 75684 22820
rect 74844 21980 74900 22036
rect 74732 21756 74788 21812
rect 74844 21532 74900 21588
rect 73948 21420 74004 21476
rect 73164 17500 73220 17556
rect 73388 17836 73444 17892
rect 72828 17052 72884 17108
rect 73164 15202 73220 15204
rect 73164 15150 73166 15202
rect 73166 15150 73218 15202
rect 73218 15150 73220 15202
rect 73164 15148 73220 15150
rect 72492 13692 72548 13748
rect 73948 18620 74004 18676
rect 73724 16268 73780 16324
rect 73836 16098 73892 16100
rect 73836 16046 73838 16098
rect 73838 16046 73890 16098
rect 73890 16046 73892 16098
rect 73836 16044 73892 16046
rect 74396 18172 74452 18228
rect 74620 17388 74676 17444
rect 74620 16828 74676 16884
rect 74396 16098 74452 16100
rect 74396 16046 74398 16098
rect 74398 16046 74450 16098
rect 74450 16046 74452 16098
rect 74396 16044 74452 16046
rect 74060 15260 74116 15316
rect 74396 15148 74452 15204
rect 73500 15036 73556 15092
rect 74172 14924 74228 14980
rect 73276 13858 73332 13860
rect 73276 13806 73278 13858
rect 73278 13806 73330 13858
rect 73330 13806 73332 13858
rect 73276 13804 73332 13806
rect 73388 13746 73444 13748
rect 73388 13694 73390 13746
rect 73390 13694 73442 13746
rect 73442 13694 73444 13746
rect 73388 13692 73444 13694
rect 72380 12236 72436 12292
rect 72604 11282 72660 11284
rect 72604 11230 72606 11282
rect 72606 11230 72658 11282
rect 72658 11230 72660 11282
rect 72604 11228 72660 11230
rect 72268 9324 72324 9380
rect 72380 10892 72436 10948
rect 72604 10668 72660 10724
rect 72716 10444 72772 10500
rect 72380 10108 72436 10164
rect 72492 9772 72548 9828
rect 72156 8316 72212 8372
rect 72380 8092 72436 8148
rect 73276 12738 73332 12740
rect 73276 12686 73278 12738
rect 73278 12686 73330 12738
rect 73330 12686 73332 12738
rect 73276 12684 73332 12686
rect 72940 9996 72996 10052
rect 72940 9660 72996 9716
rect 73052 12572 73108 12628
rect 72268 7308 72324 7364
rect 72940 7308 72996 7364
rect 73388 10668 73444 10724
rect 73724 13804 73780 13860
rect 73948 12962 74004 12964
rect 73948 12910 73950 12962
rect 73950 12910 74002 12962
rect 74002 12910 74004 12962
rect 73948 12908 74004 12910
rect 74620 14924 74676 14980
rect 74732 15260 74788 15316
rect 74508 14028 74564 14084
rect 74620 13916 74676 13972
rect 74396 13858 74452 13860
rect 74396 13806 74398 13858
rect 74398 13806 74450 13858
rect 74450 13806 74452 13858
rect 74396 13804 74452 13806
rect 75180 21868 75236 21924
rect 76300 21756 76356 21812
rect 75852 21698 75908 21700
rect 75852 21646 75854 21698
rect 75854 21646 75906 21698
rect 75906 21646 75908 21698
rect 75852 21644 75908 21646
rect 75068 20748 75124 20804
rect 75292 20188 75348 20244
rect 75740 20188 75796 20244
rect 74956 19346 75012 19348
rect 74956 19294 74958 19346
rect 74958 19294 75010 19346
rect 75010 19294 75012 19346
rect 74956 19292 75012 19294
rect 76188 19404 76244 19460
rect 75628 19122 75684 19124
rect 75628 19070 75630 19122
rect 75630 19070 75682 19122
rect 75682 19070 75684 19122
rect 75628 19068 75684 19070
rect 75292 19010 75348 19012
rect 75292 18958 75294 19010
rect 75294 18958 75346 19010
rect 75346 18958 75348 19010
rect 75292 18956 75348 18958
rect 75068 18620 75124 18676
rect 75292 18396 75348 18452
rect 76412 17836 76468 17892
rect 75516 17778 75572 17780
rect 75516 17726 75518 17778
rect 75518 17726 75570 17778
rect 75570 17726 75572 17778
rect 75516 17724 75572 17726
rect 74956 17612 75012 17668
rect 75180 17442 75236 17444
rect 75180 17390 75182 17442
rect 75182 17390 75234 17442
rect 75234 17390 75236 17442
rect 75180 17388 75236 17390
rect 76188 17442 76244 17444
rect 76188 17390 76190 17442
rect 76190 17390 76242 17442
rect 76242 17390 76244 17442
rect 76188 17388 76244 17390
rect 76636 22764 76692 22820
rect 76972 22652 77028 22708
rect 77420 25394 77476 25396
rect 77420 25342 77422 25394
rect 77422 25342 77474 25394
rect 77474 25342 77476 25394
rect 77420 25340 77476 25342
rect 78204 25340 78260 25396
rect 78492 25114 78548 25116
rect 78492 25062 78494 25114
rect 78494 25062 78546 25114
rect 78546 25062 78548 25114
rect 78492 25060 78548 25062
rect 78596 25114 78652 25116
rect 78596 25062 78598 25114
rect 78598 25062 78650 25114
rect 78650 25062 78652 25114
rect 78596 25060 78652 25062
rect 78700 25114 78756 25116
rect 78700 25062 78702 25114
rect 78702 25062 78754 25114
rect 78754 25062 78756 25114
rect 78700 25060 78756 25062
rect 78492 23546 78548 23548
rect 78492 23494 78494 23546
rect 78494 23494 78546 23546
rect 78546 23494 78548 23546
rect 78492 23492 78548 23494
rect 78596 23546 78652 23548
rect 78596 23494 78598 23546
rect 78598 23494 78650 23546
rect 78650 23494 78652 23546
rect 78596 23492 78652 23494
rect 78700 23546 78756 23548
rect 78700 23494 78702 23546
rect 78702 23494 78754 23546
rect 78754 23494 78756 23546
rect 78700 23492 78756 23494
rect 77196 22988 77252 23044
rect 77644 22764 77700 22820
rect 77980 22652 78036 22708
rect 77868 21644 77924 21700
rect 78492 21978 78548 21980
rect 78492 21926 78494 21978
rect 78494 21926 78546 21978
rect 78546 21926 78548 21978
rect 78492 21924 78548 21926
rect 78596 21978 78652 21980
rect 78596 21926 78598 21978
rect 78598 21926 78650 21978
rect 78650 21926 78652 21978
rect 78596 21924 78652 21926
rect 78700 21978 78756 21980
rect 78700 21926 78702 21978
rect 78702 21926 78754 21978
rect 78754 21926 78756 21978
rect 78700 21924 78756 21926
rect 77980 21084 78036 21140
rect 78492 20410 78548 20412
rect 78492 20358 78494 20410
rect 78494 20358 78546 20410
rect 78546 20358 78548 20410
rect 78492 20356 78548 20358
rect 78596 20410 78652 20412
rect 78596 20358 78598 20410
rect 78598 20358 78650 20410
rect 78650 20358 78652 20410
rect 78596 20356 78652 20358
rect 78700 20410 78756 20412
rect 78700 20358 78702 20410
rect 78702 20358 78754 20410
rect 78754 20358 78756 20410
rect 78700 20356 78756 20358
rect 76860 19292 76916 19348
rect 78092 19346 78148 19348
rect 78092 19294 78094 19346
rect 78094 19294 78146 19346
rect 78146 19294 78148 19346
rect 78092 19292 78148 19294
rect 77644 19122 77700 19124
rect 77644 19070 77646 19122
rect 77646 19070 77698 19122
rect 77698 19070 77700 19122
rect 77644 19068 77700 19070
rect 77196 19010 77252 19012
rect 77196 18958 77198 19010
rect 77198 18958 77250 19010
rect 77250 18958 77252 19010
rect 77196 18956 77252 18958
rect 78492 18842 78548 18844
rect 78492 18790 78494 18842
rect 78494 18790 78546 18842
rect 78546 18790 78548 18842
rect 78492 18788 78548 18790
rect 78596 18842 78652 18844
rect 78596 18790 78598 18842
rect 78598 18790 78650 18842
rect 78650 18790 78652 18842
rect 78596 18788 78652 18790
rect 78700 18842 78756 18844
rect 78700 18790 78702 18842
rect 78702 18790 78754 18842
rect 78754 18790 78756 18842
rect 78700 18788 78756 18790
rect 77308 17836 77364 17892
rect 76636 17724 76692 17780
rect 77196 17612 77252 17668
rect 77308 17388 77364 17444
rect 78492 17274 78548 17276
rect 78492 17222 78494 17274
rect 78494 17222 78546 17274
rect 78546 17222 78548 17274
rect 78492 17220 78548 17222
rect 78596 17274 78652 17276
rect 78596 17222 78598 17274
rect 78598 17222 78650 17274
rect 78650 17222 78652 17274
rect 78596 17220 78652 17222
rect 78700 17274 78756 17276
rect 78700 17222 78702 17274
rect 78702 17222 78754 17274
rect 78754 17222 78756 17274
rect 78700 17220 78756 17222
rect 76412 16210 76468 16212
rect 76412 16158 76414 16210
rect 76414 16158 76466 16210
rect 76466 16158 76468 16210
rect 76412 16156 76468 16158
rect 76972 16156 77028 16212
rect 76188 15036 76244 15092
rect 75628 14530 75684 14532
rect 75628 14478 75630 14530
rect 75630 14478 75682 14530
rect 75682 14478 75684 14530
rect 75628 14476 75684 14478
rect 76860 14476 76916 14532
rect 76300 14364 76356 14420
rect 74172 12572 74228 12628
rect 75628 12738 75684 12740
rect 75628 12686 75630 12738
rect 75630 12686 75682 12738
rect 75682 12686 75684 12738
rect 75628 12684 75684 12686
rect 75628 11394 75684 11396
rect 75628 11342 75630 11394
rect 75630 11342 75682 11394
rect 75682 11342 75684 11394
rect 75628 11340 75684 11342
rect 74620 11170 74676 11172
rect 74620 11118 74622 11170
rect 74622 11118 74674 11170
rect 74674 11118 74676 11170
rect 74620 11116 74676 11118
rect 73388 10220 73444 10276
rect 74172 10668 74228 10724
rect 74060 10220 74116 10276
rect 73612 10108 73668 10164
rect 73500 9826 73556 9828
rect 73500 9774 73502 9826
rect 73502 9774 73554 9826
rect 73554 9774 73556 9826
rect 73500 9772 73556 9774
rect 73612 9884 73668 9940
rect 73500 9436 73556 9492
rect 73276 9324 73332 9380
rect 73836 9324 73892 9380
rect 74060 9436 74116 9492
rect 73164 7644 73220 7700
rect 73276 7362 73332 7364
rect 73276 7310 73278 7362
rect 73278 7310 73330 7362
rect 73330 7310 73332 7362
rect 73276 7308 73332 7310
rect 71596 6524 71652 6580
rect 71708 6300 71764 6356
rect 72156 6636 72212 6692
rect 72268 5740 72324 5796
rect 72940 6130 72996 6132
rect 72940 6078 72942 6130
rect 72942 6078 72994 6130
rect 72994 6078 72996 6130
rect 72940 6076 72996 6078
rect 75516 10498 75572 10500
rect 75516 10446 75518 10498
rect 75518 10446 75570 10498
rect 75570 10446 75572 10498
rect 75516 10444 75572 10446
rect 74284 9996 74340 10052
rect 74172 6076 74228 6132
rect 72380 5404 72436 5460
rect 71484 2492 71540 2548
rect 72156 3500 72212 3556
rect 76076 10332 76132 10388
rect 76524 14306 76580 14308
rect 76524 14254 76526 14306
rect 76526 14254 76578 14306
rect 76578 14254 76580 14306
rect 76524 14252 76580 14254
rect 76860 13858 76916 13860
rect 76860 13806 76862 13858
rect 76862 13806 76914 13858
rect 76914 13806 76916 13858
rect 76860 13804 76916 13806
rect 77196 14418 77252 14420
rect 77196 14366 77198 14418
rect 77198 14366 77250 14418
rect 77250 14366 77252 14418
rect 77196 14364 77252 14366
rect 77644 14418 77700 14420
rect 77644 14366 77646 14418
rect 77646 14366 77698 14418
rect 77698 14366 77700 14418
rect 77644 14364 77700 14366
rect 77980 16156 78036 16212
rect 78492 15706 78548 15708
rect 78492 15654 78494 15706
rect 78494 15654 78546 15706
rect 78546 15654 78548 15706
rect 78492 15652 78548 15654
rect 78596 15706 78652 15708
rect 78596 15654 78598 15706
rect 78598 15654 78650 15706
rect 78650 15654 78652 15706
rect 78596 15652 78652 15654
rect 78700 15706 78756 15708
rect 78700 15654 78702 15706
rect 78702 15654 78754 15706
rect 78754 15654 78756 15706
rect 78700 15652 78756 15654
rect 77756 14252 77812 14308
rect 78492 14138 78548 14140
rect 78492 14086 78494 14138
rect 78494 14086 78546 14138
rect 78546 14086 78548 14138
rect 78492 14084 78548 14086
rect 78596 14138 78652 14140
rect 78596 14086 78598 14138
rect 78598 14086 78650 14138
rect 78650 14086 78652 14138
rect 78596 14084 78652 14086
rect 78700 14138 78756 14140
rect 78700 14086 78702 14138
rect 78702 14086 78754 14138
rect 78754 14086 78756 14138
rect 78700 14084 78756 14086
rect 76860 12684 76916 12740
rect 76524 11564 76580 11620
rect 76412 10780 76468 10836
rect 76748 11340 76804 11396
rect 76972 10780 77028 10836
rect 76300 9548 76356 9604
rect 76972 7868 77028 7924
rect 76972 7196 77028 7252
rect 72604 3554 72660 3556
rect 72604 3502 72606 3554
rect 72606 3502 72658 3554
rect 72658 3502 72660 3554
rect 72604 3500 72660 3502
rect 75516 1372 75572 1428
rect 78492 12570 78548 12572
rect 78492 12518 78494 12570
rect 78494 12518 78546 12570
rect 78546 12518 78548 12570
rect 78492 12516 78548 12518
rect 78596 12570 78652 12572
rect 78596 12518 78598 12570
rect 78598 12518 78650 12570
rect 78650 12518 78652 12570
rect 78596 12516 78652 12518
rect 78700 12570 78756 12572
rect 78700 12518 78702 12570
rect 78702 12518 78754 12570
rect 78754 12518 78756 12570
rect 78700 12516 78756 12518
rect 78492 11002 78548 11004
rect 78492 10950 78494 11002
rect 78494 10950 78546 11002
rect 78546 10950 78548 11002
rect 78492 10948 78548 10950
rect 78596 11002 78652 11004
rect 78596 10950 78598 11002
rect 78598 10950 78650 11002
rect 78650 10950 78652 11002
rect 78596 10948 78652 10950
rect 78700 11002 78756 11004
rect 78700 10950 78702 11002
rect 78702 10950 78754 11002
rect 78754 10950 78756 11002
rect 78700 10948 78756 10950
rect 77196 7308 77252 7364
rect 77644 10332 77700 10388
rect 78492 9434 78548 9436
rect 78492 9382 78494 9434
rect 78494 9382 78546 9434
rect 78546 9382 78548 9434
rect 78492 9380 78548 9382
rect 78596 9434 78652 9436
rect 78596 9382 78598 9434
rect 78598 9382 78650 9434
rect 78650 9382 78652 9434
rect 78596 9380 78652 9382
rect 78700 9434 78756 9436
rect 78700 9382 78702 9434
rect 78702 9382 78754 9434
rect 78754 9382 78756 9434
rect 78700 9380 78756 9382
rect 77980 8818 78036 8820
rect 77980 8766 77982 8818
rect 77982 8766 78034 8818
rect 78034 8766 78036 8818
rect 77980 8764 78036 8766
rect 78492 7866 78548 7868
rect 78492 7814 78494 7866
rect 78494 7814 78546 7866
rect 78546 7814 78548 7866
rect 78492 7812 78548 7814
rect 78596 7866 78652 7868
rect 78596 7814 78598 7866
rect 78598 7814 78650 7866
rect 78650 7814 78652 7866
rect 78596 7812 78652 7814
rect 78700 7866 78756 7868
rect 78700 7814 78702 7866
rect 78702 7814 78754 7866
rect 78754 7814 78756 7866
rect 78700 7812 78756 7814
rect 78492 6298 78548 6300
rect 78492 6246 78494 6298
rect 78494 6246 78546 6298
rect 78546 6246 78548 6298
rect 78492 6244 78548 6246
rect 78596 6298 78652 6300
rect 78596 6246 78598 6298
rect 78598 6246 78650 6298
rect 78650 6246 78652 6298
rect 78596 6244 78652 6246
rect 78700 6298 78756 6300
rect 78700 6246 78702 6298
rect 78702 6246 78754 6298
rect 78754 6246 78756 6298
rect 78700 6244 78756 6246
rect 77980 6076 78036 6132
rect 78492 4730 78548 4732
rect 78492 4678 78494 4730
rect 78494 4678 78546 4730
rect 78546 4678 78548 4730
rect 78492 4676 78548 4678
rect 78596 4730 78652 4732
rect 78596 4678 78598 4730
rect 78598 4678 78650 4730
rect 78650 4678 78652 4730
rect 78596 4676 78652 4678
rect 78700 4730 78756 4732
rect 78700 4678 78702 4730
rect 78702 4678 78754 4730
rect 78754 4678 78756 4730
rect 78700 4676 78756 4678
rect 77980 3836 78036 3892
rect 77084 3276 77140 3332
rect 78492 3162 78548 3164
rect 78492 3110 78494 3162
rect 78494 3110 78546 3162
rect 78546 3110 78548 3162
rect 78492 3108 78548 3110
rect 78596 3162 78652 3164
rect 78596 3110 78598 3162
rect 78598 3110 78650 3162
rect 78650 3110 78652 3162
rect 78596 3108 78652 3110
rect 78700 3162 78756 3164
rect 78700 3110 78702 3162
rect 78702 3110 78754 3162
rect 78754 3110 78756 3162
rect 78700 3108 78756 3110
<< metal3 >>
rect 0 38388 800 38416
rect 79200 38388 80000 38416
rect 0 38332 3388 38388
rect 3444 38332 3454 38388
rect 73938 38332 73948 38388
rect 74004 38332 80000 38388
rect 0 38304 800 38332
rect 79200 38304 80000 38332
rect 14466 37548 14476 37604
rect 14532 37548 39564 37604
rect 39620 37548 39630 37604
rect 21634 37436 21644 37492
rect 21700 37436 41580 37492
rect 41636 37436 41646 37492
rect 20850 37324 20860 37380
rect 20916 37324 42476 37380
rect 42532 37324 42542 37380
rect 34962 37212 34972 37268
rect 35028 37212 44380 37268
rect 44436 37212 44446 37268
rect 23548 37100 52556 37156
rect 52612 37100 52622 37156
rect 23548 36932 23604 37100
rect 26338 36988 26348 37044
rect 26404 36988 29596 37044
rect 29652 36988 72772 37044
rect 22082 36876 22092 36932
rect 22148 36876 23604 36932
rect 72716 36932 72772 36988
rect 72716 36876 73724 36932
rect 73780 36876 74060 36932
rect 74116 36876 74126 36932
rect 10862 36820 10872 36876
rect 10928 36820 10976 36876
rect 11032 36820 11080 36876
rect 11136 36820 11146 36876
rect 30182 36820 30192 36876
rect 30248 36820 30296 36876
rect 30352 36820 30400 36876
rect 30456 36820 30466 36876
rect 49502 36820 49512 36876
rect 49568 36820 49616 36876
rect 49672 36820 49720 36876
rect 49776 36820 49786 36876
rect 68822 36820 68832 36876
rect 68888 36820 68936 36876
rect 68992 36820 69040 36876
rect 69096 36820 69106 36876
rect 19618 36652 19628 36708
rect 19684 36652 52444 36708
rect 52500 36652 52510 36708
rect 53330 36652 53340 36708
rect 53396 36652 56028 36708
rect 56084 36652 56094 36708
rect 67172 36652 68348 36708
rect 68404 36652 68414 36708
rect 73042 36652 73052 36708
rect 73108 36652 75068 36708
rect 75124 36652 75134 36708
rect 67172 36596 67228 36652
rect 29138 36540 29148 36596
rect 29204 36540 31164 36596
rect 31220 36540 31230 36596
rect 31602 36540 31612 36596
rect 31668 36540 32844 36596
rect 32900 36540 32910 36596
rect 38612 36540 67228 36596
rect 38612 36484 38668 36540
rect 16370 36428 16380 36484
rect 16436 36428 17052 36484
rect 17108 36428 17118 36484
rect 24770 36428 24780 36484
rect 24836 36428 26236 36484
rect 26292 36428 27356 36484
rect 27412 36428 27422 36484
rect 28242 36428 28252 36484
rect 28308 36428 38668 36484
rect 43026 36428 43036 36484
rect 43092 36428 45836 36484
rect 45892 36428 45902 36484
rect 52322 36428 52332 36484
rect 52388 36428 62636 36484
rect 62692 36428 62702 36484
rect 65874 36428 65884 36484
rect 65940 36428 66556 36484
rect 66612 36428 66622 36484
rect 28252 36372 28308 36428
rect 7298 36316 7308 36372
rect 7364 36316 22092 36372
rect 22148 36316 22158 36372
rect 24098 36316 24108 36372
rect 24164 36316 27020 36372
rect 27076 36316 28308 36372
rect 28802 36316 28812 36372
rect 28868 36316 29820 36372
rect 29876 36316 72380 36372
rect 72436 36316 72446 36372
rect 13794 36204 13804 36260
rect 13860 36204 17724 36260
rect 17780 36204 17790 36260
rect 25330 36204 25340 36260
rect 25396 36204 28700 36260
rect 28756 36204 28766 36260
rect 28914 36204 28924 36260
rect 28980 36204 29372 36260
rect 29428 36204 29438 36260
rect 46274 36204 46284 36260
rect 46340 36204 50428 36260
rect 50484 36204 50494 36260
rect 56252 36204 70476 36260
rect 70532 36204 70812 36260
rect 70868 36204 70878 36260
rect 20522 36036 20532 36092
rect 20588 36036 20636 36092
rect 20692 36036 20740 36092
rect 20796 36036 20806 36092
rect 39842 36036 39852 36092
rect 39908 36036 39956 36092
rect 40012 36036 40060 36092
rect 40116 36036 40126 36092
rect 56252 36036 56308 36204
rect 59162 36036 59172 36092
rect 59228 36036 59276 36092
rect 59332 36036 59380 36092
rect 59436 36036 59446 36092
rect 78482 36036 78492 36092
rect 78548 36036 78596 36092
rect 78652 36036 78700 36092
rect 78756 36036 78766 36092
rect 44492 35980 56308 36036
rect 0 35924 800 35952
rect 44492 35924 44548 35980
rect 79200 35924 80000 35952
rect 0 35868 1932 35924
rect 1988 35868 1998 35924
rect 17266 35868 17276 35924
rect 17332 35868 27188 35924
rect 29474 35868 29484 35924
rect 29540 35868 44548 35924
rect 46274 35868 46284 35924
rect 46340 35868 46844 35924
rect 46900 35868 62188 35924
rect 63186 35868 63196 35924
rect 63252 35868 65436 35924
rect 65492 35868 65502 35924
rect 75506 35868 75516 35924
rect 75572 35868 76636 35924
rect 76692 35868 76702 35924
rect 76860 35868 80000 35924
rect 0 35840 800 35868
rect 27132 35812 27188 35868
rect 62132 35812 62188 35868
rect 76860 35812 76916 35868
rect 79200 35840 80000 35868
rect 14690 35756 14700 35812
rect 14756 35756 25900 35812
rect 25956 35756 27076 35812
rect 27132 35756 46228 35812
rect 48178 35756 48188 35812
rect 48244 35756 48972 35812
rect 49028 35756 52332 35812
rect 52388 35756 52398 35812
rect 62132 35756 63868 35812
rect 63924 35756 64428 35812
rect 64484 35756 64494 35812
rect 75058 35756 75068 35812
rect 75124 35756 76916 35812
rect 27020 35700 27076 35756
rect 21858 35644 21868 35700
rect 21924 35644 26348 35700
rect 26404 35644 26414 35700
rect 27020 35644 29484 35700
rect 29540 35644 29550 35700
rect 29932 35644 31276 35700
rect 31332 35644 33292 35700
rect 33348 35644 33358 35700
rect 29932 35588 29988 35644
rect 13234 35532 13244 35588
rect 13300 35532 15372 35588
rect 15428 35532 15438 35588
rect 29250 35532 29260 35588
rect 29316 35532 29988 35588
rect 30146 35532 30156 35588
rect 30212 35532 31948 35588
rect 32004 35532 32014 35588
rect 37538 35532 37548 35588
rect 37604 35532 37772 35588
rect 37828 35532 40572 35588
rect 40628 35532 40638 35588
rect 43250 35532 43260 35588
rect 43316 35532 44268 35588
rect 44324 35532 44334 35588
rect 16594 35420 16604 35476
rect 16660 35420 17052 35476
rect 17108 35420 18284 35476
rect 18340 35420 18956 35476
rect 19012 35420 28700 35476
rect 28756 35420 28766 35476
rect 29138 35420 29148 35476
rect 29204 35420 29596 35476
rect 29652 35420 29662 35476
rect 30482 35420 30492 35476
rect 30548 35420 32172 35476
rect 32228 35420 32238 35476
rect 33506 35420 33516 35476
rect 33572 35420 36540 35476
rect 36596 35420 36988 35476
rect 37044 35420 37054 35476
rect 37212 35420 45164 35476
rect 45220 35420 45230 35476
rect 32172 35364 32228 35420
rect 37212 35364 37268 35420
rect 46172 35364 46228 35756
rect 47618 35644 47628 35700
rect 47684 35644 49084 35700
rect 49140 35644 49150 35700
rect 50418 35644 50428 35700
rect 50484 35644 50988 35700
rect 51044 35644 54908 35700
rect 54964 35644 54974 35700
rect 57138 35644 57148 35700
rect 57204 35644 65884 35700
rect 65940 35644 65950 35700
rect 47954 35420 47964 35476
rect 48020 35420 48860 35476
rect 48916 35420 58044 35476
rect 58100 35420 61068 35476
rect 61124 35420 61134 35476
rect 12226 35308 12236 35364
rect 12292 35308 28756 35364
rect 29026 35308 29036 35364
rect 29092 35308 29372 35364
rect 29428 35308 29438 35364
rect 32172 35308 33068 35364
rect 33124 35308 33134 35364
rect 33618 35308 33628 35364
rect 33684 35308 37268 35364
rect 37324 35308 39228 35364
rect 39284 35308 39294 35364
rect 42130 35308 42140 35364
rect 42196 35308 44156 35364
rect 44212 35308 44222 35364
rect 46162 35308 46172 35364
rect 46228 35308 46238 35364
rect 67172 35308 67452 35364
rect 67508 35308 67518 35364
rect 10862 35252 10872 35308
rect 10928 35252 10976 35308
rect 11032 35252 11080 35308
rect 11136 35252 11146 35308
rect 28700 35252 28756 35308
rect 30182 35252 30192 35308
rect 30248 35252 30296 35308
rect 30352 35252 30400 35308
rect 30456 35252 30466 35308
rect 37324 35252 37380 35308
rect 49502 35252 49512 35308
rect 49568 35252 49616 35308
rect 49672 35252 49720 35308
rect 49776 35252 49786 35308
rect 67172 35252 67228 35308
rect 68822 35252 68832 35308
rect 68888 35252 68936 35308
rect 68992 35252 69040 35308
rect 69096 35252 69106 35308
rect 28690 35196 28700 35252
rect 28756 35196 28766 35252
rect 36754 35196 36764 35252
rect 36820 35196 37380 35252
rect 37874 35196 37884 35252
rect 37940 35196 38444 35252
rect 38500 35196 38510 35252
rect 38770 35196 38780 35252
rect 38836 35196 40236 35252
rect 40292 35196 40302 35252
rect 44370 35196 44380 35252
rect 44436 35196 45612 35252
rect 45668 35196 45678 35252
rect 50642 35196 50652 35252
rect 50708 35196 51324 35252
rect 51380 35196 51390 35252
rect 55794 35196 55804 35252
rect 55860 35196 60620 35252
rect 60676 35196 60686 35252
rect 65650 35196 65660 35252
rect 65716 35196 67228 35252
rect 2930 35084 2940 35140
rect 2996 35084 3948 35140
rect 4004 35084 4014 35140
rect 21522 35084 21532 35140
rect 21588 35084 25004 35140
rect 25060 35084 25340 35140
rect 25396 35084 25406 35140
rect 26562 35084 26572 35140
rect 26628 35084 27356 35140
rect 27412 35084 30996 35140
rect 36866 35084 36876 35140
rect 36932 35084 38892 35140
rect 38948 35084 38958 35140
rect 39106 35084 39116 35140
rect 39172 35084 40460 35140
rect 40516 35084 40526 35140
rect 45836 35084 47908 35140
rect 48402 35084 48412 35140
rect 48468 35084 52220 35140
rect 52276 35084 52286 35140
rect 53106 35084 53116 35140
rect 53172 35084 57148 35140
rect 57204 35084 57214 35140
rect 58258 35084 58268 35140
rect 58324 35084 64092 35140
rect 64148 35084 64158 35140
rect 68114 35084 68124 35140
rect 68180 35084 69356 35140
rect 69412 35084 69422 35140
rect 30940 35028 30996 35084
rect 45836 35028 45892 35084
rect 1810 34972 1820 35028
rect 1876 34972 3500 35028
rect 3556 34972 3566 35028
rect 9874 34972 9884 35028
rect 9940 34972 27804 35028
rect 27860 34972 27870 35028
rect 30940 34972 43036 35028
rect 43092 34972 44268 35028
rect 44324 34972 44940 35028
rect 44996 34972 45388 35028
rect 45444 34972 45454 35028
rect 45714 34972 45724 35028
rect 45780 34972 45892 35028
rect 46386 34972 46396 35028
rect 46452 34972 47628 35028
rect 47684 34972 47694 35028
rect 47852 34916 47908 35084
rect 51538 34972 51548 35028
rect 51604 34972 54348 35028
rect 54404 34972 54414 35028
rect 15362 34860 15372 34916
rect 15428 34860 16268 34916
rect 16324 34860 16940 34916
rect 16996 34860 18060 34916
rect 18116 34860 21868 34916
rect 21924 34860 21934 34916
rect 28914 34860 28924 34916
rect 28980 34860 29484 34916
rect 29540 34860 30604 34916
rect 30660 34860 30670 34916
rect 34738 34860 34748 34916
rect 34804 34860 35420 34916
rect 35476 34860 35486 34916
rect 36194 34860 36204 34916
rect 36260 34860 37100 34916
rect 37156 34860 38444 34916
rect 38500 34860 38510 34916
rect 40002 34860 40012 34916
rect 40068 34860 41244 34916
rect 41300 34860 41310 34916
rect 43698 34860 43708 34916
rect 43764 34860 45948 34916
rect 46004 34860 46732 34916
rect 46788 34860 46798 34916
rect 47852 34860 53116 34916
rect 53172 34860 53182 34916
rect 53340 34860 57260 34916
rect 57316 34860 57326 34916
rect 60610 34860 60620 34916
rect 60676 34860 60956 34916
rect 61012 34860 61022 34916
rect 53340 34804 53396 34860
rect 22194 34748 22204 34804
rect 22260 34748 24220 34804
rect 24276 34748 24286 34804
rect 24444 34748 27748 34804
rect 28802 34748 28812 34804
rect 28868 34748 29708 34804
rect 29764 34748 30828 34804
rect 30884 34748 30894 34804
rect 40338 34748 40348 34804
rect 40404 34748 41132 34804
rect 41188 34748 41198 34804
rect 42578 34748 42588 34804
rect 42644 34748 43484 34804
rect 43540 34748 44044 34804
rect 44100 34748 45612 34804
rect 45668 34748 45678 34804
rect 45826 34748 45836 34804
rect 45892 34748 53396 34804
rect 53554 34748 53564 34804
rect 53620 34748 55132 34804
rect 55188 34748 55198 34804
rect 57922 34748 57932 34804
rect 57988 34748 60284 34804
rect 60340 34748 60350 34804
rect 24444 34692 24500 34748
rect 27692 34692 27748 34748
rect 15922 34636 15932 34692
rect 15988 34636 17500 34692
rect 17556 34636 17566 34692
rect 24434 34636 24444 34692
rect 24500 34636 24510 34692
rect 26852 34636 27132 34692
rect 27188 34636 27198 34692
rect 27682 34636 27692 34692
rect 27748 34636 28364 34692
rect 28420 34636 44548 34692
rect 45154 34636 45164 34692
rect 45220 34636 49196 34692
rect 49252 34636 50652 34692
rect 50708 34636 50718 34692
rect 50988 34636 70588 34692
rect 20522 34468 20532 34524
rect 20588 34468 20636 34524
rect 20692 34468 20740 34524
rect 20796 34468 20806 34524
rect 26852 34468 26908 34636
rect 44492 34580 44548 34636
rect 50988 34580 51044 34636
rect 70532 34580 70588 34636
rect 27458 34524 27468 34580
rect 27524 34524 29820 34580
rect 29876 34524 29886 34580
rect 30706 34524 30716 34580
rect 30772 34524 31500 34580
rect 31556 34524 31566 34580
rect 44492 34524 51044 34580
rect 51762 34524 51772 34580
rect 51828 34524 58940 34580
rect 58996 34524 59006 34580
rect 70532 34524 76300 34580
rect 76356 34524 76366 34580
rect 39842 34468 39852 34524
rect 39908 34468 39956 34524
rect 40012 34468 40060 34524
rect 40116 34468 40126 34524
rect 51772 34468 51828 34524
rect 59162 34468 59172 34524
rect 59228 34468 59276 34524
rect 59332 34468 59380 34524
rect 59436 34468 59446 34524
rect 78482 34468 78492 34524
rect 78548 34468 78596 34524
rect 78652 34468 78700 34524
rect 78756 34468 78766 34524
rect 14466 34412 14476 34468
rect 14532 34412 15820 34468
rect 15876 34412 15886 34468
rect 23426 34412 23436 34468
rect 23492 34412 26908 34468
rect 30044 34412 35644 34468
rect 35700 34412 36428 34468
rect 36484 34412 36494 34468
rect 48066 34412 48076 34468
rect 48132 34412 49420 34468
rect 49476 34412 51828 34468
rect 53666 34412 53676 34468
rect 53732 34412 58828 34468
rect 58884 34412 58894 34468
rect 70532 34412 70924 34468
rect 70980 34412 70990 34468
rect 30044 34356 30100 34412
rect 3042 34300 3052 34356
rect 3108 34300 23660 34356
rect 23716 34300 24444 34356
rect 24500 34300 24510 34356
rect 28354 34300 28364 34356
rect 28420 34300 30044 34356
rect 30100 34300 30110 34356
rect 31938 34300 31948 34356
rect 32004 34300 33292 34356
rect 33348 34300 33358 34356
rect 36530 34300 36540 34356
rect 36596 34300 36876 34356
rect 36932 34300 36942 34356
rect 41234 34300 41244 34356
rect 41300 34300 41916 34356
rect 41972 34300 41982 34356
rect 44146 34300 44156 34356
rect 44212 34300 45724 34356
rect 45780 34300 45790 34356
rect 54450 34300 54460 34356
rect 54516 34300 55580 34356
rect 55636 34300 55646 34356
rect 62132 34300 63532 34356
rect 63588 34300 63598 34356
rect 17602 34188 17612 34244
rect 17668 34188 18284 34244
rect 18340 34188 28588 34244
rect 28644 34188 28654 34244
rect 29922 34188 29932 34244
rect 29988 34188 43484 34244
rect 43540 34188 43550 34244
rect 44706 34188 44716 34244
rect 44772 34188 45836 34244
rect 45892 34188 45902 34244
rect 60050 34188 60060 34244
rect 60116 34188 60732 34244
rect 60788 34188 60798 34244
rect 62132 34132 62188 34300
rect 70532 34244 70588 34412
rect 66434 34188 66444 34244
rect 66500 34188 67340 34244
rect 67396 34188 67406 34244
rect 70018 34188 70028 34244
rect 70084 34188 70588 34244
rect 10322 34076 10332 34132
rect 10388 34076 11004 34132
rect 11060 34076 13804 34132
rect 13860 34076 13870 34132
rect 16034 34076 16044 34132
rect 16100 34076 17836 34132
rect 17892 34076 17902 34132
rect 20514 34076 20524 34132
rect 20580 34076 21420 34132
rect 21476 34076 21486 34132
rect 22306 34076 22316 34132
rect 22372 34076 22988 34132
rect 23044 34076 25900 34132
rect 25956 34076 26908 34132
rect 31490 34076 31500 34132
rect 31556 34076 32060 34132
rect 32116 34076 34076 34132
rect 34132 34076 34142 34132
rect 36530 34076 36540 34132
rect 36596 34076 39340 34132
rect 39396 34076 39406 34132
rect 49858 34076 49868 34132
rect 49924 34076 58044 34132
rect 58100 34076 62188 34132
rect 64754 34076 64764 34132
rect 64820 34076 65660 34132
rect 65716 34076 65726 34132
rect 69682 34076 69692 34132
rect 69748 34076 70476 34132
rect 70532 34076 70542 34132
rect 70802 34076 70812 34132
rect 70868 34076 73052 34132
rect 73108 34076 73118 34132
rect 75058 34076 75068 34132
rect 75124 34076 77980 34132
rect 78036 34076 78046 34132
rect 4274 33964 4284 34020
rect 4340 33964 4844 34020
rect 4900 33964 18172 34020
rect 18228 33964 18238 34020
rect 18722 33964 18732 34020
rect 18788 33964 19516 34020
rect 19572 33964 24108 34020
rect 24164 33964 25340 34020
rect 25396 33964 25564 34020
rect 25620 33964 25630 34020
rect 26852 33908 26908 34076
rect 28018 33964 28028 34020
rect 28084 33964 31948 34020
rect 32004 33964 32014 34020
rect 32386 33964 32396 34020
rect 32452 33964 33852 34020
rect 33908 33964 37436 34020
rect 37492 33964 37502 34020
rect 39666 33964 39676 34020
rect 39732 33964 41468 34020
rect 41524 33964 42028 34020
rect 42084 33964 42094 34020
rect 51986 33964 51996 34020
rect 52052 33964 54124 34020
rect 54180 33964 55356 34020
rect 55412 33964 55422 34020
rect 58818 33964 58828 34020
rect 58884 33964 63644 34020
rect 63700 33964 63710 34020
rect 69346 33964 69356 34020
rect 69412 33964 71036 34020
rect 71092 33964 71102 34020
rect 26852 33852 38668 33908
rect 41122 33852 41132 33908
rect 41188 33852 53228 33908
rect 53284 33852 53294 33908
rect 38612 33796 38668 33852
rect 32498 33740 32508 33796
rect 32564 33740 34300 33796
rect 34356 33740 34366 33796
rect 38612 33740 42588 33796
rect 42644 33740 42654 33796
rect 10862 33684 10872 33740
rect 10928 33684 10976 33740
rect 11032 33684 11080 33740
rect 11136 33684 11146 33740
rect 30182 33684 30192 33740
rect 30248 33684 30296 33740
rect 30352 33684 30400 33740
rect 30456 33684 30466 33740
rect 49502 33684 49512 33740
rect 49568 33684 49616 33740
rect 49672 33684 49720 33740
rect 49776 33684 49786 33740
rect 68822 33684 68832 33740
rect 68888 33684 68936 33740
rect 68992 33684 69040 33740
rect 69096 33684 69106 33740
rect 33954 33628 33964 33684
rect 34020 33628 34524 33684
rect 34580 33628 34590 33684
rect 11666 33516 11676 33572
rect 11732 33516 12572 33572
rect 12628 33516 12638 33572
rect 19730 33516 19740 33572
rect 19796 33516 38668 33572
rect 47730 33516 47740 33572
rect 47796 33516 48860 33572
rect 48916 33516 48926 33572
rect 58818 33516 58828 33572
rect 58884 33516 59276 33572
rect 59332 33516 59342 33572
rect 60834 33516 60844 33572
rect 60900 33516 61964 33572
rect 62020 33516 62030 33572
rect 65090 33516 65100 33572
rect 65156 33516 66444 33572
rect 66500 33516 66510 33572
rect 0 33460 800 33488
rect 38612 33460 38668 33516
rect 79200 33460 80000 33488
rect 0 33404 1932 33460
rect 1988 33404 1998 33460
rect 11218 33404 11228 33460
rect 11284 33404 13468 33460
rect 13524 33404 13534 33460
rect 20850 33404 20860 33460
rect 20916 33404 21868 33460
rect 21924 33404 21934 33460
rect 23538 33404 23548 33460
rect 23604 33404 24780 33460
rect 24836 33404 26908 33460
rect 28578 33404 28588 33460
rect 28644 33404 31388 33460
rect 31444 33404 31454 33460
rect 31826 33404 31836 33460
rect 31892 33404 33180 33460
rect 33236 33404 33246 33460
rect 33506 33404 33516 33460
rect 33572 33404 36204 33460
rect 36260 33404 37212 33460
rect 37268 33404 37772 33460
rect 37828 33404 37838 33460
rect 38612 33404 43036 33460
rect 43092 33404 43484 33460
rect 43540 33404 44828 33460
rect 44884 33404 44894 33460
rect 45378 33404 45388 33460
rect 45444 33404 57596 33460
rect 57652 33404 57662 33460
rect 72930 33404 72940 33460
rect 72996 33404 73276 33460
rect 73332 33404 73342 33460
rect 77970 33404 77980 33460
rect 78036 33404 80000 33460
rect 0 33376 800 33404
rect 4722 33292 4732 33348
rect 4788 33292 14476 33348
rect 14532 33292 14542 33348
rect 18498 33292 18508 33348
rect 18564 33292 22876 33348
rect 22932 33292 22942 33348
rect 25554 33292 25564 33348
rect 25620 33292 26684 33348
rect 26740 33292 26750 33348
rect 13570 33180 13580 33236
rect 13636 33180 18620 33236
rect 18676 33180 18686 33236
rect 20514 33180 20524 33236
rect 20580 33180 21644 33236
rect 21700 33180 21710 33236
rect 15698 33068 15708 33124
rect 15764 33068 16716 33124
rect 16772 33068 16782 33124
rect 20290 33068 20300 33124
rect 20356 33068 20636 33124
rect 20692 33068 20702 33124
rect 22082 33068 22092 33124
rect 22148 33068 23324 33124
rect 23380 33068 24332 33124
rect 24388 33068 25228 33124
rect 25284 33068 26348 33124
rect 26404 33068 26414 33124
rect 20300 33012 20356 33068
rect 26852 33012 26908 33404
rect 44828 33348 44884 33404
rect 79200 33376 80000 33404
rect 28242 33292 28252 33348
rect 28308 33292 30380 33348
rect 30436 33292 30446 33348
rect 36642 33292 36652 33348
rect 36708 33292 37548 33348
rect 37604 33292 37614 33348
rect 38882 33292 38892 33348
rect 38948 33292 39452 33348
rect 39508 33292 39518 33348
rect 44828 33292 45836 33348
rect 45892 33292 45902 33348
rect 49186 33292 49196 33348
rect 49252 33292 51660 33348
rect 51716 33292 51726 33348
rect 53666 33292 53676 33348
rect 53732 33292 54348 33348
rect 54404 33292 54908 33348
rect 54964 33292 55804 33348
rect 55860 33292 55870 33348
rect 56354 33292 56364 33348
rect 56420 33292 58044 33348
rect 58100 33292 59052 33348
rect 59108 33292 59118 33348
rect 66770 33292 66780 33348
rect 66836 33292 67676 33348
rect 67732 33292 67742 33348
rect 28130 33180 28140 33236
rect 28196 33180 29260 33236
rect 29316 33180 29326 33236
rect 31154 33180 31164 33236
rect 31220 33180 32060 33236
rect 32116 33180 33852 33236
rect 33908 33180 34748 33236
rect 34804 33180 34814 33236
rect 36418 33180 36428 33236
rect 36484 33180 37324 33236
rect 37380 33180 37996 33236
rect 38052 33180 38062 33236
rect 50530 33180 50540 33236
rect 50596 33180 57148 33236
rect 57204 33180 57214 33236
rect 73154 33180 73164 33236
rect 73220 33180 76300 33236
rect 76356 33180 76366 33236
rect 29260 33124 29316 33180
rect 29260 33068 29820 33124
rect 29876 33068 29886 33124
rect 32386 33068 32396 33124
rect 32452 33068 33180 33124
rect 33236 33068 33246 33124
rect 38434 33068 38444 33124
rect 38500 33068 49868 33124
rect 49924 33068 50652 33124
rect 50708 33068 50718 33124
rect 65986 33068 65996 33124
rect 66052 33068 67004 33124
rect 67060 33068 69356 33124
rect 69412 33068 69422 33124
rect 69682 33068 69692 33124
rect 69748 33068 75404 33124
rect 75460 33068 75470 33124
rect 16370 32956 16380 33012
rect 16436 32956 20356 33012
rect 20962 32956 20972 33012
rect 21028 32956 21532 33012
rect 21588 32956 21598 33012
rect 22866 32956 22876 33012
rect 22932 32956 23772 33012
rect 23828 32956 23838 33012
rect 26852 32956 36876 33012
rect 36932 32956 36942 33012
rect 20522 32900 20532 32956
rect 20588 32900 20636 32956
rect 20692 32900 20740 32956
rect 20796 32900 20806 32956
rect 39842 32900 39852 32956
rect 39908 32900 39956 32956
rect 40012 32900 40060 32956
rect 40116 32900 40126 32956
rect 59162 32900 59172 32956
rect 59228 32900 59276 32956
rect 59332 32900 59380 32956
rect 59436 32900 59446 32956
rect 78482 32900 78492 32956
rect 78548 32900 78596 32956
rect 78652 32900 78700 32956
rect 78756 32900 78766 32956
rect 14914 32844 14924 32900
rect 14980 32844 19292 32900
rect 19348 32844 19358 32900
rect 25106 32844 25116 32900
rect 25172 32844 27468 32900
rect 27524 32844 27534 32900
rect 36418 32844 36428 32900
rect 36484 32844 37212 32900
rect 37268 32844 38556 32900
rect 38612 32844 38622 32900
rect 12674 32732 12684 32788
rect 12740 32732 14252 32788
rect 14308 32732 14318 32788
rect 14578 32732 14588 32788
rect 14644 32732 16268 32788
rect 16324 32732 20972 32788
rect 21028 32732 21038 32788
rect 26674 32732 26684 32788
rect 26740 32732 39452 32788
rect 39508 32732 39518 32788
rect 39676 32732 42700 32788
rect 42756 32732 43036 32788
rect 43092 32732 43932 32788
rect 43988 32732 43998 32788
rect 45266 32732 45276 32788
rect 45332 32732 45612 32788
rect 45668 32732 46284 32788
rect 46340 32732 46350 32788
rect 57362 32732 57372 32788
rect 57428 32732 58156 32788
rect 58212 32732 59500 32788
rect 59556 32732 59566 32788
rect 59826 32732 59836 32788
rect 59892 32732 61292 32788
rect 61348 32732 61358 32788
rect 14588 32676 14644 32732
rect 39676 32676 39732 32732
rect 13906 32620 13916 32676
rect 13972 32620 14644 32676
rect 21298 32620 21308 32676
rect 21364 32620 22540 32676
rect 22596 32620 22606 32676
rect 26338 32620 26348 32676
rect 26404 32620 39732 32676
rect 39890 32620 39900 32676
rect 39956 32620 40236 32676
rect 40292 32620 41692 32676
rect 41748 32620 41758 32676
rect 14578 32508 14588 32564
rect 14644 32508 15148 32564
rect 15204 32508 15214 32564
rect 19282 32508 19292 32564
rect 19348 32508 19964 32564
rect 20020 32508 25452 32564
rect 25508 32508 26124 32564
rect 26180 32508 27356 32564
rect 27412 32508 30828 32564
rect 30884 32508 30894 32564
rect 37314 32508 37324 32564
rect 37380 32508 38892 32564
rect 38948 32508 38958 32564
rect 39666 32508 39676 32564
rect 39732 32508 41356 32564
rect 41412 32508 41422 32564
rect 15362 32396 15372 32452
rect 15428 32396 15932 32452
rect 15988 32396 16380 32452
rect 16436 32396 16446 32452
rect 19506 32396 19516 32452
rect 19572 32396 20412 32452
rect 20468 32396 25228 32452
rect 25284 32396 26572 32452
rect 26628 32396 26638 32452
rect 31826 32396 31836 32452
rect 31892 32396 34188 32452
rect 34244 32396 34254 32452
rect 37202 32396 37212 32452
rect 37268 32396 38444 32452
rect 38500 32396 38510 32452
rect 39442 32396 39452 32452
rect 39508 32396 42364 32452
rect 42420 32396 42700 32452
rect 42756 32396 42766 32452
rect 44818 32396 44828 32452
rect 44884 32396 45164 32452
rect 45220 32396 45230 32452
rect 57586 32396 57596 32452
rect 57652 32396 58492 32452
rect 58548 32396 58558 32452
rect 64418 32396 64428 32452
rect 64484 32396 66220 32452
rect 66276 32396 66668 32452
rect 66724 32396 69244 32452
rect 69300 32396 70476 32452
rect 70532 32396 70542 32452
rect 16706 32284 16716 32340
rect 16772 32284 33628 32340
rect 33684 32284 33694 32340
rect 71250 32284 71260 32340
rect 71316 32284 73276 32340
rect 73332 32284 73342 32340
rect 10862 32116 10872 32172
rect 10928 32116 10976 32172
rect 11032 32116 11080 32172
rect 11136 32116 11146 32172
rect 30182 32116 30192 32172
rect 30248 32116 30296 32172
rect 30352 32116 30400 32172
rect 30456 32116 30466 32172
rect 49502 32116 49512 32172
rect 49568 32116 49616 32172
rect 49672 32116 49720 32172
rect 49776 32116 49786 32172
rect 68822 32116 68832 32172
rect 68888 32116 68936 32172
rect 68992 32116 69040 32172
rect 69096 32116 69106 32172
rect 31378 32060 31388 32116
rect 31444 32060 33404 32116
rect 33460 32060 33470 32116
rect 34738 32060 34748 32116
rect 34804 32060 38668 32116
rect 59602 32060 59612 32116
rect 59668 32060 63644 32116
rect 63700 32060 63710 32116
rect 38612 32004 38668 32060
rect 25442 31948 25452 32004
rect 25508 31948 27916 32004
rect 27972 31948 27982 32004
rect 29474 31948 29484 32004
rect 29540 31948 30604 32004
rect 30660 31948 31836 32004
rect 31892 31948 31902 32004
rect 32274 31948 32284 32004
rect 32340 31948 34076 32004
rect 34132 31948 37436 32004
rect 37492 31948 37502 32004
rect 38612 31948 48524 32004
rect 48580 31948 48590 32004
rect 50642 31948 50652 32004
rect 50708 31948 51212 32004
rect 51268 31948 51278 32004
rect 18498 31836 18508 31892
rect 18564 31836 18956 31892
rect 19012 31836 19022 31892
rect 23314 31836 23324 31892
rect 23380 31836 24668 31892
rect 24724 31836 24734 31892
rect 30156 31780 30212 31948
rect 31378 31836 31388 31892
rect 31444 31836 33740 31892
rect 33796 31836 33806 31892
rect 39442 31836 39452 31892
rect 39508 31836 39788 31892
rect 39844 31836 39854 31892
rect 42354 31836 42364 31892
rect 42420 31836 46172 31892
rect 46228 31836 46238 31892
rect 46396 31836 47964 31892
rect 48020 31836 48030 31892
rect 48962 31836 48972 31892
rect 49028 31836 50092 31892
rect 50148 31836 50158 31892
rect 60386 31836 60396 31892
rect 60452 31836 64652 31892
rect 64708 31836 64876 31892
rect 64932 31836 64942 31892
rect 46396 31780 46452 31836
rect 4274 31724 4284 31780
rect 4340 31724 14140 31780
rect 14196 31724 15036 31780
rect 15092 31724 15102 31780
rect 22754 31724 22764 31780
rect 22820 31724 23660 31780
rect 23716 31724 23726 31780
rect 23874 31724 23884 31780
rect 23940 31724 25004 31780
rect 25060 31724 25070 31780
rect 30146 31724 30156 31780
rect 30212 31724 30222 31780
rect 31490 31724 31500 31780
rect 31556 31724 32172 31780
rect 32228 31724 32238 31780
rect 33394 31724 33404 31780
rect 33460 31724 35756 31780
rect 35812 31724 36540 31780
rect 36596 31724 36606 31780
rect 36978 31724 36988 31780
rect 37044 31724 46452 31780
rect 46610 31724 46620 31780
rect 46676 31724 53900 31780
rect 53956 31724 59948 31780
rect 60004 31724 60844 31780
rect 60900 31724 61516 31780
rect 61572 31724 61582 31780
rect 17826 31612 17836 31668
rect 17892 31612 27356 31668
rect 27412 31612 28588 31668
rect 28644 31612 28654 31668
rect 30370 31612 30380 31668
rect 30436 31612 31388 31668
rect 31444 31612 31454 31668
rect 32274 31612 32284 31668
rect 32340 31612 33180 31668
rect 33236 31612 39004 31668
rect 39060 31612 39070 31668
rect 43474 31612 43484 31668
rect 43540 31612 45052 31668
rect 45108 31612 49644 31668
rect 49700 31612 51436 31668
rect 51492 31612 51502 31668
rect 60050 31612 60060 31668
rect 60116 31612 60620 31668
rect 60676 31612 60686 31668
rect 14802 31500 14812 31556
rect 14868 31500 16044 31556
rect 16100 31500 16110 31556
rect 23538 31500 23548 31556
rect 23604 31500 24220 31556
rect 24276 31500 26460 31556
rect 26516 31500 26526 31556
rect 27122 31500 27132 31556
rect 27188 31500 29596 31556
rect 29652 31500 30492 31556
rect 30548 31500 30558 31556
rect 31042 31500 31052 31556
rect 31108 31500 32396 31556
rect 32452 31500 32462 31556
rect 33506 31500 33516 31556
rect 33572 31500 39116 31556
rect 39172 31500 39182 31556
rect 43698 31500 43708 31556
rect 43764 31500 43932 31556
rect 43988 31500 44940 31556
rect 44996 31500 45388 31556
rect 45444 31500 45454 31556
rect 46722 31500 46732 31556
rect 46788 31500 47516 31556
rect 47572 31500 48636 31556
rect 48692 31500 48702 31556
rect 48962 31500 48972 31556
rect 49028 31500 49420 31556
rect 49476 31500 50876 31556
rect 50932 31500 50942 31556
rect 65202 31500 65212 31556
rect 65268 31500 66332 31556
rect 66388 31500 69132 31556
rect 69188 31500 69916 31556
rect 69972 31500 69982 31556
rect 33516 31444 33572 31500
rect 9538 31388 9548 31444
rect 9604 31388 9996 31444
rect 10052 31388 19068 31444
rect 19124 31388 19134 31444
rect 28242 31388 28252 31444
rect 28308 31388 30940 31444
rect 30996 31388 33572 31444
rect 50978 31388 50988 31444
rect 51044 31388 51548 31444
rect 51604 31388 51614 31444
rect 20522 31332 20532 31388
rect 20588 31332 20636 31388
rect 20692 31332 20740 31388
rect 20796 31332 20806 31388
rect 39842 31332 39852 31388
rect 39908 31332 39956 31388
rect 40012 31332 40060 31388
rect 40116 31332 40126 31388
rect 59162 31332 59172 31388
rect 59228 31332 59276 31388
rect 59332 31332 59380 31388
rect 59436 31332 59446 31388
rect 78482 31332 78492 31388
rect 78548 31332 78596 31388
rect 78652 31332 78700 31388
rect 78756 31332 78766 31388
rect 18386 31276 18396 31332
rect 18452 31276 19404 31332
rect 19460 31276 19470 31332
rect 31266 31276 31276 31332
rect 31332 31276 32396 31332
rect 32452 31276 32462 31332
rect 33740 31276 38668 31332
rect 40786 31276 40796 31332
rect 40852 31276 50540 31332
rect 50596 31276 50606 31332
rect 33740 31220 33796 31276
rect 4050 31164 4060 31220
rect 4116 31164 33740 31220
rect 33796 31164 33806 31220
rect 35634 31164 35644 31220
rect 35700 31164 36988 31220
rect 37044 31164 37054 31220
rect 38612 31108 38668 31276
rect 40002 31164 40012 31220
rect 40068 31164 41244 31220
rect 41300 31164 41310 31220
rect 43708 31164 45220 31220
rect 45378 31164 45388 31220
rect 45444 31164 73948 31220
rect 74004 31164 74014 31220
rect 43708 31108 43764 31164
rect 45164 31108 45220 31164
rect 5170 31052 5180 31108
rect 5236 31052 8428 31108
rect 19842 31052 19852 31108
rect 19908 31052 20076 31108
rect 20132 31052 20142 31108
rect 24994 31052 25004 31108
rect 25060 31052 26236 31108
rect 26292 31052 26302 31108
rect 30146 31052 30156 31108
rect 30212 31052 31612 31108
rect 31668 31052 31678 31108
rect 38612 31052 43764 31108
rect 43820 31052 44604 31108
rect 44660 31052 44670 31108
rect 45164 31052 48972 31108
rect 49028 31052 49308 31108
rect 49364 31052 49374 31108
rect 69906 31052 69916 31108
rect 69972 31052 74172 31108
rect 74228 31052 74238 31108
rect 0 30996 800 31024
rect 8372 30996 8428 31052
rect 43820 30996 43876 31052
rect 79200 30996 80000 31024
rect 0 30940 1932 30996
rect 1988 30940 1998 30996
rect 8372 30940 17668 30996
rect 17938 30940 17948 30996
rect 18004 30940 23548 30996
rect 23604 30940 23614 30996
rect 23874 30940 23884 30996
rect 23940 30940 28588 30996
rect 28644 30940 28654 30996
rect 36530 30940 36540 30996
rect 36596 30940 37436 30996
rect 37492 30940 37502 30996
rect 38210 30940 38220 30996
rect 38276 30940 38892 30996
rect 38948 30940 39788 30996
rect 39844 30940 41020 30996
rect 41076 30940 41086 30996
rect 42466 30940 42476 30996
rect 42532 30940 43820 30996
rect 43876 30940 43886 30996
rect 44258 30940 44268 30996
rect 44324 30940 46844 30996
rect 46900 30940 46910 30996
rect 51314 30940 51324 30996
rect 51380 30940 53564 30996
rect 53620 30940 53630 30996
rect 58706 30940 58716 30996
rect 58772 30940 59948 30996
rect 60004 30940 60396 30996
rect 60452 30940 60462 30996
rect 77970 30940 77980 30996
rect 78036 30940 80000 30996
rect 0 30912 800 30940
rect 17612 30884 17668 30940
rect 79200 30912 80000 30940
rect 14914 30828 14924 30884
rect 14980 30828 17052 30884
rect 17108 30828 17118 30884
rect 17612 30828 21308 30884
rect 21364 30828 21374 30884
rect 24658 30828 24668 30884
rect 24724 30828 25564 30884
rect 25620 30828 26012 30884
rect 26068 30828 26078 30884
rect 36642 30828 36652 30884
rect 36708 30828 37212 30884
rect 37268 30828 37996 30884
rect 38052 30828 38062 30884
rect 39116 30828 42252 30884
rect 42308 30828 42318 30884
rect 47954 30828 47964 30884
rect 48020 30828 56700 30884
rect 56756 30828 56766 30884
rect 75282 30828 75292 30884
rect 75348 30828 77756 30884
rect 77812 30828 77822 30884
rect 39116 30772 39172 30828
rect 15092 30716 15260 30772
rect 15316 30716 20076 30772
rect 20132 30716 21420 30772
rect 21476 30716 21486 30772
rect 32610 30716 32620 30772
rect 32676 30716 39172 30772
rect 39228 30716 43148 30772
rect 43204 30716 43214 30772
rect 15092 30660 15148 30716
rect 39228 30660 39284 30716
rect 14466 30604 14476 30660
rect 14532 30604 15148 30660
rect 30706 30604 30716 30660
rect 30772 30604 39284 30660
rect 39442 30604 39452 30660
rect 39508 30604 42252 30660
rect 42308 30604 42318 30660
rect 55458 30604 55468 30660
rect 55524 30604 58604 30660
rect 58660 30604 59724 30660
rect 59780 30604 61068 30660
rect 61124 30604 61134 30660
rect 10862 30548 10872 30604
rect 10928 30548 10976 30604
rect 11032 30548 11080 30604
rect 11136 30548 11146 30604
rect 30182 30548 30192 30604
rect 30248 30548 30296 30604
rect 30352 30548 30400 30604
rect 30456 30548 30466 30604
rect 49502 30548 49512 30604
rect 49568 30548 49616 30604
rect 49672 30548 49720 30604
rect 49776 30548 49786 30604
rect 68822 30548 68832 30604
rect 68888 30548 68936 30604
rect 68992 30548 69040 30604
rect 69096 30548 69106 30604
rect 20178 30492 20188 30548
rect 20244 30492 20748 30548
rect 20804 30492 28140 30548
rect 28196 30492 28206 30548
rect 37874 30492 37884 30548
rect 37940 30492 38668 30548
rect 38612 30436 38668 30492
rect 50372 30492 60284 30548
rect 60340 30492 60350 30548
rect 50372 30436 50428 30492
rect 16482 30380 16492 30436
rect 16548 30380 17388 30436
rect 17444 30380 17454 30436
rect 22418 30380 22428 30436
rect 22484 30380 23324 30436
rect 23380 30380 24108 30436
rect 24164 30380 26684 30436
rect 26740 30380 29652 30436
rect 36082 30380 36092 30436
rect 36148 30380 36652 30436
rect 36708 30380 37660 30436
rect 37716 30380 37726 30436
rect 38612 30380 50428 30436
rect 53778 30380 53788 30436
rect 53844 30380 54908 30436
rect 54964 30380 54974 30436
rect 59490 30380 59500 30436
rect 59556 30380 59836 30436
rect 59892 30380 59902 30436
rect 69122 30380 69132 30436
rect 69188 30380 69916 30436
rect 69972 30380 69982 30436
rect 29596 30324 29652 30380
rect 16146 30268 16156 30324
rect 16212 30268 16222 30324
rect 19058 30268 19068 30324
rect 19124 30268 22652 30324
rect 22708 30268 22718 30324
rect 24882 30268 24892 30324
rect 24948 30268 29428 30324
rect 29586 30268 29596 30324
rect 29652 30268 29662 30324
rect 33506 30268 33516 30324
rect 33572 30268 34524 30324
rect 34580 30268 34590 30324
rect 35308 30268 41804 30324
rect 41860 30268 42476 30324
rect 42532 30268 42542 30324
rect 56690 30268 56700 30324
rect 56756 30268 58156 30324
rect 58212 30268 58716 30324
rect 58772 30268 58782 30324
rect 68562 30268 68572 30324
rect 68628 30268 76636 30324
rect 76692 30268 77308 30324
rect 77364 30268 77980 30324
rect 78036 30268 78046 30324
rect 16156 30212 16212 30268
rect 29372 30212 29428 30268
rect 13122 30156 13132 30212
rect 13188 30156 14700 30212
rect 14756 30156 15596 30212
rect 15652 30156 15662 30212
rect 16156 30156 17276 30212
rect 17332 30156 18116 30212
rect 19282 30156 19292 30212
rect 19348 30156 19516 30212
rect 19572 30156 20188 30212
rect 20244 30156 22876 30212
rect 22932 30156 22942 30212
rect 23986 30156 23996 30212
rect 24052 30156 25452 30212
rect 25508 30156 25518 30212
rect 26002 30156 26012 30212
rect 26068 30156 27692 30212
rect 27748 30156 28252 30212
rect 28308 30156 29148 30212
rect 29204 30156 29214 30212
rect 29362 30156 29372 30212
rect 29428 30156 29438 30212
rect 29922 30156 29932 30212
rect 29988 30156 31724 30212
rect 31780 30156 31790 30212
rect 18060 30100 18116 30156
rect 3714 30044 3724 30100
rect 3780 30044 5740 30100
rect 5796 30044 5806 30100
rect 13794 30044 13804 30100
rect 13860 30044 14364 30100
rect 14420 30044 15036 30100
rect 15092 30044 15484 30100
rect 15540 30044 15550 30100
rect 16370 30044 16380 30100
rect 16436 30044 17612 30100
rect 17668 30044 17678 30100
rect 18060 30044 19180 30100
rect 19236 30044 20300 30100
rect 20356 30044 20366 30100
rect 20514 30044 20524 30100
rect 20580 30044 21196 30100
rect 21252 30044 21262 30100
rect 26786 30044 26796 30100
rect 26852 30044 29708 30100
rect 29764 30044 29774 30100
rect 34066 30044 34076 30100
rect 34132 30044 35084 30100
rect 35140 30044 35150 30100
rect 20524 29988 20580 30044
rect 15922 29932 15932 29988
rect 15988 29932 16716 29988
rect 16772 29932 16782 29988
rect 19058 29932 19068 29988
rect 19124 29932 19628 29988
rect 19684 29932 20580 29988
rect 21970 29932 21980 29988
rect 22036 29932 22540 29988
rect 22596 29932 22606 29988
rect 28354 29932 28364 29988
rect 28420 29932 29260 29988
rect 29316 29932 34860 29988
rect 34916 29932 34926 29988
rect 35308 29876 35364 30268
rect 36418 30156 36428 30212
rect 36484 30156 37436 30212
rect 37492 30156 37502 30212
rect 37650 30156 37660 30212
rect 37716 30156 37996 30212
rect 38052 30156 38062 30212
rect 38612 30156 39452 30212
rect 39508 30156 39518 30212
rect 41570 30156 41580 30212
rect 41636 30156 42588 30212
rect 42644 30156 43876 30212
rect 48066 30156 48076 30212
rect 48132 30156 48748 30212
rect 48804 30156 48972 30212
rect 49028 30156 49038 30212
rect 57362 30156 57372 30212
rect 57428 30156 58940 30212
rect 58996 30156 59006 30212
rect 59490 30156 59500 30212
rect 59556 30156 60508 30212
rect 60564 30156 60574 30212
rect 60946 30156 60956 30212
rect 61012 30156 62636 30212
rect 62692 30156 62702 30212
rect 66658 30156 66668 30212
rect 66724 30156 67564 30212
rect 67620 30156 67630 30212
rect 71362 30156 71372 30212
rect 71428 30156 73724 30212
rect 73780 30156 73790 30212
rect 74498 30156 74508 30212
rect 74564 30156 75628 30212
rect 75684 30156 75694 30212
rect 37314 30044 37324 30100
rect 37380 30044 37772 30100
rect 37828 30044 37838 30100
rect 38612 29988 38668 30156
rect 43820 30100 43876 30156
rect 43138 30044 43148 30100
rect 43204 30044 43596 30100
rect 43652 30044 43662 30100
rect 43810 30044 43820 30100
rect 43876 30044 43886 30100
rect 58818 30044 58828 30100
rect 58884 30044 59724 30100
rect 59780 30044 59790 30100
rect 60162 30044 60172 30100
rect 60228 30044 61740 30100
rect 61796 30044 61806 30100
rect 75394 30044 75404 30100
rect 75460 30044 76300 30100
rect 76356 30044 76366 30100
rect 38098 29932 38108 29988
rect 38164 29932 38668 29988
rect 39330 29932 39340 29988
rect 39396 29932 40236 29988
rect 40292 29932 40302 29988
rect 44034 29932 44044 29988
rect 44100 29932 46060 29988
rect 46116 29932 46126 29988
rect 46946 29932 46956 29988
rect 47012 29932 47740 29988
rect 47796 29932 47806 29988
rect 52210 29932 52220 29988
rect 52276 29932 52892 29988
rect 52948 29932 52958 29988
rect 60386 29932 60396 29988
rect 60452 29932 61404 29988
rect 61460 29932 61470 29988
rect 66546 29932 66556 29988
rect 66612 29932 67564 29988
rect 67620 29932 71484 29988
rect 71540 29932 71550 29988
rect 75506 29932 75516 29988
rect 75572 29932 76972 29988
rect 77028 29932 77038 29988
rect 22418 29820 22428 29876
rect 22484 29820 23660 29876
rect 23716 29820 25116 29876
rect 25172 29820 25182 29876
rect 26852 29820 35364 29876
rect 43250 29820 43260 29876
rect 43316 29820 43820 29876
rect 43876 29820 43886 29876
rect 44930 29820 44940 29876
rect 44996 29820 45724 29876
rect 45780 29820 45790 29876
rect 52770 29820 52780 29876
rect 52836 29820 53452 29876
rect 53508 29820 53518 29876
rect 60274 29820 60284 29876
rect 60340 29820 61180 29876
rect 61236 29820 61246 29876
rect 67218 29820 67228 29876
rect 67284 29820 68348 29876
rect 68404 29820 68414 29876
rect 20522 29764 20532 29820
rect 20588 29764 20636 29820
rect 20692 29764 20740 29820
rect 20796 29764 20806 29820
rect 26852 29764 26908 29820
rect 39842 29764 39852 29820
rect 39908 29764 39956 29820
rect 40012 29764 40060 29820
rect 40116 29764 40126 29820
rect 59162 29764 59172 29820
rect 59228 29764 59276 29820
rect 59332 29764 59380 29820
rect 59436 29764 59446 29820
rect 78482 29764 78492 29820
rect 78548 29764 78596 29820
rect 78652 29764 78700 29820
rect 78756 29764 78766 29820
rect 21634 29708 21644 29764
rect 21700 29708 26908 29764
rect 29932 29708 30828 29764
rect 30884 29708 30894 29764
rect 34178 29708 34188 29764
rect 34244 29708 38668 29764
rect 41906 29708 41916 29764
rect 41972 29708 57148 29764
rect 57204 29708 57820 29764
rect 57876 29708 57886 29764
rect 29932 29652 29988 29708
rect 38612 29652 38668 29708
rect 15474 29596 15484 29652
rect 15540 29596 16268 29652
rect 16324 29596 16334 29652
rect 17490 29596 17500 29652
rect 17556 29596 18620 29652
rect 18676 29596 18686 29652
rect 20290 29596 20300 29652
rect 20356 29596 20748 29652
rect 20804 29596 21756 29652
rect 21812 29596 21822 29652
rect 23426 29596 23436 29652
rect 23492 29596 28308 29652
rect 29362 29596 29372 29652
rect 29428 29596 29932 29652
rect 29988 29596 29998 29652
rect 30146 29596 30156 29652
rect 30212 29596 31052 29652
rect 31108 29596 31118 29652
rect 32834 29596 32844 29652
rect 32900 29596 34580 29652
rect 35858 29596 35868 29652
rect 35924 29596 38276 29652
rect 38612 29596 39844 29652
rect 40002 29596 40012 29652
rect 40068 29596 41468 29652
rect 41524 29596 41534 29652
rect 46172 29596 48412 29652
rect 48468 29596 49084 29652
rect 49140 29596 49150 29652
rect 49858 29596 49868 29652
rect 49924 29596 50428 29652
rect 50484 29596 50494 29652
rect 51762 29596 51772 29652
rect 51828 29596 53116 29652
rect 53172 29596 54684 29652
rect 54740 29596 54750 29652
rect 64978 29596 64988 29652
rect 65044 29596 65772 29652
rect 65828 29596 65838 29652
rect 28252 29540 28308 29596
rect 4946 29484 4956 29540
rect 5012 29484 6748 29540
rect 6804 29484 6814 29540
rect 20626 29484 20636 29540
rect 20692 29484 22092 29540
rect 22148 29484 22158 29540
rect 26114 29484 26124 29540
rect 26180 29484 26796 29540
rect 26852 29484 26862 29540
rect 28252 29484 29708 29540
rect 29764 29484 29774 29540
rect 30034 29484 30044 29540
rect 30100 29484 33180 29540
rect 33236 29484 33246 29540
rect 34524 29428 34580 29596
rect 35522 29484 35532 29540
rect 35588 29484 36988 29540
rect 37044 29484 37054 29540
rect 2482 29372 2492 29428
rect 2548 29372 8540 29428
rect 8596 29372 8606 29428
rect 9986 29372 9996 29428
rect 10052 29372 11340 29428
rect 11396 29372 11406 29428
rect 16706 29372 16716 29428
rect 16772 29372 26460 29428
rect 26516 29372 26526 29428
rect 27122 29372 27132 29428
rect 27188 29372 28644 29428
rect 31490 29372 31500 29428
rect 31556 29372 32172 29428
rect 32228 29372 33292 29428
rect 33348 29372 33358 29428
rect 34524 29372 36204 29428
rect 36260 29372 36270 29428
rect 28588 29316 28644 29372
rect 38220 29316 38276 29596
rect 39788 29540 39844 29596
rect 46172 29540 46228 29596
rect 38434 29484 38444 29540
rect 38500 29484 39004 29540
rect 39060 29484 39070 29540
rect 39788 29484 45108 29540
rect 45266 29484 45276 29540
rect 45332 29484 46172 29540
rect 46228 29484 46238 29540
rect 47170 29484 47180 29540
rect 47236 29484 47740 29540
rect 47796 29484 47806 29540
rect 48290 29484 48300 29540
rect 48356 29484 49756 29540
rect 49812 29484 49822 29540
rect 59266 29484 59276 29540
rect 59332 29484 60844 29540
rect 60900 29484 60910 29540
rect 61180 29484 62748 29540
rect 62804 29484 62814 29540
rect 71026 29484 71036 29540
rect 71092 29484 72268 29540
rect 72324 29484 72716 29540
rect 72772 29484 72782 29540
rect 45052 29428 45108 29484
rect 61180 29428 61236 29484
rect 38658 29372 38668 29428
rect 38724 29372 39340 29428
rect 39396 29372 39788 29428
rect 39844 29372 40348 29428
rect 40404 29372 40414 29428
rect 42578 29372 42588 29428
rect 42644 29372 43932 29428
rect 43988 29372 44716 29428
rect 44772 29372 44782 29428
rect 45052 29372 46732 29428
rect 46788 29372 46798 29428
rect 47842 29372 47852 29428
rect 47908 29372 48636 29428
rect 48692 29372 48702 29428
rect 54786 29372 54796 29428
rect 54852 29372 55580 29428
rect 55636 29372 55646 29428
rect 58146 29372 58156 29428
rect 58212 29372 59948 29428
rect 60004 29372 60014 29428
rect 61170 29372 61180 29428
rect 61236 29372 61246 29428
rect 62066 29372 62076 29428
rect 62132 29372 62412 29428
rect 62468 29372 62478 29428
rect 62636 29372 72772 29428
rect 6514 29260 6524 29316
rect 6580 29260 7420 29316
rect 7476 29260 10220 29316
rect 10276 29260 11788 29316
rect 11844 29260 11854 29316
rect 16594 29260 16604 29316
rect 16660 29260 17836 29316
rect 17892 29260 17902 29316
rect 18274 29260 18284 29316
rect 18340 29260 19740 29316
rect 19796 29260 24220 29316
rect 24276 29260 25228 29316
rect 25284 29260 26684 29316
rect 26740 29260 26750 29316
rect 28018 29260 28028 29316
rect 28084 29260 28094 29316
rect 28578 29260 28588 29316
rect 28644 29260 33404 29316
rect 33460 29260 33470 29316
rect 34290 29260 34300 29316
rect 34356 29260 34860 29316
rect 34916 29260 34926 29316
rect 35746 29260 35756 29316
rect 35812 29260 36988 29316
rect 37044 29260 37054 29316
rect 38220 29260 38444 29316
rect 38500 29260 38510 29316
rect 44258 29260 44268 29316
rect 44324 29260 45948 29316
rect 46004 29260 46956 29316
rect 47012 29260 47022 29316
rect 5282 29148 5292 29204
rect 5348 29148 6076 29204
rect 6132 29148 6748 29204
rect 6804 29148 6814 29204
rect 13234 29148 13244 29204
rect 13300 29148 15708 29204
rect 15764 29148 15774 29204
rect 20514 29148 20524 29204
rect 20580 29148 21532 29204
rect 21588 29148 21598 29204
rect 16146 29036 16156 29092
rect 16212 29036 17500 29092
rect 17556 29036 19292 29092
rect 19348 29036 22428 29092
rect 22484 29036 22494 29092
rect 10862 28980 10872 29036
rect 10928 28980 10976 29036
rect 11032 28980 11080 29036
rect 11136 28980 11146 29036
rect 23492 28980 23548 29260
rect 28028 29204 28084 29260
rect 33404 29204 33460 29260
rect 28028 29148 33348 29204
rect 33404 29148 44940 29204
rect 44996 29148 45006 29204
rect 49746 29148 49756 29204
rect 49812 29148 51436 29204
rect 51492 29148 54124 29204
rect 54180 29148 54190 29204
rect 57474 29148 57484 29204
rect 57540 29148 59612 29204
rect 59668 29148 59678 29204
rect 33292 29092 33348 29148
rect 62636 29092 62692 29372
rect 72716 29316 72772 29372
rect 66882 29260 66892 29316
rect 66948 29260 67900 29316
rect 67956 29260 67966 29316
rect 69682 29260 69692 29316
rect 69748 29260 70700 29316
rect 70756 29260 70766 29316
rect 72706 29260 72716 29316
rect 72772 29260 72782 29316
rect 73826 29260 73836 29316
rect 73892 29260 74732 29316
rect 74788 29260 74798 29316
rect 67900 29204 67956 29260
rect 65202 29148 65212 29204
rect 65268 29148 66556 29204
rect 66612 29148 66622 29204
rect 67900 29148 72828 29204
rect 72884 29148 72894 29204
rect 32386 29036 32396 29092
rect 32452 29036 33068 29092
rect 33124 29036 33134 29092
rect 33292 29036 41804 29092
rect 41860 29036 41870 29092
rect 50372 29036 52052 29092
rect 54450 29036 54460 29092
rect 54516 29036 62692 29092
rect 70466 29036 70476 29092
rect 70532 29036 72044 29092
rect 72100 29036 72110 29092
rect 73938 29036 73948 29092
rect 74004 29036 76524 29092
rect 76580 29036 76590 29092
rect 30182 28980 30192 29036
rect 30248 28980 30296 29036
rect 30352 28980 30400 29036
rect 30456 28980 30466 29036
rect 49502 28980 49512 29036
rect 49568 28980 49616 29036
rect 49672 28980 49720 29036
rect 49776 28980 49786 29036
rect 15092 28924 16828 28980
rect 16884 28924 20748 28980
rect 20804 28924 21644 28980
rect 21700 28924 21710 28980
rect 22866 28924 22876 28980
rect 22932 28924 23548 28980
rect 37090 28924 37100 28980
rect 37156 28924 46956 28980
rect 47012 28924 47022 28980
rect 15092 28756 15148 28924
rect 50372 28868 50428 29036
rect 51996 28980 52052 29036
rect 68822 28980 68832 29036
rect 68888 28980 68936 29036
rect 68992 28980 69040 29036
rect 69096 28980 69106 29036
rect 51762 28924 51772 28980
rect 51828 28924 51838 28980
rect 51996 28924 57148 28980
rect 57204 28924 57214 28980
rect 59602 28924 59612 28980
rect 59668 28924 60172 28980
rect 60228 28924 60238 28980
rect 20962 28812 20972 28868
rect 21028 28812 23100 28868
rect 23156 28812 23166 28868
rect 30370 28812 30380 28868
rect 30436 28812 31500 28868
rect 31556 28812 35196 28868
rect 35252 28812 35262 28868
rect 35410 28812 35420 28868
rect 35476 28812 36092 28868
rect 36148 28812 36158 28868
rect 40114 28812 40124 28868
rect 40180 28812 40684 28868
rect 40740 28812 41692 28868
rect 41748 28812 42364 28868
rect 42420 28812 50428 28868
rect 51772 28756 51828 28924
rect 2258 28700 2268 28756
rect 2324 28700 7084 28756
rect 7140 28700 10668 28756
rect 10724 28700 10734 28756
rect 14690 28700 14700 28756
rect 14756 28700 14924 28756
rect 14980 28700 15148 28756
rect 21074 28700 21084 28756
rect 21140 28700 23212 28756
rect 23268 28700 24892 28756
rect 24948 28700 26236 28756
rect 26292 28700 26302 28756
rect 32050 28700 32060 28756
rect 32116 28700 33180 28756
rect 33236 28700 33246 28756
rect 38994 28700 39004 28756
rect 39060 28700 39788 28756
rect 39844 28700 41580 28756
rect 41636 28700 41646 28756
rect 44930 28700 44940 28756
rect 44996 28700 46844 28756
rect 46900 28700 47292 28756
rect 47348 28700 48860 28756
rect 48916 28700 48926 28756
rect 49970 28700 49980 28756
rect 50036 28700 51828 28756
rect 51884 28812 59052 28868
rect 59108 28812 59118 28868
rect 59938 28812 59948 28868
rect 60004 28812 60956 28868
rect 61012 28812 61022 28868
rect 51884 28644 51940 28812
rect 58482 28700 58492 28756
rect 58548 28700 59332 28756
rect 59276 28644 59332 28700
rect 2930 28588 2940 28644
rect 2996 28588 5628 28644
rect 5684 28588 5694 28644
rect 11330 28588 11340 28644
rect 11396 28588 20860 28644
rect 20916 28588 20926 28644
rect 22082 28588 22092 28644
rect 22148 28588 22540 28644
rect 22596 28588 22606 28644
rect 22754 28588 22764 28644
rect 22820 28588 23884 28644
rect 23940 28588 23950 28644
rect 31602 28588 31612 28644
rect 31668 28588 32396 28644
rect 32452 28588 32462 28644
rect 33282 28588 33292 28644
rect 33348 28588 35308 28644
rect 35364 28588 35374 28644
rect 36642 28588 36652 28644
rect 36708 28588 38220 28644
rect 38276 28588 38668 28644
rect 38724 28588 38734 28644
rect 39106 28588 39116 28644
rect 39172 28588 39564 28644
rect 39620 28588 39630 28644
rect 40450 28588 40460 28644
rect 40516 28588 41020 28644
rect 41076 28588 41086 28644
rect 46386 28588 46396 28644
rect 46452 28588 47852 28644
rect 47908 28588 51940 28644
rect 51996 28588 52780 28644
rect 52836 28588 52846 28644
rect 57922 28588 57932 28644
rect 57988 28588 58716 28644
rect 58772 28588 58782 28644
rect 59266 28588 59276 28644
rect 59332 28588 59612 28644
rect 59668 28588 59678 28644
rect 61394 28588 61404 28644
rect 61460 28588 62076 28644
rect 62132 28588 62142 28644
rect 65874 28588 65884 28644
rect 65940 28588 67116 28644
rect 67172 28588 69692 28644
rect 69748 28588 69758 28644
rect 71922 28588 71932 28644
rect 71988 28588 72492 28644
rect 72548 28588 73836 28644
rect 73892 28588 73902 28644
rect 0 28532 800 28560
rect 51996 28532 52052 28588
rect 79200 28532 80000 28560
rect 0 28476 1932 28532
rect 1988 28476 1998 28532
rect 22642 28476 22652 28532
rect 22708 28476 24836 28532
rect 26450 28476 26460 28532
rect 26516 28476 27580 28532
rect 27636 28476 27646 28532
rect 30930 28476 30940 28532
rect 30996 28476 31006 28532
rect 33730 28476 33740 28532
rect 33796 28476 35644 28532
rect 35700 28476 35710 28532
rect 48514 28476 48524 28532
rect 48580 28476 48972 28532
rect 49028 28476 49038 28532
rect 50306 28476 50316 28532
rect 50372 28476 52052 28532
rect 52108 28476 53788 28532
rect 53844 28476 54572 28532
rect 54628 28476 54638 28532
rect 54898 28476 54908 28532
rect 54964 28476 55916 28532
rect 55972 28476 55982 28532
rect 58258 28476 58268 28532
rect 58324 28476 59052 28532
rect 59108 28476 59118 28532
rect 61282 28476 61292 28532
rect 61348 28476 62972 28532
rect 63028 28476 63038 28532
rect 75394 28476 75404 28532
rect 75460 28476 80000 28532
rect 0 28448 800 28476
rect 24780 28420 24836 28476
rect 30940 28420 30996 28476
rect 52108 28420 52164 28476
rect 79200 28448 80000 28476
rect 15586 28364 15596 28420
rect 15652 28364 17164 28420
rect 17220 28364 18396 28420
rect 18452 28364 18462 28420
rect 23090 28364 23100 28420
rect 23156 28364 23772 28420
rect 23828 28364 24556 28420
rect 24612 28364 24622 28420
rect 24780 28364 30996 28420
rect 33618 28364 33628 28420
rect 33684 28364 34748 28420
rect 34804 28364 36092 28420
rect 36148 28364 36158 28420
rect 36418 28364 36428 28420
rect 36484 28364 37324 28420
rect 37380 28364 38780 28420
rect 38836 28364 39900 28420
rect 39956 28364 39966 28420
rect 43474 28364 43484 28420
rect 43540 28364 51436 28420
rect 51492 28364 52108 28420
rect 52164 28364 52174 28420
rect 52882 28364 52892 28420
rect 52948 28364 53564 28420
rect 53620 28364 53630 28420
rect 57586 28364 57596 28420
rect 57652 28364 58940 28420
rect 58996 28364 59006 28420
rect 59378 28364 59388 28420
rect 59444 28364 60284 28420
rect 60340 28364 60350 28420
rect 60498 28364 60508 28420
rect 60564 28364 61628 28420
rect 61684 28364 62524 28420
rect 62580 28364 62590 28420
rect 22306 28252 22316 28308
rect 22372 28252 22876 28308
rect 22932 28252 22942 28308
rect 26562 28252 26572 28308
rect 26628 28252 26908 28308
rect 26964 28252 26974 28308
rect 27458 28252 27468 28308
rect 27524 28252 31164 28308
rect 31220 28252 31230 28308
rect 34402 28252 34412 28308
rect 34468 28252 35084 28308
rect 35140 28252 35150 28308
rect 52210 28252 52220 28308
rect 52276 28252 52668 28308
rect 52724 28252 52734 28308
rect 52994 28252 53004 28308
rect 53060 28252 53676 28308
rect 53732 28252 53742 28308
rect 60834 28252 60844 28308
rect 60900 28252 61516 28308
rect 61572 28252 62076 28308
rect 62132 28252 62636 28308
rect 62692 28252 62702 28308
rect 20522 28196 20532 28252
rect 20588 28196 20636 28252
rect 20692 28196 20740 28252
rect 20796 28196 20806 28252
rect 39842 28196 39852 28252
rect 39908 28196 39956 28252
rect 40012 28196 40060 28252
rect 40116 28196 40126 28252
rect 59162 28196 59172 28252
rect 59228 28196 59276 28252
rect 59332 28196 59380 28252
rect 59436 28196 59446 28252
rect 78482 28196 78492 28252
rect 78548 28196 78596 28252
rect 78652 28196 78700 28252
rect 78756 28196 78766 28252
rect 25218 28140 25228 28196
rect 25284 28140 28364 28196
rect 28420 28140 37548 28196
rect 37604 28140 37614 28196
rect 38098 28140 38108 28196
rect 38164 28140 38892 28196
rect 38948 28140 38958 28196
rect 43250 28140 43260 28196
rect 43316 28140 50428 28196
rect 52882 28140 52892 28196
rect 52948 28140 53340 28196
rect 53396 28140 53406 28196
rect 67172 28140 73724 28196
rect 73780 28140 75180 28196
rect 75236 28140 75246 28196
rect 50372 28084 50428 28140
rect 67172 28084 67228 28140
rect 8306 28028 8316 28084
rect 8372 28028 9660 28084
rect 9716 28028 9726 28084
rect 14242 28028 14252 28084
rect 14308 28028 14924 28084
rect 14980 28028 19292 28084
rect 19348 28028 19358 28084
rect 20738 28028 20748 28084
rect 20804 28028 21308 28084
rect 21364 28028 21374 28084
rect 24546 28028 24556 28084
rect 24612 28028 25564 28084
rect 25620 28028 25630 28084
rect 26338 28028 26348 28084
rect 26404 28028 27132 28084
rect 27188 28028 27804 28084
rect 27860 28028 27870 28084
rect 28018 28028 28028 28084
rect 28084 28028 28700 28084
rect 28756 28028 28924 28084
rect 28980 28028 35140 28084
rect 35410 28028 35420 28084
rect 35476 28028 36764 28084
rect 36820 28028 36830 28084
rect 39218 28028 39228 28084
rect 39284 28028 39900 28084
rect 39956 28028 39966 28084
rect 43922 28028 43932 28084
rect 43988 28028 44380 28084
rect 44436 28028 44446 28084
rect 46946 28028 46956 28084
rect 47012 28028 49756 28084
rect 49812 28028 49980 28084
rect 50036 28028 50046 28084
rect 50372 28028 67228 28084
rect 35084 27972 35140 28028
rect 4274 27916 4284 27972
rect 4340 27916 15148 27972
rect 18722 27916 18732 27972
rect 18788 27916 20076 27972
rect 20132 27916 20142 27972
rect 21084 27916 21868 27972
rect 21924 27916 22876 27972
rect 22932 27916 24332 27972
rect 24388 27916 24398 27972
rect 30706 27916 30716 27972
rect 30772 27916 31836 27972
rect 31892 27916 32172 27972
rect 32228 27916 34860 27972
rect 34916 27916 34926 27972
rect 35084 27916 37100 27972
rect 37156 27916 37166 27972
rect 38658 27916 38668 27972
rect 38724 27916 39564 27972
rect 39620 27916 39630 27972
rect 46162 27916 46172 27972
rect 46228 27916 47404 27972
rect 47460 27916 50876 27972
rect 50932 27916 57036 27972
rect 57092 27916 57484 27972
rect 57540 27916 57550 27972
rect 69468 27916 71372 27972
rect 71428 27916 71438 27972
rect 5282 27804 5292 27860
rect 5348 27804 6580 27860
rect 6738 27804 6748 27860
rect 6804 27804 13804 27860
rect 13860 27804 13870 27860
rect 6524 27748 6580 27804
rect 6524 27692 6860 27748
rect 6916 27692 10220 27748
rect 10276 27692 11004 27748
rect 11060 27692 11070 27748
rect 9986 27580 9996 27636
rect 10052 27580 12124 27636
rect 12180 27580 12190 27636
rect 10862 27412 10872 27468
rect 10928 27412 10976 27468
rect 11032 27412 11080 27468
rect 11136 27412 11146 27468
rect 15092 27300 15148 27916
rect 21084 27860 21140 27916
rect 69468 27860 69524 27916
rect 16818 27804 16828 27860
rect 16884 27804 17836 27860
rect 17892 27804 19068 27860
rect 19124 27804 19134 27860
rect 21074 27804 21084 27860
rect 21140 27804 21150 27860
rect 28130 27804 28140 27860
rect 28196 27804 29036 27860
rect 29092 27804 29102 27860
rect 30482 27804 30492 27860
rect 30548 27804 31724 27860
rect 31780 27804 31790 27860
rect 33842 27804 33852 27860
rect 33908 27804 34972 27860
rect 35028 27804 35038 27860
rect 37426 27804 37436 27860
rect 37492 27804 38780 27860
rect 38836 27804 38846 27860
rect 41458 27804 41468 27860
rect 41524 27804 42476 27860
rect 42532 27804 42542 27860
rect 55010 27804 55020 27860
rect 55076 27804 55692 27860
rect 55748 27804 55758 27860
rect 56242 27804 56252 27860
rect 56308 27804 61180 27860
rect 61236 27804 61246 27860
rect 68562 27804 68572 27860
rect 68628 27804 69468 27860
rect 69524 27804 69534 27860
rect 70354 27804 70364 27860
rect 70420 27804 71260 27860
rect 71316 27804 71326 27860
rect 71586 27804 71596 27860
rect 71652 27804 72828 27860
rect 72884 27804 75292 27860
rect 75348 27804 75358 27860
rect 15586 27692 15596 27748
rect 15652 27692 16268 27748
rect 16324 27692 20524 27748
rect 20580 27692 20590 27748
rect 23986 27692 23996 27748
rect 24052 27692 25900 27748
rect 25956 27692 26796 27748
rect 26852 27692 27020 27748
rect 27076 27692 27086 27748
rect 34178 27692 34188 27748
rect 34244 27692 35420 27748
rect 35476 27692 35486 27748
rect 37986 27692 37996 27748
rect 38052 27692 39340 27748
rect 39396 27692 40684 27748
rect 40740 27692 40750 27748
rect 44482 27692 44492 27748
rect 44548 27692 45388 27748
rect 45444 27692 45454 27748
rect 50978 27692 50988 27748
rect 51044 27692 51884 27748
rect 51940 27692 53116 27748
rect 53172 27692 55244 27748
rect 55300 27692 55310 27748
rect 66994 27692 67004 27748
rect 67060 27692 68796 27748
rect 68852 27692 68862 27748
rect 69010 27692 69020 27748
rect 69076 27692 70252 27748
rect 70308 27692 70318 27748
rect 71138 27692 71148 27748
rect 71204 27692 73500 27748
rect 73556 27692 75180 27748
rect 75236 27692 75246 27748
rect 34524 27636 34580 27692
rect 16482 27580 16492 27636
rect 16548 27580 17612 27636
rect 17668 27580 18284 27636
rect 18340 27580 18350 27636
rect 19282 27580 19292 27636
rect 19348 27580 21532 27636
rect 21588 27580 21598 27636
rect 27122 27580 27132 27636
rect 27188 27580 30492 27636
rect 30548 27580 30558 27636
rect 30818 27580 30828 27636
rect 30884 27580 32172 27636
rect 32228 27580 32238 27636
rect 34514 27580 34524 27636
rect 34580 27580 34590 27636
rect 38546 27580 38556 27636
rect 38612 27580 40124 27636
rect 40180 27580 40190 27636
rect 46274 27580 46284 27636
rect 46340 27580 46956 27636
rect 47012 27580 47022 27636
rect 63522 27580 63532 27636
rect 63588 27580 70028 27636
rect 70084 27580 70094 27636
rect 18610 27468 18620 27524
rect 18676 27468 19628 27524
rect 19684 27468 24444 27524
rect 24500 27468 25900 27524
rect 25956 27468 25966 27524
rect 37426 27468 37436 27524
rect 37492 27468 39004 27524
rect 39060 27468 39070 27524
rect 39330 27468 39340 27524
rect 39396 27468 39676 27524
rect 39732 27468 39742 27524
rect 30182 27412 30192 27468
rect 30248 27412 30296 27468
rect 30352 27412 30400 27468
rect 30456 27412 30466 27468
rect 49502 27412 49512 27468
rect 49568 27412 49616 27468
rect 49672 27412 49720 27468
rect 49776 27412 49786 27468
rect 68822 27412 68832 27468
rect 68888 27412 68936 27468
rect 68992 27412 69040 27468
rect 69096 27412 69106 27468
rect 18162 27356 18172 27412
rect 18228 27356 20188 27412
rect 20244 27356 26684 27412
rect 26740 27356 26750 27412
rect 35858 27356 35868 27412
rect 35924 27356 37100 27412
rect 37156 27356 38332 27412
rect 38388 27356 39116 27412
rect 39172 27356 40796 27412
rect 40852 27356 41636 27412
rect 44482 27356 44492 27412
rect 44548 27356 45164 27412
rect 45220 27356 45230 27412
rect 52546 27356 52556 27412
rect 52612 27356 53564 27412
rect 53620 27356 53630 27412
rect 59042 27356 59052 27412
rect 59108 27356 61404 27412
rect 61460 27356 61470 27412
rect 41580 27300 41636 27356
rect 15092 27244 25004 27300
rect 25060 27244 26572 27300
rect 26628 27244 26638 27300
rect 31154 27244 31164 27300
rect 31220 27244 35364 27300
rect 35746 27244 35756 27300
rect 35812 27244 41356 27300
rect 41412 27244 41422 27300
rect 41580 27244 62300 27300
rect 62356 27244 62366 27300
rect 63410 27244 63420 27300
rect 63476 27244 66220 27300
rect 66276 27244 66286 27300
rect 35308 27188 35364 27244
rect 20514 27132 20524 27188
rect 20580 27132 24612 27188
rect 25106 27132 25116 27188
rect 25172 27132 25788 27188
rect 25844 27132 25854 27188
rect 26786 27132 26796 27188
rect 26852 27132 27356 27188
rect 27412 27132 35084 27188
rect 35140 27132 35150 27188
rect 35308 27132 60172 27188
rect 60228 27132 60620 27188
rect 60676 27132 60686 27188
rect 62402 27132 62412 27188
rect 62468 27132 69356 27188
rect 69412 27132 69422 27188
rect 6738 27020 6748 27076
rect 6804 27020 10108 27076
rect 10164 27020 10174 27076
rect 19954 27020 19964 27076
rect 20020 27020 20748 27076
rect 20804 27020 20814 27076
rect 21634 27020 21644 27076
rect 21700 27020 23548 27076
rect 23604 27020 23614 27076
rect 24556 26964 24612 27132
rect 27010 27020 27020 27076
rect 27076 27020 27468 27076
rect 27524 27020 27534 27076
rect 29810 27020 29820 27076
rect 29876 27020 31724 27076
rect 31780 27020 34300 27076
rect 34356 27020 34366 27076
rect 34738 27020 34748 27076
rect 34804 27020 37660 27076
rect 37716 27020 37726 27076
rect 37874 27020 37884 27076
rect 37940 27020 39340 27076
rect 39396 27020 39406 27076
rect 41346 27020 41356 27076
rect 41412 27020 43484 27076
rect 43540 27020 46844 27076
rect 46900 27020 46910 27076
rect 50372 27020 52836 27076
rect 60274 27020 60284 27076
rect 60340 27020 61628 27076
rect 61684 27020 61694 27076
rect 72146 27020 72156 27076
rect 72212 27020 72604 27076
rect 72660 27020 72670 27076
rect 50372 26964 50428 27020
rect 52780 26964 52836 27020
rect 16818 26908 16828 26964
rect 16884 26908 17388 26964
rect 17444 26908 21084 26964
rect 21140 26908 21150 26964
rect 21410 26908 21420 26964
rect 21476 26908 22652 26964
rect 22708 26908 22718 26964
rect 24546 26908 24556 26964
rect 24612 26908 25564 26964
rect 25620 26908 25630 26964
rect 30370 26908 30380 26964
rect 30436 26908 31276 26964
rect 31332 26908 35756 26964
rect 35812 26908 35822 26964
rect 39340 26908 39900 26964
rect 39956 26908 39966 26964
rect 41682 26908 41692 26964
rect 41748 26908 43372 26964
rect 43428 26908 43438 26964
rect 44818 26908 44828 26964
rect 44884 26908 45500 26964
rect 45556 26908 45566 26964
rect 45826 26908 45836 26964
rect 45892 26908 50428 26964
rect 50642 26908 50652 26964
rect 50708 26908 51100 26964
rect 51156 26908 52556 26964
rect 52612 26908 52622 26964
rect 52780 26908 56700 26964
rect 56756 26908 56766 26964
rect 57138 26908 57148 26964
rect 57204 26908 61292 26964
rect 61348 26908 61358 26964
rect 65314 26908 65324 26964
rect 65380 26908 66556 26964
rect 66612 26908 66622 26964
rect 68674 26908 68684 26964
rect 68740 26908 69356 26964
rect 69412 26908 77756 26964
rect 77812 26908 77822 26964
rect 39340 26852 39396 26908
rect 3332 26796 32732 26852
rect 32788 26796 32798 26852
rect 39330 26796 39340 26852
rect 39396 26796 39406 26852
rect 39778 26796 39788 26852
rect 39844 26796 40292 26852
rect 47282 26796 47292 26852
rect 47348 26796 48412 26852
rect 48468 26796 48478 26852
rect 49186 26796 49196 26852
rect 49252 26796 50540 26852
rect 50596 26796 51660 26852
rect 51716 26796 53116 26852
rect 53172 26796 53182 26852
rect 53554 26796 53564 26852
rect 53620 26796 61628 26852
rect 61684 26796 61694 26852
rect 3332 26740 3388 26796
rect 1810 26684 1820 26740
rect 1876 26684 3388 26740
rect 9874 26684 9884 26740
rect 9940 26684 11228 26740
rect 11284 26684 11788 26740
rect 11844 26684 11854 26740
rect 21074 26684 21084 26740
rect 21140 26684 21868 26740
rect 21924 26684 21934 26740
rect 28578 26684 28588 26740
rect 28644 26684 35532 26740
rect 35588 26684 36316 26740
rect 36372 26684 36382 26740
rect 38770 26684 38780 26740
rect 38836 26684 39676 26740
rect 39732 26684 39742 26740
rect 20522 26628 20532 26684
rect 20588 26628 20636 26684
rect 20692 26628 20740 26684
rect 20796 26628 20806 26684
rect 39842 26628 39852 26684
rect 39908 26628 39956 26684
rect 40012 26628 40060 26684
rect 40116 26628 40126 26684
rect 29698 26572 29708 26628
rect 29764 26572 35308 26628
rect 35364 26572 35374 26628
rect 38658 26572 38668 26628
rect 38724 26572 39564 26628
rect 39620 26572 39630 26628
rect 40236 26516 40292 26796
rect 53564 26740 53620 26796
rect 44818 26684 44828 26740
rect 44884 26684 44894 26740
rect 47292 26684 47852 26740
rect 47908 26684 49532 26740
rect 49588 26684 53620 26740
rect 57138 26684 57148 26740
rect 57204 26684 58940 26740
rect 58996 26684 59006 26740
rect 19842 26460 19852 26516
rect 19908 26460 22092 26516
rect 22148 26460 33124 26516
rect 36642 26460 36652 26516
rect 36708 26460 38668 26516
rect 40114 26460 40124 26516
rect 40180 26460 40292 26516
rect 40674 26460 40684 26516
rect 40740 26460 42700 26516
rect 42756 26460 42766 26516
rect 8866 26348 8876 26404
rect 8932 26348 9884 26404
rect 9940 26348 10556 26404
rect 10612 26348 10622 26404
rect 26226 26348 26236 26404
rect 26292 26348 26908 26404
rect 27682 26348 27692 26404
rect 27748 26348 28252 26404
rect 28308 26348 28318 26404
rect 30706 26348 30716 26404
rect 30772 26348 31164 26404
rect 31220 26348 31230 26404
rect 31826 26348 31836 26404
rect 31892 26348 32620 26404
rect 32676 26348 32686 26404
rect 26852 26292 26908 26348
rect 33068 26292 33124 26460
rect 38612 26404 38668 26460
rect 44828 26404 44884 26684
rect 47292 26628 47348 26684
rect 59162 26628 59172 26684
rect 59228 26628 59276 26684
rect 59332 26628 59380 26684
rect 59436 26628 59446 26684
rect 78482 26628 78492 26684
rect 78548 26628 78596 26684
rect 78652 26628 78700 26684
rect 78756 26628 78766 26684
rect 47282 26572 47292 26628
rect 47348 26572 47358 26628
rect 70018 26572 70028 26628
rect 70084 26572 70364 26628
rect 70420 26572 70430 26628
rect 56690 26460 56700 26516
rect 56756 26460 58604 26516
rect 58660 26460 59948 26516
rect 60004 26460 60732 26516
rect 60788 26460 60798 26516
rect 61282 26460 61292 26516
rect 61348 26460 75628 26516
rect 75684 26460 75694 26516
rect 38612 26348 44884 26404
rect 47012 26348 55468 26404
rect 55524 26348 55534 26404
rect 65426 26348 65436 26404
rect 65492 26348 70812 26404
rect 70868 26348 70878 26404
rect 71026 26348 71036 26404
rect 71092 26348 73948 26404
rect 74004 26348 74014 26404
rect 47012 26292 47068 26348
rect 8082 26236 8092 26292
rect 8148 26236 9548 26292
rect 9604 26236 11564 26292
rect 11620 26236 11630 26292
rect 19394 26236 19404 26292
rect 19460 26236 19852 26292
rect 19908 26236 20076 26292
rect 20132 26236 26684 26292
rect 26740 26236 26750 26292
rect 26852 26236 27132 26292
rect 27188 26236 27804 26292
rect 27860 26236 29372 26292
rect 29428 26236 29438 26292
rect 33058 26236 33068 26292
rect 33124 26236 33134 26292
rect 33282 26236 33292 26292
rect 33348 26236 38668 26292
rect 39666 26236 39676 26292
rect 39732 26236 40684 26292
rect 40740 26236 47068 26292
rect 50194 26236 50204 26292
rect 50260 26236 50428 26292
rect 50484 26236 52108 26292
rect 52164 26236 52174 26292
rect 52658 26236 52668 26292
rect 52724 26236 55580 26292
rect 55636 26236 55646 26292
rect 58930 26236 58940 26292
rect 58996 26236 59724 26292
rect 59780 26236 59790 26292
rect 62178 26236 62188 26292
rect 62244 26236 63308 26292
rect 63364 26236 63374 26292
rect 69122 26236 69132 26292
rect 69188 26236 69580 26292
rect 69636 26236 69646 26292
rect 38612 26180 38668 26236
rect 18722 26124 18732 26180
rect 18788 26124 37604 26180
rect 38612 26124 43932 26180
rect 43988 26124 43998 26180
rect 48178 26124 48188 26180
rect 48244 26124 49084 26180
rect 49140 26124 49308 26180
rect 49364 26124 49374 26180
rect 69458 26124 69468 26180
rect 69524 26124 69916 26180
rect 69972 26124 69982 26180
rect 70466 26124 70476 26180
rect 70532 26124 72492 26180
rect 72548 26124 72558 26180
rect 75282 26124 75292 26180
rect 75348 26124 77084 26180
rect 77140 26124 77150 26180
rect 0 26068 800 26096
rect 0 26012 1932 26068
rect 1988 26012 1998 26068
rect 18162 26012 18172 26068
rect 18228 26012 19068 26068
rect 19124 26012 20076 26068
rect 20132 26012 20636 26068
rect 20692 26012 20702 26068
rect 21186 26012 21196 26068
rect 21252 26012 22428 26068
rect 22484 26012 22494 26068
rect 0 25984 800 26012
rect 37548 25956 37604 26124
rect 79200 26068 80000 26096
rect 38108 26012 40012 26068
rect 40068 26012 40348 26068
rect 40404 26012 40414 26068
rect 45714 26012 45724 26068
rect 45780 26012 46284 26068
rect 46340 26012 46350 26068
rect 48402 26012 48412 26068
rect 48468 26012 51492 26068
rect 68114 26012 68124 26068
rect 68180 26012 71932 26068
rect 71988 26012 71998 26068
rect 77970 26012 77980 26068
rect 78036 26012 80000 26068
rect 38108 25956 38164 26012
rect 18722 25900 18732 25956
rect 18788 25900 18956 25956
rect 19012 25900 19022 25956
rect 28018 25900 28028 25956
rect 28084 25900 28700 25956
rect 28756 25900 28766 25956
rect 37538 25900 37548 25956
rect 37604 25900 37614 25956
rect 38098 25900 38108 25956
rect 38164 25900 38174 25956
rect 38658 25900 38668 25956
rect 38724 25900 39004 25956
rect 39060 25900 39070 25956
rect 39340 25900 43372 25956
rect 43428 25900 43438 25956
rect 43810 25900 43820 25956
rect 43876 25900 45052 25956
rect 45108 25900 45118 25956
rect 10862 25844 10872 25900
rect 10928 25844 10976 25900
rect 11032 25844 11080 25900
rect 11136 25844 11146 25900
rect 30182 25844 30192 25900
rect 30248 25844 30296 25900
rect 30352 25844 30400 25900
rect 30456 25844 30466 25900
rect 39340 25844 39396 25900
rect 49502 25844 49512 25900
rect 49568 25844 49616 25900
rect 49672 25844 49720 25900
rect 49776 25844 49786 25900
rect 28578 25788 28588 25844
rect 28644 25788 28654 25844
rect 37986 25788 37996 25844
rect 38052 25788 38444 25844
rect 38500 25788 38510 25844
rect 38770 25788 38780 25844
rect 38836 25788 39396 25844
rect 39554 25788 39564 25844
rect 39620 25788 41916 25844
rect 41972 25788 41982 25844
rect 44930 25788 44940 25844
rect 44996 25788 45612 25844
rect 45668 25788 45678 25844
rect 50642 25788 50652 25844
rect 50708 25788 51212 25844
rect 51268 25788 51278 25844
rect 12002 25676 12012 25732
rect 12068 25676 12908 25732
rect 12964 25676 16492 25732
rect 16548 25676 16558 25732
rect 28588 25620 28644 25788
rect 51436 25732 51492 26012
rect 79200 25984 80000 26012
rect 53778 25900 53788 25956
rect 53844 25900 64540 25956
rect 64596 25900 64606 25956
rect 72370 25900 72380 25956
rect 72436 25900 72446 25956
rect 68822 25844 68832 25900
rect 68888 25844 68936 25900
rect 68992 25844 69040 25900
rect 69096 25844 69106 25900
rect 72380 25844 72436 25900
rect 52882 25788 52892 25844
rect 52948 25788 56924 25844
rect 56980 25788 56990 25844
rect 69794 25788 69804 25844
rect 69860 25788 72436 25844
rect 35186 25676 35196 25732
rect 35252 25676 47516 25732
rect 47572 25676 47852 25732
rect 47908 25676 47918 25732
rect 51436 25676 63084 25732
rect 63140 25676 63150 25732
rect 68562 25676 68572 25732
rect 68628 25676 72156 25732
rect 72212 25676 72222 25732
rect 76626 25676 76636 25732
rect 76692 25676 77308 25732
rect 77364 25676 77980 25732
rect 78036 25676 78046 25732
rect 15474 25564 15484 25620
rect 15540 25564 15820 25620
rect 15876 25564 15886 25620
rect 24210 25564 24220 25620
rect 24276 25564 25732 25620
rect 26338 25564 26348 25620
rect 26404 25564 26908 25620
rect 26964 25564 26974 25620
rect 27244 25564 28644 25620
rect 29250 25564 29260 25620
rect 29316 25564 30268 25620
rect 30324 25564 34412 25620
rect 34468 25564 34478 25620
rect 35522 25564 35532 25620
rect 35588 25564 35756 25620
rect 35812 25564 41356 25620
rect 41412 25564 41422 25620
rect 43474 25564 43484 25620
rect 43540 25564 47068 25620
rect 15484 25508 15540 25564
rect 25676 25508 25732 25564
rect 27244 25508 27300 25564
rect 47012 25508 47068 25564
rect 50540 25564 62412 25620
rect 62468 25564 62478 25620
rect 69346 25564 69356 25620
rect 69412 25564 71148 25620
rect 71204 25564 73164 25620
rect 73220 25564 73230 25620
rect 50540 25508 50596 25564
rect 12786 25452 12796 25508
rect 12852 25452 13580 25508
rect 13636 25452 14588 25508
rect 14644 25452 14654 25508
rect 15092 25452 15540 25508
rect 15698 25452 15708 25508
rect 15764 25452 16716 25508
rect 16772 25452 16782 25508
rect 20738 25452 20748 25508
rect 20804 25452 21644 25508
rect 21700 25452 21710 25508
rect 22642 25452 22652 25508
rect 22708 25452 22988 25508
rect 23044 25452 25004 25508
rect 25060 25452 25070 25508
rect 25676 25452 27300 25508
rect 27458 25452 27468 25508
rect 27524 25452 28476 25508
rect 28532 25452 31052 25508
rect 31108 25452 31118 25508
rect 32722 25452 32732 25508
rect 32788 25452 38780 25508
rect 38836 25452 38846 25508
rect 39778 25452 39788 25508
rect 39844 25452 39854 25508
rect 44258 25452 44268 25508
rect 44324 25452 44828 25508
rect 44884 25452 44894 25508
rect 47012 25452 50596 25508
rect 53218 25452 53228 25508
rect 53284 25452 53676 25508
rect 53732 25452 54572 25508
rect 54628 25452 54638 25508
rect 65202 25452 65212 25508
rect 65268 25452 66220 25508
rect 66276 25452 67340 25508
rect 67396 25452 68348 25508
rect 68404 25452 68414 25508
rect 70690 25452 70700 25508
rect 70756 25452 72380 25508
rect 72436 25452 72446 25508
rect 72706 25452 72716 25508
rect 72772 25452 73500 25508
rect 73556 25452 75292 25508
rect 75348 25452 75358 25508
rect 75506 25452 75516 25508
rect 75572 25452 76860 25508
rect 76916 25452 76926 25508
rect 15092 25396 15148 25452
rect 39788 25396 39844 25452
rect 6066 25340 6076 25396
rect 6132 25340 12572 25396
rect 12628 25340 15148 25396
rect 22306 25340 22316 25396
rect 22372 25340 25900 25396
rect 25956 25340 25966 25396
rect 26898 25340 26908 25396
rect 26964 25340 29596 25396
rect 29652 25340 29662 25396
rect 29810 25340 29820 25396
rect 29876 25340 33404 25396
rect 33460 25340 38108 25396
rect 38164 25340 38174 25396
rect 38546 25340 38556 25396
rect 38612 25340 38892 25396
rect 38948 25340 38958 25396
rect 39106 25340 39116 25396
rect 39172 25340 39844 25396
rect 40338 25340 40348 25396
rect 40404 25340 40908 25396
rect 40964 25340 40974 25396
rect 50754 25340 50764 25396
rect 50820 25340 50830 25396
rect 65986 25340 65996 25396
rect 66052 25340 66780 25396
rect 66836 25340 69356 25396
rect 69412 25340 69422 25396
rect 69570 25340 69580 25396
rect 69636 25340 77420 25396
rect 77476 25340 78204 25396
rect 78260 25340 78270 25396
rect 50764 25284 50820 25340
rect 4274 25228 4284 25284
rect 4340 25228 4844 25284
rect 4900 25228 21980 25284
rect 22036 25228 22046 25284
rect 28130 25228 28140 25284
rect 28196 25228 28700 25284
rect 28756 25228 28924 25284
rect 28980 25228 29708 25284
rect 29764 25228 29774 25284
rect 30146 25228 30156 25284
rect 30212 25228 38220 25284
rect 38276 25228 38286 25284
rect 38444 25228 45948 25284
rect 46004 25228 46014 25284
rect 47730 25228 47740 25284
rect 47796 25228 50820 25284
rect 51762 25228 51772 25284
rect 51828 25228 52892 25284
rect 52948 25228 52958 25284
rect 54114 25228 54124 25284
rect 54180 25228 55132 25284
rect 55188 25228 57372 25284
rect 57428 25228 57438 25284
rect 57810 25228 57820 25284
rect 57876 25228 59388 25284
rect 59444 25228 59454 25284
rect 68226 25228 68236 25284
rect 68292 25228 68302 25284
rect 68562 25228 68572 25284
rect 68628 25228 69972 25284
rect 70130 25228 70140 25284
rect 70196 25228 72156 25284
rect 72212 25228 72222 25284
rect 72380 25228 73276 25284
rect 73332 25228 73342 25284
rect 38444 25172 38500 25228
rect 68236 25172 68292 25228
rect 8418 25116 8428 25172
rect 8484 25116 9660 25172
rect 9716 25116 9726 25172
rect 14802 25116 14812 25172
rect 14868 25116 15484 25172
rect 15540 25116 15550 25172
rect 27234 25116 27244 25172
rect 27300 25116 38500 25172
rect 40898 25116 40908 25172
rect 40964 25116 41692 25172
rect 41748 25116 41758 25172
rect 44146 25116 44156 25172
rect 44212 25116 56308 25172
rect 64754 25116 64764 25172
rect 64820 25116 65996 25172
rect 66052 25116 68292 25172
rect 69916 25172 69972 25228
rect 72380 25172 72436 25228
rect 69916 25116 70476 25172
rect 70532 25116 70542 25172
rect 72258 25116 72268 25172
rect 72324 25116 72436 25172
rect 20522 25060 20532 25116
rect 20588 25060 20636 25116
rect 20692 25060 20740 25116
rect 20796 25060 20806 25116
rect 39842 25060 39852 25116
rect 39908 25060 39956 25116
rect 40012 25060 40060 25116
rect 40116 25060 40126 25116
rect 28914 25004 28924 25060
rect 28980 25004 29932 25060
rect 29988 25004 35308 25060
rect 35364 25004 37212 25060
rect 37268 25004 37278 25060
rect 44492 25004 50764 25060
rect 50820 25004 50830 25060
rect 53890 25004 53900 25060
rect 53956 25004 55132 25060
rect 55188 25004 55198 25060
rect 44492 24948 44548 25004
rect 56252 24948 56308 25116
rect 59162 25060 59172 25116
rect 59228 25060 59276 25116
rect 59332 25060 59380 25116
rect 59436 25060 59446 25116
rect 78482 25060 78492 25116
rect 78548 25060 78596 25116
rect 78652 25060 78700 25116
rect 78756 25060 78766 25116
rect 59602 25004 59612 25060
rect 59668 25004 59948 25060
rect 60004 25004 60014 25060
rect 9538 24892 9548 24948
rect 9604 24892 10220 24948
rect 10276 24892 14812 24948
rect 14868 24892 14878 24948
rect 15810 24892 15820 24948
rect 15876 24892 16716 24948
rect 16772 24892 16782 24948
rect 19730 24892 19740 24948
rect 19796 24892 29036 24948
rect 29092 24892 29102 24948
rect 29586 24892 29596 24948
rect 29652 24892 30044 24948
rect 30100 24892 44548 24948
rect 46610 24892 46620 24948
rect 46676 24892 48636 24948
rect 48692 24892 48702 24948
rect 48860 24892 54292 24948
rect 56252 24892 73332 24948
rect 73714 24892 73724 24948
rect 73780 24892 74620 24948
rect 74676 24892 74686 24948
rect 48860 24836 48916 24892
rect 4722 24780 4732 24836
rect 4788 24780 5516 24836
rect 5572 24780 5582 24836
rect 15484 24780 20188 24836
rect 20244 24780 20254 24836
rect 21298 24780 21308 24836
rect 21364 24780 27468 24836
rect 27524 24780 27534 24836
rect 27794 24780 27804 24836
rect 27860 24780 28140 24836
rect 28196 24780 28206 24836
rect 33618 24780 33628 24836
rect 33684 24780 34076 24836
rect 34132 24780 34142 24836
rect 38434 24780 38444 24836
rect 38500 24780 40012 24836
rect 40068 24780 40908 24836
rect 40964 24780 40974 24836
rect 41580 24780 48916 24836
rect 51650 24780 51660 24836
rect 51716 24780 53788 24836
rect 53844 24780 53854 24836
rect 15484 24612 15540 24780
rect 18722 24668 18732 24724
rect 18788 24668 19404 24724
rect 19460 24668 19470 24724
rect 22316 24668 23548 24724
rect 23604 24668 24444 24724
rect 24500 24668 24510 24724
rect 27906 24668 27916 24724
rect 27972 24668 28588 24724
rect 28644 24668 29036 24724
rect 29092 24668 29372 24724
rect 29428 24668 29438 24724
rect 33730 24668 33740 24724
rect 33796 24668 34412 24724
rect 34468 24668 34478 24724
rect 38210 24668 38220 24724
rect 38276 24668 39340 24724
rect 39396 24668 39676 24724
rect 39732 24668 39742 24724
rect 22316 24612 22372 24668
rect 41580 24612 41636 24780
rect 42466 24668 42476 24724
rect 42532 24668 43036 24724
rect 43092 24668 43102 24724
rect 45266 24668 45276 24724
rect 45332 24668 46172 24724
rect 46228 24668 46238 24724
rect 46946 24668 46956 24724
rect 47012 24668 52780 24724
rect 52836 24668 53900 24724
rect 53956 24668 53966 24724
rect 4834 24556 4844 24612
rect 4900 24556 6188 24612
rect 6244 24556 8428 24612
rect 8484 24556 8494 24612
rect 13458 24556 13468 24612
rect 13524 24556 14252 24612
rect 14308 24556 14318 24612
rect 15474 24556 15484 24612
rect 15540 24556 15550 24612
rect 16594 24556 16604 24612
rect 16660 24556 17724 24612
rect 17780 24556 17790 24612
rect 17938 24556 17948 24612
rect 18004 24556 22372 24612
rect 31938 24556 31948 24612
rect 32004 24556 33068 24612
rect 33124 24556 41636 24612
rect 44034 24556 44044 24612
rect 44100 24556 44716 24612
rect 44772 24556 45388 24612
rect 45444 24556 45836 24612
rect 45892 24556 45902 24612
rect 54236 24500 54292 24892
rect 73276 24836 73332 24892
rect 56242 24780 56252 24836
rect 56308 24780 57932 24836
rect 57988 24780 57998 24836
rect 58380 24780 59612 24836
rect 59668 24780 60396 24836
rect 60452 24780 60462 24836
rect 69010 24780 69020 24836
rect 69076 24780 71260 24836
rect 71316 24780 73052 24836
rect 73108 24780 73118 24836
rect 73276 24780 73836 24836
rect 73892 24780 73902 24836
rect 58380 24724 58436 24780
rect 54786 24668 54796 24724
rect 54852 24668 55356 24724
rect 55412 24668 56588 24724
rect 56644 24668 56654 24724
rect 57250 24668 57260 24724
rect 57316 24668 58436 24724
rect 58706 24668 58716 24724
rect 58772 24668 59724 24724
rect 59780 24668 59790 24724
rect 63634 24668 63644 24724
rect 63700 24668 64876 24724
rect 64932 24668 64942 24724
rect 71586 24668 71596 24724
rect 71652 24668 72604 24724
rect 72660 24668 72670 24724
rect 57810 24556 57820 24612
rect 57876 24556 59836 24612
rect 59892 24556 59902 24612
rect 61842 24556 61852 24612
rect 61908 24556 62300 24612
rect 62356 24556 62748 24612
rect 62804 24556 62814 24612
rect 11666 24444 11676 24500
rect 11732 24444 13916 24500
rect 13972 24444 13982 24500
rect 16706 24444 16716 24500
rect 16772 24444 19068 24500
rect 19124 24444 19134 24500
rect 23426 24444 23436 24500
rect 23492 24444 28924 24500
rect 28980 24444 28990 24500
rect 33618 24444 33628 24500
rect 33684 24444 36316 24500
rect 36372 24444 36382 24500
rect 37426 24444 37436 24500
rect 37492 24444 37884 24500
rect 37940 24444 40180 24500
rect 40898 24444 40908 24500
rect 40964 24444 41356 24500
rect 41412 24444 41422 24500
rect 50754 24444 50764 24500
rect 50820 24444 51100 24500
rect 51156 24444 51166 24500
rect 54236 24444 62188 24500
rect 17490 24332 17500 24388
rect 17556 24332 19628 24388
rect 19684 24332 19694 24388
rect 22082 24332 22092 24388
rect 22148 24332 23884 24388
rect 23940 24332 23950 24388
rect 10862 24276 10872 24332
rect 10928 24276 10976 24332
rect 11032 24276 11080 24332
rect 11136 24276 11146 24332
rect 30182 24276 30192 24332
rect 30248 24276 30296 24332
rect 30352 24276 30400 24332
rect 30456 24276 30466 24332
rect 36316 24276 36372 24444
rect 40124 24388 40180 24444
rect 51100 24388 51156 24444
rect 62132 24388 62188 24444
rect 40124 24332 41804 24388
rect 41860 24332 41870 24388
rect 51100 24332 54796 24388
rect 54852 24332 54862 24388
rect 56354 24332 56364 24388
rect 56420 24332 59948 24388
rect 60004 24332 61628 24388
rect 61684 24332 61694 24388
rect 62132 24332 66276 24388
rect 49502 24276 49512 24332
rect 49568 24276 49616 24332
rect 49672 24276 49720 24332
rect 49776 24276 49786 24332
rect 14802 24220 14812 24276
rect 14868 24220 15484 24276
rect 15540 24220 15550 24276
rect 18722 24220 18732 24276
rect 18788 24220 19852 24276
rect 19908 24220 19918 24276
rect 22530 24220 22540 24276
rect 22596 24220 25228 24276
rect 25284 24220 26012 24276
rect 26068 24220 26078 24276
rect 36316 24220 41300 24276
rect 41458 24220 41468 24276
rect 41524 24220 42700 24276
rect 42756 24220 43260 24276
rect 43316 24220 43326 24276
rect 50306 24220 50316 24276
rect 50372 24220 54460 24276
rect 54516 24220 54526 24276
rect 57810 24220 57820 24276
rect 57876 24220 58828 24276
rect 58884 24220 58894 24276
rect 41244 24164 41300 24220
rect 43260 24164 43316 24220
rect 66220 24164 66276 24332
rect 68822 24276 68832 24332
rect 68888 24276 68936 24332
rect 68992 24276 69040 24332
rect 69096 24276 69106 24332
rect 71810 24220 71820 24276
rect 71876 24220 72268 24276
rect 72324 24220 72334 24276
rect 4274 24108 4284 24164
rect 4340 24108 4844 24164
rect 4900 24108 31724 24164
rect 31780 24108 31790 24164
rect 34178 24108 34188 24164
rect 34244 24108 36316 24164
rect 36372 24108 36382 24164
rect 38546 24108 38556 24164
rect 38612 24108 39900 24164
rect 39956 24108 40908 24164
rect 40964 24108 40974 24164
rect 41244 24108 42588 24164
rect 42644 24108 42654 24164
rect 43260 24108 61404 24164
rect 61460 24108 61470 24164
rect 66220 24108 71708 24164
rect 71764 24108 73052 24164
rect 73108 24108 73118 24164
rect 17938 23996 17948 24052
rect 18004 23996 18396 24052
rect 18452 23996 18462 24052
rect 21746 23996 21756 24052
rect 21812 23996 23100 24052
rect 23156 23996 23166 24052
rect 29810 23996 29820 24052
rect 29876 23996 30940 24052
rect 30996 23996 33852 24052
rect 33908 23996 35532 24052
rect 35588 23996 35598 24052
rect 37202 23996 37212 24052
rect 37268 23996 44044 24052
rect 44100 23996 44110 24052
rect 49410 23996 49420 24052
rect 49476 23996 50876 24052
rect 50932 23996 50942 24052
rect 54114 23996 54124 24052
rect 54180 23996 56252 24052
rect 56308 23996 57036 24052
rect 57092 23996 58044 24052
rect 58100 23996 58380 24052
rect 58436 23996 58446 24052
rect 60386 23996 60396 24052
rect 60452 23996 64764 24052
rect 64820 23996 64830 24052
rect 1810 23884 1820 23940
rect 1876 23884 5740 23940
rect 5796 23884 5806 23940
rect 16146 23884 16156 23940
rect 16212 23884 16716 23940
rect 16772 23884 20524 23940
rect 20580 23884 20590 23940
rect 21298 23884 21308 23940
rect 21364 23884 21980 23940
rect 22036 23884 23436 23940
rect 23492 23884 23502 23940
rect 26124 23884 28308 23940
rect 28466 23884 28476 23940
rect 28532 23884 29708 23940
rect 29764 23884 30492 23940
rect 30548 23884 30558 23940
rect 33394 23884 33404 23940
rect 33460 23884 34524 23940
rect 34580 23884 34590 23940
rect 37650 23884 37660 23940
rect 37716 23884 38780 23940
rect 38836 23884 38846 23940
rect 39106 23884 39116 23940
rect 39172 23884 39508 23940
rect 40450 23884 40460 23940
rect 40516 23884 41692 23940
rect 41748 23884 41758 23940
rect 43026 23884 43036 23940
rect 43092 23884 43708 23940
rect 43764 23884 43774 23940
rect 53218 23884 53228 23940
rect 53284 23884 54460 23940
rect 54516 23884 55468 23940
rect 55524 23884 55534 23940
rect 59938 23884 59948 23940
rect 60004 23884 61292 23940
rect 61348 23884 61358 23940
rect 20178 23772 20188 23828
rect 20244 23772 21756 23828
rect 21812 23772 21822 23828
rect 22978 23772 22988 23828
rect 23044 23772 23324 23828
rect 23380 23772 23390 23828
rect 26124 23716 26180 23884
rect 26338 23772 26348 23828
rect 26404 23772 26908 23828
rect 21858 23660 21868 23716
rect 21924 23660 23436 23716
rect 23492 23660 26180 23716
rect 26852 23716 26908 23772
rect 28252 23716 28308 23884
rect 39452 23828 39508 23884
rect 30594 23772 30604 23828
rect 30660 23772 31164 23828
rect 31220 23772 32396 23828
rect 32452 23772 32462 23828
rect 38098 23772 38108 23828
rect 38164 23772 39228 23828
rect 39284 23772 39294 23828
rect 39452 23772 40684 23828
rect 40740 23772 40750 23828
rect 41234 23772 41244 23828
rect 41300 23772 43596 23828
rect 43652 23772 43662 23828
rect 50372 23772 51660 23828
rect 51716 23772 51726 23828
rect 51986 23772 51996 23828
rect 52052 23772 57372 23828
rect 57428 23772 59052 23828
rect 59108 23772 59118 23828
rect 50372 23716 50428 23772
rect 26852 23660 28196 23716
rect 28252 23660 50428 23716
rect 51314 23660 51324 23716
rect 51380 23660 57932 23716
rect 57988 23660 58492 23716
rect 58548 23660 58558 23716
rect 58940 23660 59388 23716
rect 59444 23660 60620 23716
rect 60676 23660 60686 23716
rect 0 23604 800 23632
rect 28140 23604 28196 23660
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 15362 23548 15372 23604
rect 15428 23548 15820 23604
rect 15876 23548 15886 23604
rect 21410 23548 21420 23604
rect 21476 23548 22988 23604
rect 23044 23548 23054 23604
rect 23762 23548 23772 23604
rect 23828 23548 25452 23604
rect 25508 23548 25518 23604
rect 25666 23548 25676 23604
rect 25732 23548 27244 23604
rect 27300 23548 27310 23604
rect 28140 23548 28364 23604
rect 28420 23548 28430 23604
rect 33394 23548 33404 23604
rect 33460 23548 33684 23604
rect 35970 23548 35980 23604
rect 36036 23548 37100 23604
rect 37156 23548 38108 23604
rect 38164 23548 38174 23604
rect 40236 23548 43204 23604
rect 43362 23548 43372 23604
rect 43428 23548 44156 23604
rect 44212 23548 44222 23604
rect 44380 23548 47516 23604
rect 47572 23548 47582 23604
rect 0 23520 800 23548
rect 20522 23492 20532 23548
rect 20588 23492 20636 23548
rect 20692 23492 20740 23548
rect 20796 23492 20806 23548
rect 22204 23492 22260 23548
rect 33618 23492 33628 23548
rect 33684 23492 33694 23548
rect 39842 23492 39852 23548
rect 39908 23492 39956 23548
rect 40012 23492 40060 23548
rect 40116 23492 40126 23548
rect 3332 23436 20188 23492
rect 20244 23436 20254 23492
rect 22194 23436 22204 23492
rect 22260 23436 22270 23492
rect 25554 23436 25564 23492
rect 25620 23436 26124 23492
rect 26180 23436 26684 23492
rect 26740 23436 27916 23492
rect 27972 23436 27982 23492
rect 31490 23436 31500 23492
rect 31556 23436 32620 23492
rect 32676 23436 33460 23492
rect 34850 23436 34860 23492
rect 34916 23436 36540 23492
rect 36596 23436 36606 23492
rect 39330 23436 39340 23492
rect 39396 23436 39732 23492
rect 3332 23380 3388 23436
rect 33404 23380 33460 23436
rect 39676 23380 39732 23436
rect 40236 23380 40292 23548
rect 43148 23492 43204 23548
rect 44380 23492 44436 23548
rect 58940 23492 58996 23660
rect 66220 23604 66276 24108
rect 70242 23884 70252 23940
rect 70308 23884 71036 23940
rect 71092 23884 72604 23940
rect 72660 23884 72670 23940
rect 67106 23772 67116 23828
rect 67172 23772 69580 23828
rect 69636 23772 72044 23828
rect 72100 23772 72110 23828
rect 72258 23772 72268 23828
rect 72324 23772 72828 23828
rect 72884 23772 72894 23828
rect 75394 23660 75404 23716
rect 75460 23660 78932 23716
rect 78876 23604 78932 23660
rect 79200 23604 80000 23632
rect 60050 23548 60060 23604
rect 60116 23548 64204 23604
rect 64260 23548 65436 23604
rect 65492 23548 65502 23604
rect 66210 23548 66220 23604
rect 66276 23548 66286 23604
rect 71810 23548 71820 23604
rect 71876 23548 72156 23604
rect 72212 23548 72222 23604
rect 72370 23548 72380 23604
rect 72436 23548 74284 23604
rect 74340 23548 74350 23604
rect 78876 23548 80000 23604
rect 59162 23492 59172 23548
rect 59228 23492 59276 23548
rect 59332 23492 59380 23548
rect 59436 23492 59446 23548
rect 78482 23492 78492 23548
rect 78548 23492 78596 23548
rect 78652 23492 78700 23548
rect 78756 23492 78766 23548
rect 79200 23520 80000 23548
rect 43148 23436 44436 23492
rect 45602 23436 45612 23492
rect 45668 23436 50652 23492
rect 50708 23436 50718 23492
rect 54450 23436 54460 23492
rect 54516 23436 58996 23492
rect 66882 23436 66892 23492
rect 66948 23436 68908 23492
rect 68964 23436 72268 23492
rect 72324 23436 72334 23492
rect 73602 23436 73612 23492
rect 73668 23436 74060 23492
rect 74116 23436 74844 23492
rect 74900 23436 74910 23492
rect 2370 23324 2380 23380
rect 2436 23324 3388 23380
rect 5730 23324 5740 23380
rect 5796 23324 8652 23380
rect 8708 23324 9660 23380
rect 9716 23324 9726 23380
rect 16258 23324 16268 23380
rect 16324 23324 17500 23380
rect 17556 23324 17566 23380
rect 26450 23324 26460 23380
rect 26516 23324 27244 23380
rect 27300 23324 27310 23380
rect 31602 23324 31612 23380
rect 31668 23324 32060 23380
rect 32116 23324 33180 23380
rect 33236 23324 33246 23380
rect 33404 23324 36428 23380
rect 36484 23324 39620 23380
rect 39676 23324 40292 23380
rect 40786 23324 40796 23380
rect 40852 23324 41468 23380
rect 41524 23324 42812 23380
rect 42868 23324 42878 23380
rect 44370 23324 44380 23380
rect 44436 23324 45388 23380
rect 45444 23324 45454 23380
rect 46162 23324 46172 23380
rect 46228 23324 47516 23380
rect 47572 23324 50092 23380
rect 50148 23324 51100 23380
rect 51156 23324 51660 23380
rect 51716 23324 51726 23380
rect 60610 23324 60620 23380
rect 60676 23324 61740 23380
rect 61796 23324 61806 23380
rect 65650 23324 65660 23380
rect 65716 23324 67508 23380
rect 69682 23324 69692 23380
rect 69748 23324 72156 23380
rect 72212 23324 72222 23380
rect 39564 23268 39620 23324
rect 67452 23268 67508 23324
rect 7186 23212 7196 23268
rect 7252 23212 9100 23268
rect 9156 23212 9166 23268
rect 15092 23212 16044 23268
rect 16100 23212 16110 23268
rect 19058 23212 19068 23268
rect 19124 23212 19740 23268
rect 19796 23212 19806 23268
rect 28354 23212 28364 23268
rect 28420 23212 29260 23268
rect 29316 23212 30380 23268
rect 30436 23212 30446 23268
rect 31938 23212 31948 23268
rect 32004 23212 33292 23268
rect 33348 23212 33358 23268
rect 36642 23212 36652 23268
rect 36708 23212 38780 23268
rect 38836 23212 39340 23268
rect 39396 23212 39406 23268
rect 39564 23212 39676 23268
rect 39732 23212 42476 23268
rect 42532 23212 42542 23268
rect 47170 23212 47180 23268
rect 47236 23212 47964 23268
rect 48020 23212 48030 23268
rect 61170 23212 61180 23268
rect 61236 23212 62188 23268
rect 62290 23212 62300 23268
rect 62356 23212 63196 23268
rect 63252 23212 65548 23268
rect 65604 23212 65614 23268
rect 67442 23212 67452 23268
rect 67508 23212 71484 23268
rect 71540 23212 71550 23268
rect 72706 23212 72716 23268
rect 72772 23212 73724 23268
rect 73780 23212 73790 23268
rect 8642 22988 8652 23044
rect 8708 22988 15036 23044
rect 15092 22988 15148 23212
rect 62132 23156 62188 23212
rect 15362 23100 15372 23156
rect 15428 23100 15932 23156
rect 15988 23100 15998 23156
rect 19842 23100 19852 23156
rect 19908 23100 25676 23156
rect 25732 23100 25742 23156
rect 28242 23100 28252 23156
rect 28308 23100 30716 23156
rect 30772 23100 30782 23156
rect 32498 23100 32508 23156
rect 32564 23100 34636 23156
rect 34692 23100 35420 23156
rect 35476 23100 40124 23156
rect 40180 23100 41020 23156
rect 41076 23100 41086 23156
rect 51314 23100 51324 23156
rect 51380 23100 51660 23156
rect 51716 23100 51726 23156
rect 53554 23100 53564 23156
rect 53620 23100 54236 23156
rect 54292 23100 54302 23156
rect 57698 23100 57708 23156
rect 57764 23100 59500 23156
rect 59556 23100 59566 23156
rect 60722 23100 60732 23156
rect 60788 23100 61292 23156
rect 61348 23100 61964 23156
rect 62020 23100 62030 23156
rect 62132 23100 62636 23156
rect 62692 23100 62702 23156
rect 63298 23100 63308 23156
rect 63364 23100 68348 23156
rect 68404 23100 68414 23156
rect 69234 23100 69244 23156
rect 69300 23100 70588 23156
rect 70644 23100 70654 23156
rect 72482 23100 72492 23156
rect 72548 23100 72828 23156
rect 72884 23100 72894 23156
rect 15474 22988 15484 23044
rect 15540 22988 16604 23044
rect 16660 22988 16670 23044
rect 21186 22988 21196 23044
rect 21252 22988 26012 23044
rect 26068 22988 26078 23044
rect 28802 22988 28812 23044
rect 28868 22988 34244 23044
rect 38882 22988 38892 23044
rect 38948 22988 39900 23044
rect 39956 22988 39966 23044
rect 41234 22988 41244 23044
rect 41300 22988 41916 23044
rect 41972 22988 41982 23044
rect 43810 22988 43820 23044
rect 43876 22988 45500 23044
rect 45556 22988 45948 23044
rect 46004 22988 46014 23044
rect 49410 22988 49420 23044
rect 49476 22988 50988 23044
rect 51044 22988 51054 23044
rect 53890 22988 53900 23044
rect 53956 22988 56028 23044
rect 56084 22988 58156 23044
rect 58212 22988 58222 23044
rect 60162 22988 60172 23044
rect 60228 22988 62188 23044
rect 63746 22988 63756 23044
rect 63812 22988 65996 23044
rect 66052 22988 66062 23044
rect 67330 22988 67340 23044
rect 67396 22988 70364 23044
rect 70420 22988 70430 23044
rect 70802 22988 70812 23044
rect 70868 22988 76412 23044
rect 76468 22988 77196 23044
rect 77252 22988 77262 23044
rect 34188 22932 34244 22988
rect 62132 22932 62188 22988
rect 10210 22876 10220 22932
rect 10276 22876 13580 22932
rect 13636 22876 13646 22932
rect 18162 22876 18172 22932
rect 18228 22876 20300 22932
rect 20356 22876 26908 22932
rect 29026 22876 29036 22932
rect 29092 22876 30660 22932
rect 34178 22876 34188 22932
rect 34244 22876 34254 22932
rect 34402 22876 34412 22932
rect 34468 22876 36764 22932
rect 36820 22876 36830 22932
rect 38994 22876 39004 22932
rect 39060 22876 39788 22932
rect 39844 22876 50428 22932
rect 53554 22876 53564 22932
rect 53620 22876 54572 22932
rect 54628 22876 54638 22932
rect 62132 22876 65660 22932
rect 65716 22876 65726 22932
rect 68450 22876 68460 22932
rect 68516 22876 69916 22932
rect 69972 22876 69982 22932
rect 71586 22876 71596 22932
rect 71652 22876 72268 22932
rect 72324 22876 72334 22932
rect 26852 22820 26908 22876
rect 30604 22820 30660 22876
rect 26852 22764 27804 22820
rect 27860 22764 27870 22820
rect 28018 22764 28028 22820
rect 28084 22764 29148 22820
rect 29204 22764 29214 22820
rect 30604 22764 47068 22820
rect 47124 22764 47134 22820
rect 10862 22708 10872 22764
rect 10928 22708 10976 22764
rect 11032 22708 11080 22764
rect 11136 22708 11146 22764
rect 30182 22708 30192 22764
rect 30248 22708 30296 22764
rect 30352 22708 30400 22764
rect 30456 22708 30466 22764
rect 49502 22708 49512 22764
rect 49568 22708 49616 22764
rect 49672 22708 49720 22764
rect 49776 22708 49786 22764
rect 50372 22708 50428 22876
rect 71026 22764 71036 22820
rect 71092 22764 75628 22820
rect 75684 22764 76636 22820
rect 76692 22764 77644 22820
rect 77700 22764 77710 22820
rect 68822 22708 68832 22764
rect 68888 22708 68936 22764
rect 68992 22708 69040 22764
rect 69096 22708 69106 22764
rect 26852 22652 28084 22708
rect 26852 22596 26908 22652
rect 18722 22540 18732 22596
rect 18788 22540 19852 22596
rect 19908 22540 19918 22596
rect 26338 22540 26348 22596
rect 26404 22540 26908 22596
rect 28028 22596 28084 22652
rect 38612 22652 45164 22708
rect 45220 22652 46172 22708
rect 46228 22652 46238 22708
rect 50372 22652 57036 22708
rect 57092 22652 59948 22708
rect 60004 22652 60014 22708
rect 72258 22652 72268 22708
rect 72324 22652 76972 22708
rect 77028 22652 77980 22708
rect 78036 22652 78046 22708
rect 38612 22596 38668 22652
rect 28028 22540 38668 22596
rect 39666 22540 39676 22596
rect 39732 22540 40796 22596
rect 40852 22540 40862 22596
rect 43362 22540 43372 22596
rect 43428 22540 64708 22596
rect 64866 22540 64876 22596
rect 64932 22540 73164 22596
rect 73220 22540 73500 22596
rect 73556 22540 73566 22596
rect 18274 22428 18284 22484
rect 18340 22428 19404 22484
rect 19460 22428 19470 22484
rect 25778 22428 25788 22484
rect 25844 22428 26572 22484
rect 26628 22428 26638 22484
rect 27794 22428 27804 22484
rect 27860 22428 46620 22484
rect 46676 22428 54460 22484
rect 54516 22428 54526 22484
rect 54674 22428 54684 22484
rect 54740 22428 56140 22484
rect 56196 22428 56812 22484
rect 56868 22428 62188 22484
rect 62132 22372 62188 22428
rect 64652 22372 64708 22540
rect 65762 22428 65772 22484
rect 65828 22428 67004 22484
rect 67060 22428 67070 22484
rect 69458 22428 69468 22484
rect 69524 22428 70476 22484
rect 70532 22428 70542 22484
rect 4946 22316 4956 22372
rect 5012 22316 5740 22372
rect 5796 22316 5806 22372
rect 15922 22316 15932 22372
rect 15988 22316 22092 22372
rect 22148 22316 30660 22372
rect 39890 22316 39900 22372
rect 39956 22316 40684 22372
rect 40740 22316 40750 22372
rect 42130 22316 42140 22372
rect 42196 22316 43260 22372
rect 43316 22316 50092 22372
rect 50148 22316 50158 22372
rect 50642 22316 50652 22372
rect 50708 22316 59500 22372
rect 59556 22316 59566 22372
rect 62132 22316 63084 22372
rect 63140 22316 63150 22372
rect 64652 22316 73052 22372
rect 73108 22316 73118 22372
rect 30604 22260 30660 22316
rect 3154 22204 3164 22260
rect 3220 22204 3836 22260
rect 3892 22204 3902 22260
rect 6290 22204 6300 22260
rect 6356 22204 16268 22260
rect 16324 22204 17052 22260
rect 17108 22204 17118 22260
rect 18172 22204 22036 22260
rect 26562 22204 26572 22260
rect 26628 22204 29988 22260
rect 30594 22204 30604 22260
rect 30660 22204 31052 22260
rect 31108 22204 31118 22260
rect 34626 22204 34636 22260
rect 34692 22204 36988 22260
rect 37044 22204 37054 22260
rect 39442 22204 39452 22260
rect 39508 22204 39788 22260
rect 39844 22204 39854 22260
rect 46732 22204 50204 22260
rect 50260 22204 59612 22260
rect 59668 22204 60060 22260
rect 60116 22204 60126 22260
rect 69346 22204 69356 22260
rect 69412 22204 70700 22260
rect 70756 22204 70766 22260
rect 71586 22204 71596 22260
rect 71652 22204 71932 22260
rect 71988 22204 71998 22260
rect 18172 22148 18228 22204
rect 21980 22148 22036 22204
rect 29932 22148 29988 22204
rect 46732 22148 46788 22204
rect 11330 22092 11340 22148
rect 11396 22092 13468 22148
rect 13524 22092 13534 22148
rect 13794 22092 13804 22148
rect 13860 22092 14252 22148
rect 14308 22092 18228 22148
rect 18386 22092 18396 22148
rect 18452 22092 18462 22148
rect 21970 22092 21980 22148
rect 22036 22092 22046 22148
rect 26002 22092 26012 22148
rect 26068 22092 28140 22148
rect 28196 22092 28206 22148
rect 29922 22092 29932 22148
rect 29988 22092 43708 22148
rect 43764 22092 43774 22148
rect 44930 22092 44940 22148
rect 44996 22092 46732 22148
rect 46788 22092 46798 22148
rect 50372 22092 62300 22148
rect 62356 22092 62366 22148
rect 69458 22092 69468 22148
rect 69524 22092 69534 22148
rect 69906 22092 69916 22148
rect 69972 22092 70364 22148
rect 70420 22092 70430 22148
rect 73826 22092 73836 22148
rect 73892 22092 74172 22148
rect 74228 22092 74238 22148
rect 18396 22036 18452 22092
rect 14914 21980 14924 22036
rect 14980 21980 18452 22036
rect 23538 21980 23548 22036
rect 23604 21980 24108 22036
rect 24164 21980 25004 22036
rect 25060 21980 31276 22036
rect 31332 21980 31342 22036
rect 35970 21980 35980 22036
rect 36036 21980 36540 22036
rect 36596 21980 36606 22036
rect 20522 21924 20532 21980
rect 20588 21924 20636 21980
rect 20692 21924 20740 21980
rect 20796 21924 20806 21980
rect 39842 21924 39852 21980
rect 39908 21924 39956 21980
rect 40012 21924 40060 21980
rect 40116 21924 40126 21980
rect 50372 21924 50428 22092
rect 69468 22036 69524 22092
rect 51314 21980 51324 22036
rect 51380 21980 51996 22036
rect 52052 21980 52062 22036
rect 56578 21980 56588 22036
rect 56644 21980 58268 22036
rect 58324 21980 58334 22036
rect 69468 21980 72828 22036
rect 72884 21980 74844 22036
rect 74900 21980 74910 22036
rect 59162 21924 59172 21980
rect 59228 21924 59276 21980
rect 59332 21924 59380 21980
rect 59436 21924 59446 21980
rect 78482 21924 78492 21980
rect 78548 21924 78596 21980
rect 78652 21924 78700 21980
rect 78756 21924 78766 21980
rect 14018 21868 14028 21924
rect 14084 21868 15484 21924
rect 15540 21868 15550 21924
rect 16818 21868 16828 21924
rect 16884 21868 18396 21924
rect 18452 21868 18462 21924
rect 22754 21868 22764 21924
rect 22820 21868 23884 21924
rect 23940 21868 23950 21924
rect 25666 21868 25676 21924
rect 25732 21868 26796 21924
rect 26852 21868 28364 21924
rect 28420 21868 28430 21924
rect 30930 21868 30940 21924
rect 30996 21868 31948 21924
rect 32004 21868 32014 21924
rect 40450 21868 40460 21924
rect 40516 21868 41916 21924
rect 41972 21868 50428 21924
rect 51650 21868 51660 21924
rect 51716 21868 52892 21924
rect 52948 21868 52958 21924
rect 70690 21868 70700 21924
rect 70756 21868 71036 21924
rect 71092 21868 71102 21924
rect 74050 21868 74060 21924
rect 74116 21868 75180 21924
rect 75236 21868 75246 21924
rect 4050 21756 4060 21812
rect 4116 21756 4956 21812
rect 5012 21756 5022 21812
rect 6178 21756 6188 21812
rect 6244 21756 10556 21812
rect 10612 21756 10622 21812
rect 11778 21756 11788 21812
rect 11844 21756 12684 21812
rect 12740 21756 13468 21812
rect 13524 21756 14140 21812
rect 14196 21756 14206 21812
rect 14466 21756 14476 21812
rect 14532 21756 16604 21812
rect 16660 21756 16670 21812
rect 18498 21756 18508 21812
rect 18564 21756 19292 21812
rect 19348 21756 19358 21812
rect 22978 21756 22988 21812
rect 23044 21756 24108 21812
rect 24164 21756 24174 21812
rect 25890 21756 25900 21812
rect 25956 21756 27020 21812
rect 27076 21756 27086 21812
rect 27234 21756 27244 21812
rect 27300 21756 27580 21812
rect 27636 21756 29596 21812
rect 29652 21756 29662 21812
rect 29922 21756 29932 21812
rect 29988 21756 33516 21812
rect 33572 21756 33582 21812
rect 35298 21756 35308 21812
rect 35364 21756 36204 21812
rect 36260 21756 36270 21812
rect 38770 21756 38780 21812
rect 38836 21756 40348 21812
rect 40404 21756 40414 21812
rect 40674 21756 40684 21812
rect 40740 21756 41804 21812
rect 41860 21756 42364 21812
rect 42420 21756 42430 21812
rect 49746 21756 49756 21812
rect 49812 21756 50316 21812
rect 50372 21756 50382 21812
rect 50866 21756 50876 21812
rect 50932 21756 51436 21812
rect 51492 21756 52332 21812
rect 52388 21756 52398 21812
rect 57586 21756 57596 21812
rect 57652 21756 59052 21812
rect 59108 21756 59118 21812
rect 59826 21756 59836 21812
rect 59892 21756 60508 21812
rect 60564 21756 60574 21812
rect 66210 21756 66220 21812
rect 66276 21756 66892 21812
rect 66948 21756 66958 21812
rect 68674 21756 68684 21812
rect 68740 21756 72604 21812
rect 72660 21756 72670 21812
rect 73490 21756 73500 21812
rect 73556 21756 73566 21812
rect 74722 21756 74732 21812
rect 74788 21756 76300 21812
rect 76356 21756 76366 21812
rect 73500 21700 73556 21756
rect 4162 21644 4172 21700
rect 4228 21644 9996 21700
rect 10052 21644 10062 21700
rect 10434 21644 10444 21700
rect 10500 21644 11564 21700
rect 11620 21644 11630 21700
rect 15586 21644 15596 21700
rect 15652 21644 16940 21700
rect 16996 21644 17006 21700
rect 17378 21644 17388 21700
rect 17444 21644 18732 21700
rect 18788 21644 20300 21700
rect 20356 21644 20366 21700
rect 24322 21644 24332 21700
rect 24388 21644 31164 21700
rect 31220 21644 31230 21700
rect 32722 21644 32732 21700
rect 32788 21644 37380 21700
rect 38434 21644 38444 21700
rect 38500 21644 41356 21700
rect 41412 21644 41422 21700
rect 51314 21644 51324 21700
rect 51380 21644 51772 21700
rect 51828 21644 51838 21700
rect 67106 21644 67116 21700
rect 67172 21644 67676 21700
rect 67732 21644 67742 21700
rect 71362 21644 71372 21700
rect 71428 21644 71438 21700
rect 73500 21644 73724 21700
rect 73780 21644 73790 21700
rect 75842 21644 75852 21700
rect 75908 21644 77868 21700
rect 77924 21644 77934 21700
rect 37324 21588 37380 21644
rect 9426 21532 9436 21588
rect 9492 21532 9884 21588
rect 9940 21532 10332 21588
rect 10388 21532 10398 21588
rect 11106 21532 11116 21588
rect 11172 21532 12012 21588
rect 12068 21532 12078 21588
rect 15922 21532 15932 21588
rect 15988 21532 17276 21588
rect 17332 21532 17342 21588
rect 19282 21532 19292 21588
rect 19348 21532 21420 21588
rect 21476 21532 21486 21588
rect 23426 21532 23436 21588
rect 23492 21532 23772 21588
rect 23828 21532 23838 21588
rect 24658 21532 24668 21588
rect 24724 21532 26124 21588
rect 26180 21532 26190 21588
rect 26450 21532 26460 21588
rect 26516 21532 26526 21588
rect 26852 21532 27804 21588
rect 27860 21532 29372 21588
rect 29428 21532 29438 21588
rect 29586 21532 29596 21588
rect 29652 21532 29662 21588
rect 29810 21532 29820 21588
rect 29876 21532 30380 21588
rect 30436 21532 31612 21588
rect 31668 21532 31678 21588
rect 36418 21532 36428 21588
rect 36484 21532 37100 21588
rect 37156 21532 37166 21588
rect 37324 21532 42812 21588
rect 42868 21532 43372 21588
rect 43428 21532 43438 21588
rect 43922 21532 43932 21588
rect 43988 21532 44828 21588
rect 44884 21532 45612 21588
rect 45668 21532 45678 21588
rect 47506 21532 47516 21588
rect 47572 21532 48860 21588
rect 48916 21532 49868 21588
rect 49924 21532 49934 21588
rect 51538 21532 51548 21588
rect 51604 21532 51884 21588
rect 51940 21532 51950 21588
rect 56802 21532 56812 21588
rect 56868 21532 58380 21588
rect 58436 21532 58446 21588
rect 65314 21532 65324 21588
rect 65380 21532 69692 21588
rect 69748 21532 69758 21588
rect 11116 21476 11172 21532
rect 8978 21420 8988 21476
rect 9044 21420 11172 21476
rect 11442 21420 11452 21476
rect 11508 21420 19404 21476
rect 19460 21420 19470 21476
rect 22418 21420 22428 21476
rect 22484 21420 23884 21476
rect 23940 21420 23950 21476
rect 24668 21420 25564 21476
rect 25620 21420 25788 21476
rect 25844 21420 25854 21476
rect 10546 21308 10556 21364
rect 10612 21308 11900 21364
rect 11956 21308 11966 21364
rect 14354 21308 14364 21364
rect 14420 21308 18284 21364
rect 18340 21308 18350 21364
rect 24668 21252 24724 21420
rect 26460 21364 26516 21532
rect 26852 21364 26908 21532
rect 29596 21476 29652 21532
rect 43372 21476 43428 21532
rect 71372 21476 71428 21644
rect 71698 21532 71708 21588
rect 71764 21532 72940 21588
rect 72996 21532 74844 21588
rect 74900 21532 74910 21588
rect 28578 21420 28588 21476
rect 28644 21420 29148 21476
rect 29204 21420 29214 21476
rect 29596 21420 33180 21476
rect 33236 21420 33246 21476
rect 34290 21420 34300 21476
rect 34356 21420 36316 21476
rect 36372 21420 36988 21476
rect 37044 21420 37054 21476
rect 38882 21420 38892 21476
rect 38948 21420 39228 21476
rect 39284 21420 40124 21476
rect 40180 21420 40190 21476
rect 43372 21420 44492 21476
rect 44548 21420 45500 21476
rect 45556 21420 45566 21476
rect 47170 21420 47180 21476
rect 47236 21420 48636 21476
rect 48692 21420 48702 21476
rect 59938 21420 59948 21476
rect 60004 21420 60620 21476
rect 60676 21420 60686 21476
rect 66658 21420 66668 21476
rect 66724 21420 67228 21476
rect 67284 21420 69580 21476
rect 69636 21420 69646 21476
rect 71372 21420 72492 21476
rect 72548 21420 73948 21476
rect 74004 21420 74014 21476
rect 26460 21308 26908 21364
rect 29586 21308 29596 21364
rect 29652 21308 30268 21364
rect 30324 21308 30334 21364
rect 31154 21308 31164 21364
rect 31220 21308 32284 21364
rect 32340 21308 44268 21364
rect 44324 21308 45388 21364
rect 45444 21308 45454 21364
rect 45938 21308 45948 21364
rect 46004 21308 60508 21364
rect 60564 21308 60574 21364
rect 70578 21308 70588 21364
rect 70644 21308 71148 21364
rect 71204 21308 71214 21364
rect 13570 21196 13580 21252
rect 13636 21196 14476 21252
rect 14532 21196 14542 21252
rect 16370 21196 16380 21252
rect 16436 21196 16716 21252
rect 16772 21196 16782 21252
rect 20178 21196 20188 21252
rect 20244 21196 24668 21252
rect 24724 21196 24734 21252
rect 36194 21196 36204 21252
rect 36260 21196 45780 21252
rect 0 21140 800 21168
rect 10862 21140 10872 21196
rect 10928 21140 10976 21196
rect 11032 21140 11080 21196
rect 11136 21140 11146 21196
rect 30182 21140 30192 21196
rect 30248 21140 30296 21196
rect 30352 21140 30400 21196
rect 30456 21140 30466 21196
rect 0 21084 2772 21140
rect 12114 21084 12124 21140
rect 12180 21084 17836 21140
rect 17892 21084 18620 21140
rect 18676 21084 19628 21140
rect 19684 21084 19694 21140
rect 38612 21084 44940 21140
rect 44996 21084 45500 21140
rect 45556 21084 45566 21140
rect 0 21056 800 21084
rect 2716 21028 2772 21084
rect 38612 21028 38668 21084
rect 45724 21028 45780 21196
rect 49502 21140 49512 21196
rect 49568 21140 49616 21196
rect 49672 21140 49720 21196
rect 49776 21140 49786 21196
rect 68822 21140 68832 21196
rect 68888 21140 68936 21196
rect 68992 21140 69040 21196
rect 69096 21140 69106 21196
rect 79200 21140 80000 21168
rect 70690 21084 70700 21140
rect 70756 21084 72716 21140
rect 72772 21084 72782 21140
rect 77970 21084 77980 21140
rect 78036 21084 80000 21140
rect 79200 21056 80000 21084
rect 2706 20972 2716 21028
rect 2772 20972 2782 21028
rect 20626 20972 20636 21028
rect 20692 20972 21084 21028
rect 21140 20972 25228 21028
rect 25284 20972 25294 21028
rect 26852 20972 38668 21028
rect 39330 20972 39340 21028
rect 39396 20972 42140 21028
rect 42196 20972 42700 21028
rect 42756 20972 42766 21028
rect 45724 20972 59724 21028
rect 59780 20972 59790 21028
rect 26852 20916 26908 20972
rect 4946 20860 4956 20916
rect 5012 20860 11676 20916
rect 11732 20860 11742 20916
rect 16930 20860 16940 20916
rect 16996 20860 17836 20916
rect 17892 20860 21812 20916
rect 23762 20860 23772 20916
rect 23828 20860 26908 20916
rect 31154 20860 31164 20916
rect 31220 20860 32732 20916
rect 32788 20860 32798 20916
rect 36418 20860 36428 20916
rect 36484 20860 40236 20916
rect 40292 20860 40302 20916
rect 44156 20860 49084 20916
rect 49140 20860 49150 20916
rect 61058 20860 61068 20916
rect 61124 20860 70028 20916
rect 70084 20860 70588 20916
rect 70644 20860 70812 20916
rect 70868 20860 71932 20916
rect 71988 20860 71998 20916
rect 11004 20804 11060 20860
rect 5730 20748 5740 20804
rect 5796 20748 6916 20804
rect 9986 20748 9996 20804
rect 10052 20748 10444 20804
rect 10500 20748 10510 20804
rect 10994 20748 11004 20804
rect 11060 20748 11070 20804
rect 6860 20692 6916 20748
rect 4946 20636 4956 20692
rect 5012 20636 5852 20692
rect 5908 20636 5918 20692
rect 6850 20636 6860 20692
rect 6916 20636 11228 20692
rect 11284 20636 11788 20692
rect 11844 20636 11854 20692
rect 16370 20636 16380 20692
rect 16436 20636 16716 20692
rect 16772 20636 16782 20692
rect 10098 20524 10108 20580
rect 10164 20524 10174 20580
rect 11666 20524 11676 20580
rect 11732 20524 15708 20580
rect 15764 20524 15774 20580
rect 10108 20132 10164 20524
rect 10770 20412 10780 20468
rect 10836 20412 12236 20468
rect 12292 20412 12302 20468
rect 16940 20356 16996 20860
rect 18274 20748 18284 20804
rect 18340 20748 19964 20804
rect 20020 20748 20030 20804
rect 20850 20748 20860 20804
rect 20916 20748 21532 20804
rect 21588 20748 21598 20804
rect 21756 20692 21812 20860
rect 44156 20804 44212 20860
rect 26226 20748 26236 20804
rect 26292 20748 26908 20804
rect 29810 20748 29820 20804
rect 29876 20748 30828 20804
rect 30884 20748 31388 20804
rect 31444 20748 44212 20804
rect 47842 20748 47852 20804
rect 47908 20748 48748 20804
rect 48804 20748 48814 20804
rect 49970 20748 49980 20804
rect 50036 20748 50316 20804
rect 50372 20748 50382 20804
rect 60732 20748 62412 20804
rect 62468 20748 62478 20804
rect 62850 20748 62860 20804
rect 62916 20748 67004 20804
rect 67060 20748 67070 20804
rect 73714 20748 73724 20804
rect 73780 20748 75068 20804
rect 75124 20748 75134 20804
rect 26852 20692 26908 20748
rect 60732 20692 60788 20748
rect 62860 20692 62916 20748
rect 17266 20636 17276 20692
rect 17332 20636 21308 20692
rect 21364 20636 21374 20692
rect 21746 20636 21756 20692
rect 21812 20636 22092 20692
rect 22148 20636 26180 20692
rect 26852 20636 28140 20692
rect 28196 20636 28206 20692
rect 33282 20636 33292 20692
rect 33348 20636 35420 20692
rect 35476 20636 36428 20692
rect 36484 20636 36494 20692
rect 38612 20636 40124 20692
rect 40180 20636 40190 20692
rect 48626 20636 48636 20692
rect 48692 20636 50204 20692
rect 50260 20636 50988 20692
rect 51044 20636 51772 20692
rect 51828 20636 51838 20692
rect 56802 20636 56812 20692
rect 56868 20636 60732 20692
rect 60788 20636 60798 20692
rect 60956 20636 62916 20692
rect 64306 20636 64316 20692
rect 64372 20636 65100 20692
rect 65156 20636 65166 20692
rect 71474 20636 71484 20692
rect 71540 20636 72828 20692
rect 72884 20636 72894 20692
rect 21308 20580 21364 20636
rect 26124 20580 26180 20636
rect 38612 20580 38668 20636
rect 60956 20580 61012 20636
rect 17154 20524 17164 20580
rect 17220 20524 18284 20580
rect 18340 20524 18350 20580
rect 18498 20524 18508 20580
rect 18564 20524 18956 20580
rect 19012 20524 19022 20580
rect 19394 20524 19404 20580
rect 19460 20524 19740 20580
rect 19796 20524 19806 20580
rect 21308 20524 25004 20580
rect 25060 20524 25070 20580
rect 25890 20524 25900 20580
rect 25956 20524 25966 20580
rect 26124 20524 27356 20580
rect 27412 20524 27422 20580
rect 29250 20524 29260 20580
rect 29316 20524 29988 20580
rect 30258 20524 30268 20580
rect 30324 20524 31164 20580
rect 31220 20524 31230 20580
rect 36306 20524 36316 20580
rect 36372 20524 38668 20580
rect 43026 20524 43036 20580
rect 43092 20524 43932 20580
rect 43988 20524 43998 20580
rect 45154 20524 45164 20580
rect 45220 20524 45948 20580
rect 46004 20524 46014 20580
rect 52098 20524 52108 20580
rect 52164 20524 52780 20580
rect 52836 20524 52846 20580
rect 57820 20524 60956 20580
rect 61012 20524 61022 20580
rect 61618 20524 61628 20580
rect 61684 20524 63084 20580
rect 63140 20524 63150 20580
rect 25900 20468 25956 20524
rect 29932 20468 29988 20524
rect 57820 20468 57876 20524
rect 18722 20412 18732 20468
rect 18788 20412 19068 20468
rect 19124 20412 19134 20468
rect 25900 20412 28700 20468
rect 28756 20412 29708 20468
rect 29764 20412 29774 20468
rect 29932 20412 38780 20468
rect 38836 20412 38846 20468
rect 48178 20412 48188 20468
rect 48244 20412 57876 20468
rect 60498 20412 60508 20468
rect 60564 20412 62076 20468
rect 62132 20412 62142 20468
rect 20522 20356 20532 20412
rect 20588 20356 20636 20412
rect 20692 20356 20740 20412
rect 20796 20356 20806 20412
rect 39842 20356 39852 20412
rect 39908 20356 39956 20412
rect 40012 20356 40060 20412
rect 40116 20356 40126 20412
rect 59162 20356 59172 20412
rect 59228 20356 59276 20412
rect 59332 20356 59380 20412
rect 59436 20356 59446 20412
rect 78482 20356 78492 20412
rect 78548 20356 78596 20412
rect 78652 20356 78700 20412
rect 78756 20356 78766 20412
rect 16594 20300 16604 20356
rect 16660 20300 16996 20356
rect 22530 20300 22540 20356
rect 22596 20300 23548 20356
rect 23604 20300 24668 20356
rect 24724 20300 24734 20356
rect 30146 20300 30156 20356
rect 30212 20300 37548 20356
rect 37604 20300 37614 20356
rect 52658 20300 52668 20356
rect 52724 20300 58604 20356
rect 58660 20300 58670 20356
rect 59714 20300 59724 20356
rect 59780 20300 62188 20356
rect 63298 20300 63308 20356
rect 63364 20300 68460 20356
rect 68516 20300 69020 20356
rect 69076 20300 69086 20356
rect 62132 20244 62188 20300
rect 10322 20188 10332 20244
rect 10388 20188 10668 20244
rect 10724 20188 10734 20244
rect 12562 20188 12572 20244
rect 12628 20188 29820 20244
rect 29876 20188 29886 20244
rect 32834 20188 32844 20244
rect 32900 20188 34076 20244
rect 34132 20188 34142 20244
rect 48850 20188 48860 20244
rect 48916 20188 49420 20244
rect 49476 20188 49486 20244
rect 54786 20188 54796 20244
rect 54852 20188 56700 20244
rect 56756 20188 56766 20244
rect 60610 20188 60620 20244
rect 60676 20188 61628 20244
rect 61684 20188 61694 20244
rect 62132 20188 75292 20244
rect 75348 20188 75740 20244
rect 75796 20188 75806 20244
rect 7298 20076 7308 20132
rect 7364 20076 8540 20132
rect 8596 20076 8606 20132
rect 10108 20076 11900 20132
rect 11956 20076 11966 20132
rect 15092 20076 26908 20132
rect 26964 20076 26974 20132
rect 27906 20076 27916 20132
rect 27972 20076 30940 20132
rect 30996 20076 31006 20132
rect 32162 20076 32172 20132
rect 32228 20076 32508 20132
rect 32564 20076 33404 20132
rect 33460 20076 33964 20132
rect 34020 20076 34524 20132
rect 34580 20076 34590 20132
rect 40450 20076 40460 20132
rect 40516 20076 41356 20132
rect 41412 20076 42476 20132
rect 42532 20076 42542 20132
rect 42690 20076 42700 20132
rect 42756 20076 43260 20132
rect 43316 20076 43326 20132
rect 58258 20076 58268 20132
rect 58324 20076 59164 20132
rect 59220 20076 59230 20132
rect 61170 20076 61180 20132
rect 61236 20076 62188 20132
rect 63746 20076 63756 20132
rect 63812 20076 64540 20132
rect 64596 20076 64606 20132
rect 67106 20076 67116 20132
rect 67172 20076 69356 20132
rect 69412 20076 69422 20132
rect 15092 20020 15148 20076
rect 8082 19964 8092 20020
rect 8148 19964 9660 20020
rect 9716 19964 9726 20020
rect 10098 19964 10108 20020
rect 10164 19964 11676 20020
rect 11732 19964 11742 20020
rect 11900 19964 15148 20020
rect 16370 19964 16380 20020
rect 16436 19964 17556 20020
rect 23090 19964 23100 20020
rect 23156 19964 24052 20020
rect 27122 19964 27132 20020
rect 27188 19964 27468 20020
rect 27524 19964 27804 20020
rect 27860 19964 29372 20020
rect 29428 19964 29438 20020
rect 49858 19964 49868 20020
rect 49924 19964 54348 20020
rect 54404 19964 54414 20020
rect 59378 19964 59388 20020
rect 59444 19964 60844 20020
rect 60900 19964 60910 20020
rect 62132 19964 62188 20076
rect 62244 19964 62254 20020
rect 64866 19964 64876 20020
rect 64932 19964 67228 20020
rect 67284 19964 67294 20020
rect 69570 19964 69580 20020
rect 69636 19964 71596 20020
rect 71652 19964 71662 20020
rect 11900 19796 11956 19964
rect 17500 19908 17556 19964
rect 23996 19908 24052 19964
rect 64876 19908 64932 19964
rect 15036 19852 16268 19908
rect 16324 19852 17164 19908
rect 17220 19852 17230 19908
rect 17490 19852 17500 19908
rect 17556 19852 19516 19908
rect 19572 19852 19582 19908
rect 20178 19852 20188 19908
rect 20244 19852 21868 19908
rect 21924 19852 23548 19908
rect 23604 19852 23614 19908
rect 23986 19852 23996 19908
rect 24052 19852 24062 19908
rect 25218 19852 25228 19908
rect 25284 19852 27972 19908
rect 28130 19852 28140 19908
rect 28196 19852 29036 19908
rect 29092 19852 29932 19908
rect 29988 19852 29998 19908
rect 36754 19852 36764 19908
rect 36820 19852 47068 19908
rect 47124 19852 47134 19908
rect 50306 19852 50316 19908
rect 50372 19852 50428 19908
rect 50484 19852 50494 19908
rect 52770 19852 52780 19908
rect 52836 19852 53228 19908
rect 53284 19852 56028 19908
rect 56084 19852 56094 19908
rect 58034 19852 58044 19908
rect 58100 19852 64932 19908
rect 68674 19852 68684 19908
rect 68740 19852 70476 19908
rect 70532 19852 70542 19908
rect 15036 19796 15092 19852
rect 27916 19796 27972 19852
rect 4386 19740 4396 19796
rect 4452 19740 11956 19796
rect 13906 19740 13916 19796
rect 13972 19740 15092 19796
rect 16146 19740 16156 19796
rect 16212 19740 17276 19796
rect 17332 19740 17342 19796
rect 23314 19740 23324 19796
rect 23380 19740 27244 19796
rect 27300 19740 27310 19796
rect 27916 19740 33572 19796
rect 34626 19740 34636 19796
rect 34692 19740 35420 19796
rect 35476 19740 35486 19796
rect 42018 19740 42028 19796
rect 42084 19740 43708 19796
rect 43764 19740 61068 19796
rect 61124 19740 61852 19796
rect 61908 19740 61918 19796
rect 62290 19740 62300 19796
rect 62356 19740 63196 19796
rect 63252 19740 65436 19796
rect 65492 19740 65502 19796
rect 69010 19740 69020 19796
rect 69076 19740 70812 19796
rect 70868 19740 70878 19796
rect 33516 19684 33572 19740
rect 15810 19628 15820 19684
rect 15876 19628 16604 19684
rect 16660 19628 16670 19684
rect 21970 19628 21980 19684
rect 22036 19628 30100 19684
rect 33516 19628 35308 19684
rect 35364 19628 35374 19684
rect 50372 19628 63868 19684
rect 63924 19628 64988 19684
rect 65044 19628 65054 19684
rect 10862 19572 10872 19628
rect 10928 19572 10976 19628
rect 11032 19572 11080 19628
rect 11136 19572 11146 19628
rect 21858 19516 21868 19572
rect 21924 19516 22316 19572
rect 22372 19516 22382 19572
rect 30044 19460 30100 19628
rect 30182 19572 30192 19628
rect 30248 19572 30296 19628
rect 30352 19572 30400 19628
rect 30456 19572 30466 19628
rect 49502 19572 49512 19628
rect 49568 19572 49616 19628
rect 49672 19572 49720 19628
rect 49776 19572 49786 19628
rect 30706 19516 30716 19572
rect 30772 19516 41132 19572
rect 41188 19516 41198 19572
rect 42354 19516 42364 19572
rect 42420 19516 44492 19572
rect 44548 19516 44558 19572
rect 50372 19460 50428 19628
rect 68822 19572 68832 19628
rect 68888 19572 68936 19628
rect 68992 19572 69040 19628
rect 69096 19572 69106 19628
rect 55010 19516 55020 19572
rect 55076 19516 55468 19572
rect 55524 19516 62300 19572
rect 62356 19516 62366 19572
rect 10546 19404 10556 19460
rect 10612 19404 14812 19460
rect 14868 19404 14878 19460
rect 15026 19404 15036 19460
rect 15092 19404 23100 19460
rect 23156 19404 23166 19460
rect 23986 19404 23996 19460
rect 24052 19404 24892 19460
rect 24948 19404 26236 19460
rect 26292 19404 26302 19460
rect 27010 19404 27020 19460
rect 27076 19404 28588 19460
rect 28644 19404 28654 19460
rect 30044 19404 33628 19460
rect 33684 19404 33694 19460
rect 38210 19404 38220 19460
rect 38276 19404 40572 19460
rect 40628 19404 40638 19460
rect 46722 19404 46732 19460
rect 46788 19404 50428 19460
rect 61842 19404 61852 19460
rect 61908 19404 76188 19460
rect 76244 19404 76254 19460
rect 5394 19292 5404 19348
rect 5460 19292 40460 19348
rect 40516 19292 40526 19348
rect 41682 19292 41692 19348
rect 41748 19292 50316 19348
rect 50372 19292 50382 19348
rect 69682 19292 69692 19348
rect 69748 19292 70252 19348
rect 70308 19292 70318 19348
rect 74946 19292 74956 19348
rect 75012 19292 76860 19348
rect 76916 19292 78092 19348
rect 78148 19292 78158 19348
rect 12114 19180 12124 19236
rect 12180 19180 12684 19236
rect 12740 19180 12750 19236
rect 18386 19180 18396 19236
rect 18452 19180 18620 19236
rect 18676 19180 18686 19236
rect 26114 19180 26124 19236
rect 26180 19180 26572 19236
rect 26628 19180 27132 19236
rect 27188 19180 27356 19236
rect 27412 19180 27916 19236
rect 27972 19180 27982 19236
rect 28578 19180 28588 19236
rect 28644 19180 29036 19236
rect 29092 19180 29102 19236
rect 29698 19180 29708 19236
rect 29764 19180 32396 19236
rect 32452 19180 33180 19236
rect 33236 19180 33246 19236
rect 36418 19180 36428 19236
rect 36484 19180 39452 19236
rect 39508 19180 42252 19236
rect 42308 19180 42318 19236
rect 50372 19180 57820 19236
rect 57876 19180 59276 19236
rect 59332 19180 60172 19236
rect 60228 19180 60238 19236
rect 66434 19180 66444 19236
rect 66500 19180 71820 19236
rect 71876 19180 71886 19236
rect 10098 19068 10108 19124
rect 10164 19068 10892 19124
rect 10948 19068 11340 19124
rect 11396 19068 11406 19124
rect 14802 19068 14812 19124
rect 14868 19068 16828 19124
rect 16884 19068 16894 19124
rect 17826 19068 17836 19124
rect 17892 19068 18284 19124
rect 18340 19068 18350 19124
rect 21634 19068 21644 19124
rect 21700 19068 21980 19124
rect 22036 19068 22046 19124
rect 28018 19068 28028 19124
rect 28084 19068 30268 19124
rect 30324 19068 30334 19124
rect 30930 19068 30940 19124
rect 30996 19068 39116 19124
rect 39172 19068 43932 19124
rect 43988 19068 44940 19124
rect 44996 19068 45006 19124
rect 50372 19012 50428 19180
rect 52994 19068 53004 19124
rect 53060 19068 54124 19124
rect 54180 19068 59388 19124
rect 59444 19068 59454 19124
rect 68898 19068 68908 19124
rect 68964 19068 69804 19124
rect 69860 19068 69870 19124
rect 70252 19012 70308 19180
rect 72594 19068 72604 19124
rect 72660 19068 73276 19124
rect 73332 19068 73342 19124
rect 75618 19068 75628 19124
rect 75684 19068 77644 19124
rect 77700 19068 77710 19124
rect 14354 18956 14364 19012
rect 14420 18956 16044 19012
rect 16100 18956 20188 19012
rect 20244 18956 20254 19012
rect 21858 18956 21868 19012
rect 21924 18956 22988 19012
rect 23044 18956 23436 19012
rect 23492 18956 23502 19012
rect 25218 18956 25228 19012
rect 25284 18956 25676 19012
rect 25732 18956 25742 19012
rect 29698 18956 29708 19012
rect 29764 18956 30716 19012
rect 30772 18956 30782 19012
rect 38098 18956 38108 19012
rect 38164 18956 40684 19012
rect 40740 18956 40750 19012
rect 41570 18956 41580 19012
rect 41636 18956 42476 19012
rect 42532 18956 42542 19012
rect 47506 18956 47516 19012
rect 47572 18956 49196 19012
rect 49252 18956 50428 19012
rect 54796 18956 62188 19012
rect 65202 18956 65212 19012
rect 65268 18956 69916 19012
rect 69972 18956 69982 19012
rect 70242 18956 70252 19012
rect 70308 18956 70318 19012
rect 75282 18956 75292 19012
rect 75348 18956 77196 19012
rect 77252 18956 77262 19012
rect 54796 18900 54852 18956
rect 11218 18844 11228 18900
rect 11284 18844 11294 18900
rect 16370 18844 16380 18900
rect 16436 18844 17388 18900
rect 17444 18844 17454 18900
rect 17826 18844 17836 18900
rect 17892 18844 18396 18900
rect 18452 18844 18462 18900
rect 21970 18844 21980 18900
rect 22036 18844 24220 18900
rect 24276 18844 28028 18900
rect 28084 18844 28094 18900
rect 28252 18844 37716 18900
rect 49410 18844 49420 18900
rect 49476 18844 54852 18900
rect 0 18676 800 18704
rect 0 18620 1932 18676
rect 1988 18620 1998 18676
rect 0 18592 800 18620
rect 11228 18564 11284 18844
rect 20522 18788 20532 18844
rect 20588 18788 20636 18844
rect 20692 18788 20740 18844
rect 20796 18788 20806 18844
rect 28252 18788 28308 18844
rect 37660 18788 37716 18844
rect 39842 18788 39852 18844
rect 39908 18788 39956 18844
rect 40012 18788 40060 18844
rect 40116 18788 40126 18844
rect 59162 18788 59172 18844
rect 59228 18788 59276 18844
rect 59332 18788 59380 18844
rect 59436 18788 59446 18844
rect 62132 18788 62188 18956
rect 66994 18844 67004 18900
rect 67060 18844 67564 18900
rect 67620 18844 70588 18900
rect 70644 18844 70654 18900
rect 78482 18788 78492 18844
rect 78548 18788 78596 18844
rect 78652 18788 78700 18844
rect 78756 18788 78766 18844
rect 15922 18732 15932 18788
rect 15988 18732 20356 18788
rect 23090 18732 23100 18788
rect 23156 18732 23436 18788
rect 23492 18732 23502 18788
rect 27234 18732 27244 18788
rect 27300 18732 28308 18788
rect 36866 18732 36876 18788
rect 36932 18732 37436 18788
rect 37492 18732 37502 18788
rect 37650 18732 37660 18788
rect 37716 18732 37726 18788
rect 62132 18732 72492 18788
rect 72548 18732 72558 18788
rect 13010 18620 13020 18676
rect 13076 18620 14252 18676
rect 14308 18620 14318 18676
rect 16706 18620 16716 18676
rect 16772 18620 18956 18676
rect 19012 18620 19022 18676
rect 20300 18564 20356 18732
rect 79200 18676 80000 18704
rect 23762 18620 23772 18676
rect 23828 18620 26124 18676
rect 26180 18620 26190 18676
rect 33506 18620 33516 18676
rect 33572 18620 50204 18676
rect 50260 18620 50270 18676
rect 55122 18620 55132 18676
rect 55188 18620 57036 18676
rect 57092 18620 58604 18676
rect 58660 18620 58940 18676
rect 58996 18620 59006 18676
rect 70802 18620 70812 18676
rect 70868 18620 71372 18676
rect 71428 18620 71820 18676
rect 71876 18620 71886 18676
rect 73892 18564 73948 18676
rect 74004 18620 74014 18676
rect 75058 18620 75068 18676
rect 75124 18620 80000 18676
rect 79200 18592 80000 18620
rect 11228 18508 14700 18564
rect 14756 18508 14766 18564
rect 16818 18508 16828 18564
rect 16884 18508 19068 18564
rect 19124 18508 19134 18564
rect 20300 18508 21756 18564
rect 21812 18508 21822 18564
rect 34962 18508 34972 18564
rect 35028 18508 37324 18564
rect 37380 18508 37390 18564
rect 48962 18508 48972 18564
rect 49028 18508 54236 18564
rect 54292 18508 54302 18564
rect 54898 18508 54908 18564
rect 54964 18508 55468 18564
rect 55524 18508 55534 18564
rect 59052 18508 65660 18564
rect 65716 18508 66780 18564
rect 66836 18508 66846 18564
rect 70578 18508 70588 18564
rect 70644 18508 73948 18564
rect 5730 18396 5740 18452
rect 5796 18396 6412 18452
rect 6468 18396 7532 18452
rect 7588 18396 7598 18452
rect 12338 18396 12348 18452
rect 12404 18396 13132 18452
rect 13188 18396 13198 18452
rect 18610 18396 18620 18452
rect 18676 18396 18956 18452
rect 19012 18396 19022 18452
rect 20066 18396 20076 18452
rect 20132 18396 20860 18452
rect 20916 18396 20926 18452
rect 22530 18396 22540 18452
rect 22596 18396 22876 18452
rect 22932 18396 22942 18452
rect 28242 18396 28252 18452
rect 28308 18396 29036 18452
rect 29092 18396 29102 18452
rect 30034 18396 30044 18452
rect 30100 18396 30492 18452
rect 30548 18396 31500 18452
rect 31556 18396 31566 18452
rect 34290 18396 34300 18452
rect 34356 18396 34366 18452
rect 37986 18396 37996 18452
rect 38052 18396 38892 18452
rect 38948 18396 38958 18452
rect 40002 18396 40012 18452
rect 40068 18396 41468 18452
rect 41524 18396 42028 18452
rect 42084 18396 42094 18452
rect 44034 18396 44044 18452
rect 44100 18396 44716 18452
rect 44772 18396 44782 18452
rect 34300 18340 34356 18396
rect 55468 18340 55524 18508
rect 55682 18396 55692 18452
rect 55748 18396 57260 18452
rect 57316 18396 57326 18452
rect 58034 18396 58044 18452
rect 58100 18396 58828 18452
rect 58884 18396 58894 18452
rect 14578 18284 14588 18340
rect 14644 18284 15372 18340
rect 15428 18284 16156 18340
rect 16212 18284 16222 18340
rect 16818 18284 16828 18340
rect 16884 18284 18508 18340
rect 18564 18284 18574 18340
rect 20290 18284 20300 18340
rect 20356 18284 20748 18340
rect 20804 18284 20814 18340
rect 21074 18284 21084 18340
rect 21140 18284 22652 18340
rect 22708 18284 23324 18340
rect 23380 18284 23390 18340
rect 29474 18284 29484 18340
rect 29540 18284 31052 18340
rect 31108 18284 31118 18340
rect 34300 18284 40348 18340
rect 40404 18284 40796 18340
rect 40852 18284 40862 18340
rect 43026 18284 43036 18340
rect 43092 18284 43484 18340
rect 43540 18284 43550 18340
rect 48626 18284 48636 18340
rect 48692 18284 49980 18340
rect 50036 18284 51100 18340
rect 51156 18284 51166 18340
rect 55468 18284 55804 18340
rect 55860 18284 55870 18340
rect 56690 18284 56700 18340
rect 56756 18284 57820 18340
rect 57876 18284 57886 18340
rect 59052 18228 59108 18508
rect 61394 18396 61404 18452
rect 61460 18396 62412 18452
rect 62468 18396 62478 18452
rect 62850 18396 62860 18452
rect 62916 18396 63868 18452
rect 63924 18396 63934 18452
rect 68114 18396 68124 18452
rect 68180 18396 69244 18452
rect 69300 18396 69310 18452
rect 69906 18396 69916 18452
rect 69972 18396 72268 18452
rect 72324 18396 72334 18452
rect 73892 18396 75292 18452
rect 75348 18396 75358 18452
rect 73892 18340 73948 18396
rect 63522 18284 63532 18340
rect 63588 18284 64652 18340
rect 64708 18284 64718 18340
rect 64876 18284 65884 18340
rect 65940 18284 65950 18340
rect 70018 18284 70028 18340
rect 70084 18284 70812 18340
rect 70868 18284 73948 18340
rect 64876 18228 64932 18284
rect 15026 18172 15036 18228
rect 15092 18172 17164 18228
rect 17220 18172 17230 18228
rect 21970 18172 21980 18228
rect 22036 18172 22540 18228
rect 22596 18172 22606 18228
rect 27682 18172 27692 18228
rect 27748 18172 38668 18228
rect 42690 18172 42700 18228
rect 42756 18172 47628 18228
rect 47684 18172 47694 18228
rect 49298 18172 49308 18228
rect 49364 18172 51996 18228
rect 52052 18172 52062 18228
rect 53442 18172 53452 18228
rect 53508 18172 54684 18228
rect 54740 18172 59108 18228
rect 60050 18172 60060 18228
rect 60116 18172 61964 18228
rect 62020 18172 64932 18228
rect 65314 18172 65324 18228
rect 65380 18172 74396 18228
rect 74452 18172 74462 18228
rect 16482 18060 16492 18116
rect 16548 18060 19180 18116
rect 19236 18060 23996 18116
rect 24052 18060 29484 18116
rect 29540 18060 29550 18116
rect 10862 18004 10872 18060
rect 10928 18004 10976 18060
rect 11032 18004 11080 18060
rect 11136 18004 11146 18060
rect 30182 18004 30192 18060
rect 30248 18004 30296 18060
rect 30352 18004 30400 18060
rect 30456 18004 30466 18060
rect 38612 18004 38668 18172
rect 40338 18060 40348 18116
rect 40404 18060 40684 18116
rect 40740 18060 41020 18116
rect 41076 18060 41086 18116
rect 54002 18060 54012 18116
rect 54068 18060 56476 18116
rect 56532 18060 56542 18116
rect 59938 18060 59948 18116
rect 60004 18060 60620 18116
rect 60676 18060 60686 18116
rect 49502 18004 49512 18060
rect 49568 18004 49616 18060
rect 49672 18004 49720 18060
rect 49776 18004 49786 18060
rect 68822 18004 68832 18060
rect 68888 18004 68936 18060
rect 68992 18004 69040 18060
rect 69096 18004 69106 18060
rect 13794 17948 13804 18004
rect 13860 17948 18060 18004
rect 18116 17948 18126 18004
rect 20178 17948 20188 18004
rect 20244 17948 20748 18004
rect 20804 17948 20814 18004
rect 34738 17948 34748 18004
rect 34804 17948 35868 18004
rect 35924 17948 36988 18004
rect 37044 17948 37054 18004
rect 38612 17948 41244 18004
rect 41300 17948 43092 18004
rect 57250 17948 57260 18004
rect 57316 17948 58716 18004
rect 58772 17948 58782 18004
rect 18060 17892 18116 17948
rect 43036 17892 43092 17948
rect 12898 17836 12908 17892
rect 12964 17836 13580 17892
rect 13636 17836 13646 17892
rect 13804 17836 16156 17892
rect 16212 17836 16222 17892
rect 17154 17836 17164 17892
rect 17220 17836 17500 17892
rect 17556 17836 17566 17892
rect 18060 17836 25004 17892
rect 25060 17836 25070 17892
rect 25666 17836 25676 17892
rect 25732 17836 34972 17892
rect 35028 17836 35038 17892
rect 36082 17836 36092 17892
rect 36148 17836 36540 17892
rect 36596 17836 40236 17892
rect 40292 17836 40684 17892
rect 40740 17836 40750 17892
rect 43036 17836 55020 17892
rect 55076 17836 55086 17892
rect 55906 17836 55916 17892
rect 55972 17836 58156 17892
rect 58212 17836 58222 17892
rect 68786 17836 68796 17892
rect 68852 17836 71036 17892
rect 71092 17836 71102 17892
rect 73378 17836 73388 17892
rect 73444 17836 76412 17892
rect 76468 17836 77308 17892
rect 77364 17836 77374 17892
rect 5058 17724 5068 17780
rect 5124 17724 6076 17780
rect 6132 17724 11788 17780
rect 11844 17724 11854 17780
rect 12562 17724 12572 17780
rect 12628 17724 13468 17780
rect 13524 17724 13534 17780
rect 13804 17668 13860 17836
rect 23100 17780 23156 17836
rect 14242 17724 14252 17780
rect 14308 17724 14700 17780
rect 14756 17724 18172 17780
rect 18228 17724 22372 17780
rect 23090 17724 23100 17780
rect 23156 17724 23166 17780
rect 23492 17724 29372 17780
rect 29428 17724 29438 17780
rect 33394 17724 33404 17780
rect 33460 17724 35644 17780
rect 35700 17724 35710 17780
rect 43372 17724 47404 17780
rect 47460 17724 47470 17780
rect 48738 17724 48748 17780
rect 48804 17724 49308 17780
rect 49364 17724 49374 17780
rect 53666 17724 53676 17780
rect 53732 17724 54460 17780
rect 54516 17724 62412 17780
rect 62468 17724 62478 17780
rect 65986 17724 65996 17780
rect 66052 17724 69356 17780
rect 69412 17724 69422 17780
rect 75506 17724 75516 17780
rect 75572 17724 76636 17780
rect 76692 17724 76702 17780
rect 22316 17668 22372 17724
rect 23492 17668 23548 17724
rect 5282 17612 5292 17668
rect 5348 17612 13860 17668
rect 15698 17612 15708 17668
rect 15764 17612 20356 17668
rect 20738 17612 20748 17668
rect 20804 17612 21644 17668
rect 21700 17612 22092 17668
rect 22148 17612 22158 17668
rect 22316 17612 23548 17668
rect 29810 17612 29820 17668
rect 29876 17612 32620 17668
rect 32676 17612 32686 17668
rect 34626 17612 34636 17668
rect 34692 17612 37212 17668
rect 37268 17612 37278 17668
rect 20300 17556 20356 17612
rect 5842 17500 5852 17556
rect 5908 17500 6636 17556
rect 6692 17500 6702 17556
rect 11666 17500 11676 17556
rect 11732 17500 12684 17556
rect 12740 17500 12750 17556
rect 15922 17500 15932 17556
rect 15988 17500 16716 17556
rect 16772 17500 16782 17556
rect 20290 17500 20300 17556
rect 20356 17500 21420 17556
rect 21476 17500 26796 17556
rect 26852 17500 26862 17556
rect 30370 17500 30380 17556
rect 30436 17500 31276 17556
rect 31332 17500 33628 17556
rect 33684 17500 33694 17556
rect 35522 17500 35532 17556
rect 35588 17500 36204 17556
rect 36260 17500 39340 17556
rect 39396 17500 39406 17556
rect 42914 17500 42924 17556
rect 42980 17500 42990 17556
rect 42924 17444 42980 17500
rect 43372 17444 43428 17724
rect 45042 17612 45052 17668
rect 45108 17612 46396 17668
rect 46452 17612 47068 17668
rect 47124 17612 47134 17668
rect 57586 17612 57596 17668
rect 57652 17612 59388 17668
rect 59444 17612 60956 17668
rect 61012 17612 64204 17668
rect 64260 17612 64270 17668
rect 67666 17612 67676 17668
rect 67732 17612 69804 17668
rect 69860 17612 69870 17668
rect 72258 17612 72268 17668
rect 72324 17612 74956 17668
rect 75012 17612 77196 17668
rect 77252 17612 77262 17668
rect 43586 17500 43596 17556
rect 43652 17500 44268 17556
rect 44324 17500 44334 17556
rect 51314 17500 51324 17556
rect 51380 17500 52780 17556
rect 52836 17500 52846 17556
rect 58370 17500 58380 17556
rect 58436 17500 61516 17556
rect 61572 17500 63420 17556
rect 63476 17500 63486 17556
rect 67554 17500 67564 17556
rect 67620 17500 71484 17556
rect 71540 17500 73164 17556
rect 73220 17500 73230 17556
rect 6738 17388 6748 17444
rect 6804 17388 7980 17444
rect 8036 17388 8046 17444
rect 16258 17388 16268 17444
rect 16324 17388 17052 17444
rect 17108 17388 17118 17444
rect 18834 17388 18844 17444
rect 18900 17388 19964 17444
rect 20020 17388 20030 17444
rect 20300 17388 24556 17444
rect 24612 17388 25564 17444
rect 25620 17388 25630 17444
rect 34738 17388 34748 17444
rect 34804 17388 35196 17444
rect 35252 17388 38556 17444
rect 38612 17388 38622 17444
rect 39676 17388 42980 17444
rect 43362 17388 43372 17444
rect 43428 17388 43438 17444
rect 44370 17388 44380 17444
rect 44436 17388 46956 17444
rect 47012 17388 47022 17444
rect 50372 17388 63308 17444
rect 63364 17388 63374 17444
rect 63634 17388 63644 17444
rect 63700 17388 66556 17444
rect 66612 17388 66622 17444
rect 67666 17388 67676 17444
rect 67732 17388 71148 17444
rect 71204 17388 71372 17444
rect 71428 17388 71438 17444
rect 74610 17388 74620 17444
rect 74676 17388 75180 17444
rect 75236 17388 75246 17444
rect 76178 17388 76188 17444
rect 76244 17388 77308 17444
rect 77364 17388 77374 17444
rect 20300 17332 20356 17388
rect 39676 17332 39732 17388
rect 50372 17332 50428 17388
rect 15698 17276 15708 17332
rect 15764 17276 20356 17332
rect 22306 17276 22316 17332
rect 22372 17276 23212 17332
rect 23268 17276 23278 17332
rect 24098 17276 24108 17332
rect 24164 17276 24668 17332
rect 24724 17276 27804 17332
rect 27860 17276 27870 17332
rect 37538 17276 37548 17332
rect 37604 17276 39732 17332
rect 40562 17276 40572 17332
rect 40628 17276 41020 17332
rect 41076 17276 41086 17332
rect 45500 17276 50428 17332
rect 53666 17276 53676 17332
rect 53732 17276 58380 17332
rect 58436 17276 58446 17332
rect 58594 17276 58604 17332
rect 58660 17276 58772 17332
rect 58828 17276 58838 17332
rect 68898 17276 68908 17332
rect 68964 17276 70476 17332
rect 70532 17276 70542 17332
rect 20522 17220 20532 17276
rect 20588 17220 20636 17276
rect 20692 17220 20740 17276
rect 20796 17220 20806 17276
rect 39842 17220 39852 17276
rect 39908 17220 39956 17276
rect 40012 17220 40060 17276
rect 40116 17220 40126 17276
rect 14018 17164 14028 17220
rect 14084 17164 14924 17220
rect 14980 17164 14990 17220
rect 16706 17164 16716 17220
rect 16772 17164 18396 17220
rect 18452 17164 18462 17220
rect 23090 17164 23100 17220
rect 23156 17164 25676 17220
rect 25732 17164 28028 17220
rect 28084 17164 28094 17220
rect 34178 17164 34188 17220
rect 34244 17164 36428 17220
rect 36484 17164 38668 17220
rect 38724 17164 38734 17220
rect 42466 17164 42476 17220
rect 42532 17164 42924 17220
rect 42980 17164 42990 17220
rect 43250 17164 43260 17220
rect 43316 17164 44044 17220
rect 44100 17164 44110 17220
rect 45500 17108 45556 17276
rect 59162 17220 59172 17276
rect 59228 17220 59276 17276
rect 59332 17220 59380 17276
rect 59436 17220 59446 17276
rect 78482 17220 78492 17276
rect 78548 17220 78596 17276
rect 78652 17220 78700 17276
rect 78756 17220 78766 17276
rect 46050 17164 46060 17220
rect 46116 17164 46620 17220
rect 46676 17164 58548 17220
rect 68450 17164 68460 17220
rect 68516 17164 69468 17220
rect 69524 17164 69534 17220
rect 58492 17108 58548 17164
rect 3826 17052 3836 17108
rect 3892 17052 4732 17108
rect 4788 17052 4798 17108
rect 11666 17052 11676 17108
rect 11732 17052 16324 17108
rect 24322 17052 24332 17108
rect 24388 17052 25340 17108
rect 25396 17052 25406 17108
rect 27122 17052 27132 17108
rect 27188 17052 28812 17108
rect 28868 17052 35420 17108
rect 35476 17052 35486 17108
rect 40236 17052 45500 17108
rect 45556 17052 45566 17108
rect 46162 17052 46172 17108
rect 46228 17052 46844 17108
rect 46900 17052 46910 17108
rect 48626 17052 48636 17108
rect 48692 17052 54684 17108
rect 54740 17052 54750 17108
rect 57474 17052 57484 17108
rect 57540 17052 57932 17108
rect 57988 17052 57998 17108
rect 58492 17052 60060 17108
rect 60116 17052 60126 17108
rect 65090 17052 65100 17108
rect 65156 17052 66668 17108
rect 66724 17052 66734 17108
rect 71362 17052 71372 17108
rect 71428 17052 72828 17108
rect 72884 17052 72894 17108
rect 16268 16996 16324 17052
rect 12674 16940 12684 16996
rect 12740 16940 15708 16996
rect 15764 16940 15774 16996
rect 16258 16940 16268 16996
rect 16324 16940 16334 16996
rect 18834 16940 18844 16996
rect 18900 16940 18910 16996
rect 22866 16940 22876 16996
rect 22932 16940 24444 16996
rect 24500 16940 25788 16996
rect 25844 16940 25854 16996
rect 27682 16940 27692 16996
rect 27748 16940 28252 16996
rect 28308 16940 31836 16996
rect 31892 16940 31902 16996
rect 18844 16884 18900 16940
rect 11330 16828 11340 16884
rect 11396 16828 13020 16884
rect 13076 16828 13086 16884
rect 16370 16828 16380 16884
rect 16436 16828 17164 16884
rect 17220 16828 17230 16884
rect 18844 16828 19740 16884
rect 19796 16828 26684 16884
rect 26740 16828 26750 16884
rect 29250 16828 29260 16884
rect 29316 16828 30604 16884
rect 30660 16828 30670 16884
rect 32050 16828 32060 16884
rect 32116 16828 32732 16884
rect 32788 16828 32798 16884
rect 33282 16828 33292 16884
rect 33348 16828 35588 16884
rect 36754 16828 36764 16884
rect 36820 16828 38892 16884
rect 38948 16828 38958 16884
rect 8978 16716 8988 16772
rect 9044 16716 11228 16772
rect 11284 16716 11294 16772
rect 12338 16716 12348 16772
rect 12404 16716 15708 16772
rect 15764 16716 15774 16772
rect 18844 16660 18900 16828
rect 35532 16772 35588 16828
rect 40236 16772 40292 17052
rect 40786 16940 40796 16996
rect 40852 16940 41020 16996
rect 41076 16940 42588 16996
rect 42644 16940 42654 16996
rect 43138 16940 43148 16996
rect 43204 16940 43820 16996
rect 43876 16940 43886 16996
rect 50092 16940 53340 16996
rect 53396 16940 53406 16996
rect 55010 16940 55020 16996
rect 55076 16940 55748 16996
rect 50092 16884 50148 16940
rect 42354 16828 42364 16884
rect 42420 16828 43596 16884
rect 43652 16828 43662 16884
rect 43820 16828 43932 16884
rect 43988 16828 44156 16884
rect 44212 16828 44222 16884
rect 46946 16828 46956 16884
rect 47012 16828 47628 16884
rect 47684 16828 47694 16884
rect 48962 16828 48972 16884
rect 49028 16828 49924 16884
rect 50082 16828 50092 16884
rect 50148 16828 50158 16884
rect 50316 16828 54348 16884
rect 54404 16828 55468 16884
rect 55524 16828 55534 16884
rect 43820 16772 43876 16828
rect 49868 16772 49924 16828
rect 50316 16772 50372 16828
rect 55692 16772 55748 16940
rect 59052 16940 66332 16996
rect 66388 16940 67900 16996
rect 67956 16940 67966 16996
rect 69794 16940 69804 16996
rect 69860 16940 70700 16996
rect 70756 16940 70766 16996
rect 71586 16940 71596 16996
rect 71652 16940 72268 16996
rect 72324 16940 72334 16996
rect 59052 16884 59108 16940
rect 56018 16828 56028 16884
rect 56084 16828 56588 16884
rect 56644 16828 56654 16884
rect 57474 16828 57484 16884
rect 57540 16828 58492 16884
rect 58548 16828 59052 16884
rect 59108 16828 59118 16884
rect 60834 16828 60844 16884
rect 60900 16828 63868 16884
rect 63924 16828 63934 16884
rect 65538 16828 65548 16884
rect 65604 16828 66556 16884
rect 66612 16828 66622 16884
rect 69570 16828 69580 16884
rect 69636 16828 74620 16884
rect 74676 16828 74686 16884
rect 32162 16716 32172 16772
rect 32228 16716 33516 16772
rect 33572 16716 34412 16772
rect 34468 16716 34478 16772
rect 35522 16716 35532 16772
rect 35588 16716 36988 16772
rect 37044 16716 37054 16772
rect 37426 16716 37436 16772
rect 37492 16716 40292 16772
rect 41794 16716 41804 16772
rect 41860 16716 43876 16772
rect 44370 16716 44380 16772
rect 44436 16716 44828 16772
rect 44884 16716 44894 16772
rect 49868 16716 50372 16772
rect 52882 16716 52892 16772
rect 52948 16716 53900 16772
rect 53956 16716 54684 16772
rect 54740 16716 55356 16772
rect 55412 16716 55422 16772
rect 55692 16716 64876 16772
rect 64932 16716 64942 16772
rect 66210 16716 66220 16772
rect 66276 16716 67340 16772
rect 67396 16716 71484 16772
rect 71540 16716 71550 16772
rect 10882 16604 10892 16660
rect 10948 16604 12124 16660
rect 12180 16604 12190 16660
rect 18732 16604 18900 16660
rect 23650 16604 23660 16660
rect 23716 16604 24332 16660
rect 24388 16604 28476 16660
rect 28532 16604 28542 16660
rect 30044 16604 33852 16660
rect 33908 16604 33918 16660
rect 48178 16604 48188 16660
rect 48244 16604 63532 16660
rect 63588 16604 63598 16660
rect 18732 16548 18788 16604
rect 30044 16548 30100 16604
rect 11218 16492 11228 16548
rect 11284 16492 11294 16548
rect 18722 16492 18732 16548
rect 18788 16492 18798 16548
rect 22082 16492 22092 16548
rect 22148 16492 30100 16548
rect 38658 16492 38668 16548
rect 38724 16492 43932 16548
rect 43988 16492 43998 16548
rect 52210 16492 52220 16548
rect 52276 16492 52780 16548
rect 52836 16492 52846 16548
rect 53330 16492 53340 16548
rect 53396 16492 55468 16548
rect 55524 16492 55534 16548
rect 71250 16492 71260 16548
rect 71316 16492 71820 16548
rect 71876 16492 71886 16548
rect 10862 16436 10872 16492
rect 10928 16436 10976 16492
rect 11032 16436 11080 16492
rect 11136 16436 11146 16492
rect 11228 16436 11284 16492
rect 30182 16436 30192 16492
rect 30248 16436 30296 16492
rect 30352 16436 30400 16492
rect 30456 16436 30466 16492
rect 49502 16436 49512 16492
rect 49568 16436 49616 16492
rect 49672 16436 49720 16492
rect 49776 16436 49786 16492
rect 68822 16436 68832 16492
rect 68888 16436 68936 16492
rect 68992 16436 69040 16492
rect 69096 16436 69106 16492
rect 11228 16380 11564 16436
rect 11620 16380 11630 16436
rect 18946 16380 18956 16436
rect 19012 16380 19292 16436
rect 19348 16380 19358 16436
rect 24994 16380 25004 16436
rect 25060 16380 25564 16436
rect 25620 16380 25630 16436
rect 35298 16380 35308 16436
rect 35364 16380 40964 16436
rect 40908 16324 40964 16380
rect 49980 16380 56924 16436
rect 56980 16380 56990 16436
rect 57250 16380 57260 16436
rect 57316 16380 58380 16436
rect 58436 16380 58446 16436
rect 49980 16324 50036 16380
rect 10546 16268 10556 16324
rect 10612 16268 11900 16324
rect 11956 16268 11966 16324
rect 13570 16268 13580 16324
rect 13636 16268 30828 16324
rect 30884 16268 31052 16324
rect 31108 16268 31118 16324
rect 32274 16268 32284 16324
rect 32340 16268 32956 16324
rect 33012 16268 33022 16324
rect 33618 16268 33628 16324
rect 33684 16268 34300 16324
rect 34356 16268 36316 16324
rect 36372 16268 36382 16324
rect 38612 16268 40684 16324
rect 40740 16268 40750 16324
rect 40908 16268 50036 16324
rect 50194 16268 50204 16324
rect 50260 16268 62188 16324
rect 69122 16268 69132 16324
rect 69188 16268 73724 16324
rect 73780 16268 73790 16324
rect 0 16212 800 16240
rect 13580 16212 13636 16268
rect 38612 16212 38668 16268
rect 62132 16212 62188 16268
rect 79200 16212 80000 16240
rect 0 16156 1932 16212
rect 1988 16156 1998 16212
rect 5618 16156 5628 16212
rect 5684 16156 10332 16212
rect 10388 16156 10398 16212
rect 11106 16156 11116 16212
rect 11172 16156 12460 16212
rect 12516 16156 12908 16212
rect 12964 16156 13636 16212
rect 15810 16156 15820 16212
rect 15876 16156 16828 16212
rect 16884 16156 16894 16212
rect 22082 16156 22092 16212
rect 22148 16156 24444 16212
rect 24500 16156 24510 16212
rect 26338 16156 26348 16212
rect 26404 16156 35420 16212
rect 35476 16156 38668 16212
rect 39666 16156 39676 16212
rect 39732 16156 49644 16212
rect 49700 16156 50988 16212
rect 51044 16156 51054 16212
rect 51538 16156 51548 16212
rect 51604 16156 57484 16212
rect 57540 16156 57550 16212
rect 57922 16156 57932 16212
rect 57988 16156 59388 16212
rect 59444 16156 59454 16212
rect 62132 16156 76412 16212
rect 76468 16156 76972 16212
rect 77028 16156 77038 16212
rect 77970 16156 77980 16212
rect 78036 16156 80000 16212
rect 0 16128 800 16156
rect 79200 16128 80000 16156
rect 3714 16044 3724 16100
rect 3780 16044 5740 16100
rect 5796 16044 5806 16100
rect 8530 16044 8540 16100
rect 8596 16044 9324 16100
rect 9380 16044 9390 16100
rect 14354 16044 14364 16100
rect 14420 16044 15596 16100
rect 15652 16044 18956 16100
rect 19012 16044 19022 16100
rect 31378 16044 31388 16100
rect 31444 16044 33068 16100
rect 33124 16044 33134 16100
rect 35634 16044 35644 16100
rect 35700 16044 38220 16100
rect 38276 16044 38286 16100
rect 38612 16044 39116 16100
rect 39172 16044 39182 16100
rect 42802 16044 42812 16100
rect 42868 16044 43484 16100
rect 43540 16044 43550 16100
rect 43922 16044 43932 16100
rect 43988 16044 50428 16100
rect 52546 16044 52556 16100
rect 52612 16044 54348 16100
rect 54404 16044 54414 16100
rect 71922 16044 71932 16100
rect 71988 16044 73836 16100
rect 73892 16044 74396 16100
rect 74452 16044 74462 16100
rect 33068 15988 33124 16044
rect 38612 15988 38668 16044
rect 4386 15932 4396 15988
rect 4452 15932 5292 15988
rect 5348 15932 5358 15988
rect 6178 15932 6188 15988
rect 6244 15932 7532 15988
rect 7588 15932 7598 15988
rect 10098 15932 10108 15988
rect 10164 15932 11340 15988
rect 11396 15932 12348 15988
rect 12404 15932 12414 15988
rect 16930 15932 16940 15988
rect 16996 15932 17948 15988
rect 18004 15932 19852 15988
rect 19908 15932 19918 15988
rect 25778 15932 25788 15988
rect 25844 15932 27020 15988
rect 27076 15932 27468 15988
rect 27524 15932 31164 15988
rect 31220 15932 31612 15988
rect 31668 15932 31678 15988
rect 31826 15932 31836 15988
rect 31892 15932 32508 15988
rect 32564 15932 32574 15988
rect 33068 15932 35028 15988
rect 36642 15932 36652 15988
rect 36708 15932 38668 15988
rect 42354 15932 42364 15988
rect 42420 15932 50260 15988
rect 2706 15820 2716 15876
rect 2772 15820 4060 15876
rect 4116 15820 4126 15876
rect 14690 15820 14700 15876
rect 14756 15820 14766 15876
rect 20178 15820 20188 15876
rect 20244 15820 20636 15876
rect 20692 15820 26908 15876
rect 28466 15820 28476 15876
rect 28532 15820 32060 15876
rect 32116 15820 33964 15876
rect 34020 15820 34030 15876
rect 14700 15540 14756 15820
rect 20522 15652 20532 15708
rect 20588 15652 20636 15708
rect 20692 15652 20740 15708
rect 20796 15652 20806 15708
rect 26852 15652 26908 15820
rect 31714 15708 31724 15764
rect 31780 15708 33068 15764
rect 33124 15708 33134 15764
rect 34972 15652 35028 15932
rect 35186 15820 35196 15876
rect 35252 15820 35980 15876
rect 36036 15820 41020 15876
rect 41076 15820 43036 15876
rect 43092 15820 43102 15876
rect 44370 15820 44380 15876
rect 44436 15820 44716 15876
rect 44772 15820 46396 15876
rect 46452 15820 46462 15876
rect 50204 15764 50260 15932
rect 50372 15876 50428 16044
rect 51426 15932 51436 15988
rect 51492 15932 52220 15988
rect 52276 15932 54012 15988
rect 54068 15932 54078 15988
rect 54450 15932 54460 15988
rect 54516 15932 54526 15988
rect 54460 15876 54516 15932
rect 50372 15820 54516 15876
rect 57250 15820 57260 15876
rect 57316 15820 58940 15876
rect 58996 15820 59006 15876
rect 62850 15820 62860 15876
rect 62916 15820 64988 15876
rect 65044 15820 66556 15876
rect 66612 15820 67900 15876
rect 67956 15820 67966 15876
rect 42914 15708 42924 15764
rect 42980 15708 43484 15764
rect 43540 15708 43550 15764
rect 44146 15708 44156 15764
rect 44212 15708 46116 15764
rect 47954 15708 47964 15764
rect 48020 15708 48636 15764
rect 48692 15708 48702 15764
rect 50204 15708 54908 15764
rect 54964 15708 56588 15764
rect 56644 15708 58044 15764
rect 58100 15708 58110 15764
rect 63298 15708 63308 15764
rect 63364 15708 65884 15764
rect 65940 15708 65950 15764
rect 39842 15652 39852 15708
rect 39908 15652 39956 15708
rect 40012 15652 40060 15708
rect 40116 15652 40126 15708
rect 20972 15596 23548 15652
rect 23604 15596 23614 15652
rect 26852 15596 29708 15652
rect 29764 15596 31276 15652
rect 31332 15596 33628 15652
rect 33684 15596 33694 15652
rect 33842 15596 33852 15652
rect 33908 15596 34524 15652
rect 34580 15596 34590 15652
rect 34972 15596 37436 15652
rect 37492 15596 38332 15652
rect 38388 15596 38398 15652
rect 43922 15596 43932 15652
rect 43988 15596 44492 15652
rect 44548 15596 44558 15652
rect 20972 15540 21028 15596
rect 46060 15540 46116 15708
rect 59162 15652 59172 15708
rect 59228 15652 59276 15708
rect 59332 15652 59380 15708
rect 59436 15652 59446 15708
rect 78482 15652 78492 15708
rect 78548 15652 78596 15708
rect 78652 15652 78700 15708
rect 78756 15652 78766 15708
rect 60386 15596 60396 15652
rect 60452 15596 63868 15652
rect 63924 15596 67564 15652
rect 67620 15596 68348 15652
rect 68404 15596 68414 15652
rect 5954 15484 5964 15540
rect 6020 15484 7644 15540
rect 7700 15484 7710 15540
rect 14700 15484 15708 15540
rect 15764 15484 21028 15540
rect 21522 15484 21532 15540
rect 21588 15484 22204 15540
rect 22260 15484 32284 15540
rect 32340 15484 40012 15540
rect 40068 15484 42028 15540
rect 42084 15484 42812 15540
rect 42868 15484 42878 15540
rect 43698 15484 43708 15540
rect 43764 15484 44156 15540
rect 44212 15484 44222 15540
rect 46050 15484 46060 15540
rect 46116 15484 47404 15540
rect 47460 15484 47470 15540
rect 50978 15484 50988 15540
rect 51044 15484 51436 15540
rect 51492 15484 51502 15540
rect 54450 15484 54460 15540
rect 54516 15484 54796 15540
rect 54852 15484 54862 15540
rect 56914 15484 56924 15540
rect 56980 15484 59500 15540
rect 59556 15484 59566 15540
rect 15250 15372 15260 15428
rect 15316 15372 16156 15428
rect 16212 15372 19516 15428
rect 19572 15372 22876 15428
rect 22932 15372 22942 15428
rect 23436 15372 23996 15428
rect 24052 15372 24062 15428
rect 23436 15316 23492 15372
rect 31724 15316 31780 15484
rect 42690 15372 42700 15428
rect 42756 15372 50764 15428
rect 50820 15372 50830 15428
rect 4834 15260 4844 15316
rect 4900 15260 5628 15316
rect 5684 15260 5694 15316
rect 10434 15260 10444 15316
rect 10500 15260 11564 15316
rect 11620 15260 11630 15316
rect 12226 15260 12236 15316
rect 12292 15260 13132 15316
rect 13188 15260 13198 15316
rect 13906 15260 13916 15316
rect 13972 15260 14588 15316
rect 14644 15260 16604 15316
rect 16660 15260 16670 15316
rect 23426 15260 23436 15316
rect 23492 15260 23502 15316
rect 23650 15260 23660 15316
rect 23716 15260 24556 15316
rect 24612 15260 25340 15316
rect 25396 15260 25406 15316
rect 25778 15260 25788 15316
rect 25844 15260 27132 15316
rect 27188 15260 27198 15316
rect 27346 15260 27356 15316
rect 27412 15260 27422 15316
rect 28354 15260 28364 15316
rect 28420 15260 29932 15316
rect 29988 15260 29998 15316
rect 31714 15260 31724 15316
rect 31780 15260 31790 15316
rect 43362 15260 43372 15316
rect 43428 15260 44044 15316
rect 44100 15260 44110 15316
rect 27356 15204 27412 15260
rect 29932 15204 29988 15260
rect 50988 15204 51044 15484
rect 55458 15372 55468 15428
rect 55524 15372 57372 15428
rect 57428 15372 57438 15428
rect 58482 15372 58492 15428
rect 58548 15372 59276 15428
rect 59332 15372 59342 15428
rect 62962 15372 62972 15428
rect 63028 15372 64652 15428
rect 64708 15372 64718 15428
rect 12002 15148 12012 15204
rect 12068 15148 14700 15204
rect 14756 15148 14766 15204
rect 15026 15148 15036 15204
rect 15092 15148 18396 15204
rect 18452 15148 18462 15204
rect 20402 15148 20412 15204
rect 20468 15148 27412 15204
rect 28130 15148 28140 15204
rect 28196 15148 29596 15204
rect 29652 15148 29662 15204
rect 29932 15148 36764 15204
rect 36820 15148 37772 15204
rect 37828 15148 37838 15204
rect 40338 15148 40348 15204
rect 40404 15148 47012 15204
rect 48402 15148 48412 15204
rect 48468 15148 51044 15204
rect 55412 15260 56028 15316
rect 56084 15260 56812 15316
rect 56868 15260 60396 15316
rect 60452 15260 60462 15316
rect 74050 15260 74060 15316
rect 74116 15260 74732 15316
rect 74788 15260 74798 15316
rect 26348 15092 26404 15148
rect 29596 15092 29652 15148
rect 46956 15092 47012 15148
rect 55412 15092 55468 15260
rect 57138 15148 57148 15204
rect 57204 15148 57596 15204
rect 57652 15148 57820 15204
rect 57876 15148 63308 15204
rect 63364 15148 63374 15204
rect 73154 15148 73164 15204
rect 73220 15148 74396 15204
rect 74452 15148 74462 15204
rect 7186 15036 7196 15092
rect 7252 15036 8092 15092
rect 8148 15036 10556 15092
rect 10612 15036 10622 15092
rect 26338 15036 26348 15092
rect 26404 15036 26414 15092
rect 29596 15036 34188 15092
rect 34244 15036 34254 15092
rect 46956 15036 47292 15092
rect 47348 15036 48972 15092
rect 49028 15036 49038 15092
rect 51650 15036 51660 15092
rect 51716 15036 55468 15092
rect 56802 15036 56812 15092
rect 56868 15036 58156 15092
rect 58212 15036 64092 15092
rect 64148 15036 66108 15092
rect 66164 15036 66174 15092
rect 71810 15036 71820 15092
rect 71876 15036 73500 15092
rect 73556 15036 76188 15092
rect 76244 15036 76254 15092
rect 17602 14924 17612 14980
rect 17668 14924 18060 14980
rect 18116 14924 18126 14980
rect 18386 14924 18396 14980
rect 18452 14924 19068 14980
rect 19124 14924 20860 14980
rect 20916 14924 20926 14980
rect 23762 14924 23772 14980
rect 23828 14924 24780 14980
rect 24836 14924 24846 14980
rect 50866 14924 50876 14980
rect 50932 14924 52892 14980
rect 52948 14924 56140 14980
rect 56196 14924 56206 14980
rect 74162 14924 74172 14980
rect 74228 14924 74620 14980
rect 74676 14924 74686 14980
rect 10862 14868 10872 14924
rect 10928 14868 10976 14924
rect 11032 14868 11080 14924
rect 11136 14868 11146 14924
rect 30182 14868 30192 14924
rect 30248 14868 30296 14924
rect 30352 14868 30400 14924
rect 30456 14868 30466 14924
rect 49502 14868 49512 14924
rect 49568 14868 49616 14924
rect 49672 14868 49720 14924
rect 49776 14868 49786 14924
rect 68822 14868 68832 14924
rect 68888 14868 68936 14924
rect 68992 14868 69040 14924
rect 69096 14868 69106 14924
rect 13346 14812 13356 14868
rect 13412 14812 21028 14868
rect 52770 14812 52780 14868
rect 52836 14812 57260 14868
rect 57316 14812 57326 14868
rect 60722 14812 60732 14868
rect 60788 14812 63532 14868
rect 63588 14812 63598 14868
rect 9986 14700 9996 14756
rect 10052 14700 16716 14756
rect 16772 14700 17388 14756
rect 17444 14700 17454 14756
rect 20972 14644 21028 14812
rect 28578 14700 28588 14756
rect 28644 14700 28812 14756
rect 28868 14700 29932 14756
rect 29988 14700 29998 14756
rect 30258 14700 30268 14756
rect 30324 14700 38108 14756
rect 38164 14700 38556 14756
rect 38612 14700 38622 14756
rect 57362 14700 57372 14756
rect 57428 14700 57438 14756
rect 58818 14700 58828 14756
rect 58884 14700 59276 14756
rect 59332 14700 59342 14756
rect 65314 14700 65324 14756
rect 65380 14700 66220 14756
rect 66276 14700 66286 14756
rect 57372 14644 57428 14700
rect 18274 14588 18284 14644
rect 18340 14588 18844 14644
rect 18900 14588 18910 14644
rect 20972 14588 30828 14644
rect 30884 14588 30894 14644
rect 37986 14588 37996 14644
rect 38052 14588 48860 14644
rect 48916 14588 51100 14644
rect 51156 14588 51166 14644
rect 53218 14588 53228 14644
rect 53284 14588 54348 14644
rect 54404 14588 54684 14644
rect 54740 14588 54750 14644
rect 57026 14588 57036 14644
rect 57092 14588 64540 14644
rect 64596 14588 65660 14644
rect 65716 14588 65726 14644
rect 70018 14588 70028 14644
rect 70084 14588 71036 14644
rect 71092 14588 71102 14644
rect 16818 14476 16828 14532
rect 16884 14476 17500 14532
rect 17556 14476 17566 14532
rect 17714 14476 17724 14532
rect 17780 14476 18956 14532
rect 19012 14476 19022 14532
rect 28578 14476 28588 14532
rect 28644 14476 30268 14532
rect 30324 14476 30334 14532
rect 34178 14476 34188 14532
rect 34244 14476 35644 14532
rect 35700 14476 35710 14532
rect 36194 14476 36204 14532
rect 36260 14476 39900 14532
rect 39956 14476 41020 14532
rect 41076 14476 41086 14532
rect 41906 14476 41916 14532
rect 41972 14476 48300 14532
rect 48356 14476 48366 14532
rect 49298 14476 49308 14532
rect 49364 14476 50316 14532
rect 50372 14476 52108 14532
rect 52164 14476 52174 14532
rect 56690 14476 56700 14532
rect 56756 14476 58604 14532
rect 58660 14476 59444 14532
rect 59602 14476 59612 14532
rect 59668 14476 63644 14532
rect 63700 14476 63710 14532
rect 69682 14476 69692 14532
rect 69748 14476 71820 14532
rect 71876 14476 71886 14532
rect 75618 14476 75628 14532
rect 75684 14476 76860 14532
rect 76916 14476 76926 14532
rect 59388 14420 59444 14476
rect 14914 14364 14924 14420
rect 14980 14364 15260 14420
rect 15316 14364 28812 14420
rect 28868 14364 28878 14420
rect 40674 14364 40684 14420
rect 40740 14364 41692 14420
rect 41748 14364 41758 14420
rect 45602 14364 45612 14420
rect 45668 14364 46060 14420
rect 46116 14364 46126 14420
rect 47506 14364 47516 14420
rect 47572 14364 48188 14420
rect 48244 14364 52780 14420
rect 52836 14364 52846 14420
rect 56914 14364 56924 14420
rect 56980 14364 57596 14420
rect 57652 14364 57662 14420
rect 59388 14364 61292 14420
rect 61348 14364 61358 14420
rect 62738 14364 62748 14420
rect 62804 14364 63980 14420
rect 64036 14364 68236 14420
rect 68292 14364 68302 14420
rect 68898 14364 68908 14420
rect 68964 14364 70364 14420
rect 70420 14364 70430 14420
rect 76290 14364 76300 14420
rect 76356 14364 77196 14420
rect 77252 14364 77644 14420
rect 77700 14364 77710 14420
rect 5058 14252 5068 14308
rect 5124 14252 6076 14308
rect 6132 14252 17164 14308
rect 17220 14252 17948 14308
rect 18004 14252 18014 14308
rect 20178 14252 20188 14308
rect 20244 14252 21308 14308
rect 21364 14252 21374 14308
rect 27122 14252 27132 14308
rect 27188 14252 29484 14308
rect 29540 14252 29550 14308
rect 38882 14252 38892 14308
rect 38948 14252 41412 14308
rect 41570 14252 41580 14308
rect 41636 14252 47964 14308
rect 48020 14252 48030 14308
rect 58370 14252 58380 14308
rect 58436 14252 59276 14308
rect 59332 14252 64876 14308
rect 64932 14252 64942 14308
rect 76514 14252 76524 14308
rect 76580 14252 77756 14308
rect 77812 14252 77822 14308
rect 41356 14196 41412 14252
rect 15484 14140 15932 14196
rect 15988 14140 15998 14196
rect 21858 14140 21868 14196
rect 21924 14140 22148 14196
rect 24210 14140 24220 14196
rect 24276 14140 25900 14196
rect 25956 14140 25966 14196
rect 32386 14140 32396 14196
rect 32452 14140 33068 14196
rect 33124 14140 33134 14196
rect 33394 14140 33404 14196
rect 33460 14140 34524 14196
rect 34580 14140 34590 14196
rect 37548 14140 38668 14196
rect 38724 14140 38734 14196
rect 41356 14140 45612 14196
rect 45668 14140 45678 14196
rect 48850 14140 48860 14196
rect 48916 14140 50764 14196
rect 50820 14140 53004 14196
rect 53060 14140 53070 14196
rect 55234 14140 55244 14196
rect 55300 14140 55916 14196
rect 55972 14140 56364 14196
rect 56420 14140 56430 14196
rect 63522 14140 63532 14196
rect 63588 14140 65436 14196
rect 65492 14140 65502 14196
rect 12338 14028 12348 14084
rect 12404 14028 13692 14084
rect 13748 14028 13758 14084
rect 15484 13972 15540 14140
rect 20522 14084 20532 14140
rect 20588 14084 20636 14140
rect 20692 14084 20740 14140
rect 20796 14084 20806 14140
rect 22092 14084 22148 14140
rect 4834 13916 4844 13972
rect 4900 13916 8652 13972
rect 8708 13916 8718 13972
rect 10546 13916 10556 13972
rect 10612 13916 11452 13972
rect 11508 13916 11518 13972
rect 13010 13916 13020 13972
rect 13076 13916 15540 13972
rect 15708 14028 20076 14084
rect 20132 14028 20142 14084
rect 22082 14028 22092 14084
rect 22148 14028 22158 14084
rect 31154 14028 31164 14084
rect 31220 14028 37100 14084
rect 37156 14028 37166 14084
rect 15708 13860 15764 14028
rect 37548 13972 37604 14140
rect 39842 14084 39852 14140
rect 39908 14084 39956 14140
rect 40012 14084 40060 14140
rect 40116 14084 40126 14140
rect 59162 14084 59172 14140
rect 59228 14084 59276 14140
rect 59332 14084 59380 14140
rect 59436 14084 59446 14140
rect 78482 14084 78492 14140
rect 78548 14084 78596 14140
rect 78652 14084 78700 14140
rect 78756 14084 78766 14140
rect 41020 14028 55468 14084
rect 55524 14028 58268 14084
rect 58324 14028 58334 14084
rect 63858 14028 63868 14084
rect 63924 14028 65828 14084
rect 41020 13972 41076 14028
rect 65772 13972 65828 14028
rect 73892 14028 74508 14084
rect 74564 14028 74574 14084
rect 16930 13916 16940 13972
rect 16996 13916 17836 13972
rect 17892 13916 17902 13972
rect 19170 13916 19180 13972
rect 19236 13916 25788 13972
rect 25844 13916 25854 13972
rect 30034 13916 30044 13972
rect 30100 13916 33628 13972
rect 33684 13916 33694 13972
rect 33842 13916 33852 13972
rect 33908 13916 34860 13972
rect 34916 13916 37548 13972
rect 37604 13916 37614 13972
rect 38658 13916 38668 13972
rect 38724 13916 39228 13972
rect 39284 13916 41076 13972
rect 41234 13916 41244 13972
rect 41300 13916 42588 13972
rect 42644 13916 43036 13972
rect 43092 13916 43102 13972
rect 46386 13916 46396 13972
rect 46452 13916 47292 13972
rect 47348 13916 47358 13972
rect 55570 13916 55580 13972
rect 55636 13916 56812 13972
rect 56868 13916 56878 13972
rect 63522 13916 63532 13972
rect 63588 13916 65548 13972
rect 65604 13916 65614 13972
rect 65762 13916 65772 13972
rect 65828 13916 66780 13972
rect 66836 13916 66846 13972
rect 73892 13860 73948 14028
rect 74610 13916 74620 13972
rect 74676 13916 77140 13972
rect 13234 13804 13244 13860
rect 13300 13804 13916 13860
rect 13972 13804 13982 13860
rect 15092 13804 15764 13860
rect 20850 13804 20860 13860
rect 20916 13804 23100 13860
rect 23156 13804 23324 13860
rect 23380 13804 23390 13860
rect 23986 13804 23996 13860
rect 24052 13804 24892 13860
rect 24948 13804 24958 13860
rect 25554 13804 25564 13860
rect 25620 13804 26012 13860
rect 26068 13804 26078 13860
rect 31378 13804 31388 13860
rect 31444 13804 33068 13860
rect 33124 13804 33134 13860
rect 34066 13804 34076 13860
rect 34132 13804 35420 13860
rect 35476 13804 35486 13860
rect 35634 13804 35644 13860
rect 35700 13804 40908 13860
rect 40964 13804 41692 13860
rect 41748 13804 42364 13860
rect 42420 13804 42430 13860
rect 43250 13804 43260 13860
rect 43316 13804 47684 13860
rect 47842 13804 47852 13860
rect 47908 13804 50428 13860
rect 50484 13804 50494 13860
rect 53778 13804 53788 13860
rect 53844 13804 54460 13860
rect 54516 13804 55916 13860
rect 55972 13804 60732 13860
rect 60788 13804 60798 13860
rect 62132 13804 62860 13860
rect 62916 13804 62926 13860
rect 65426 13804 65436 13860
rect 65492 13804 68684 13860
rect 68740 13804 68750 13860
rect 71138 13804 71148 13860
rect 71204 13804 73276 13860
rect 73332 13804 73724 13860
rect 73780 13804 73948 13860
rect 74386 13804 74396 13860
rect 74452 13804 76860 13860
rect 76916 13804 76926 13860
rect 0 13748 800 13776
rect 15092 13748 15148 13804
rect 35644 13748 35700 13804
rect 47628 13748 47684 13804
rect 62132 13748 62188 13804
rect 77084 13748 77140 13916
rect 79200 13748 80000 13776
rect 0 13692 1932 13748
rect 1988 13692 1998 13748
rect 8642 13692 8652 13748
rect 8708 13692 15148 13748
rect 16034 13692 16044 13748
rect 16100 13692 17724 13748
rect 17780 13692 17790 13748
rect 21522 13692 21532 13748
rect 21588 13692 25228 13748
rect 25284 13692 25294 13748
rect 25442 13692 25452 13748
rect 25508 13692 26236 13748
rect 26292 13692 28252 13748
rect 28308 13692 29036 13748
rect 29092 13692 29102 13748
rect 31042 13692 31052 13748
rect 31108 13692 31500 13748
rect 31556 13692 31566 13748
rect 32498 13692 32508 13748
rect 32564 13692 34748 13748
rect 34804 13692 34814 13748
rect 34962 13692 34972 13748
rect 35028 13692 35196 13748
rect 35252 13692 35700 13748
rect 42914 13692 42924 13748
rect 42980 13692 43820 13748
rect 43876 13692 43886 13748
rect 47628 13692 48188 13748
rect 48244 13692 50092 13748
rect 50148 13692 50158 13748
rect 51650 13692 51660 13748
rect 51716 13692 52556 13748
rect 52612 13692 53340 13748
rect 53396 13692 53406 13748
rect 54898 13692 54908 13748
rect 54964 13692 56476 13748
rect 56532 13692 58044 13748
rect 58100 13692 62188 13748
rect 63410 13692 63420 13748
rect 63476 13692 66556 13748
rect 66612 13692 66622 13748
rect 68450 13692 68460 13748
rect 68516 13692 70588 13748
rect 70644 13692 71708 13748
rect 71764 13692 71774 13748
rect 72482 13692 72492 13748
rect 72548 13692 73388 13748
rect 73444 13692 73454 13748
rect 77084 13692 80000 13748
rect 0 13664 800 13692
rect 54908 13636 54964 13692
rect 79200 13664 80000 13692
rect 17826 13580 17836 13636
rect 17892 13580 18060 13636
rect 18116 13580 20188 13636
rect 20244 13580 20254 13636
rect 20514 13580 20524 13636
rect 20580 13580 21756 13636
rect 21812 13580 22988 13636
rect 23044 13580 23054 13636
rect 24098 13580 24108 13636
rect 24164 13580 25340 13636
rect 25396 13580 25406 13636
rect 26114 13580 26124 13636
rect 26180 13580 26460 13636
rect 26516 13580 26526 13636
rect 26674 13580 26684 13636
rect 26740 13580 27804 13636
rect 27860 13580 27870 13636
rect 29474 13580 29484 13636
rect 29540 13580 30716 13636
rect 30772 13580 31164 13636
rect 31220 13580 31230 13636
rect 33170 13580 33180 13636
rect 33236 13580 34076 13636
rect 34132 13580 34142 13636
rect 38434 13580 38444 13636
rect 38500 13580 45948 13636
rect 46004 13580 48300 13636
rect 48356 13580 48366 13636
rect 51762 13580 51772 13636
rect 51828 13580 54964 13636
rect 56914 13580 56924 13636
rect 56980 13580 58380 13636
rect 58436 13580 64204 13636
rect 64260 13580 66220 13636
rect 66276 13580 66286 13636
rect 11442 13468 11452 13524
rect 11508 13468 13916 13524
rect 13972 13468 14924 13524
rect 14980 13468 14990 13524
rect 17602 13468 17612 13524
rect 17668 13468 18284 13524
rect 18340 13468 18350 13524
rect 21970 13468 21980 13524
rect 22036 13468 22876 13524
rect 22932 13468 22942 13524
rect 23538 13468 23548 13524
rect 23604 13468 26908 13524
rect 26964 13468 26974 13524
rect 31826 13468 31836 13524
rect 31892 13468 34636 13524
rect 34692 13468 34702 13524
rect 37090 13468 37100 13524
rect 37156 13468 41468 13524
rect 41524 13468 41534 13524
rect 42802 13468 42812 13524
rect 42868 13468 45724 13524
rect 45780 13468 46732 13524
rect 46788 13468 46798 13524
rect 51986 13468 51996 13524
rect 52052 13468 54348 13524
rect 54404 13468 54414 13524
rect 67106 13468 67116 13524
rect 67172 13468 69580 13524
rect 69636 13468 69646 13524
rect 46732 13412 46788 13468
rect 15026 13356 15036 13412
rect 15092 13356 25452 13412
rect 25508 13356 25518 13412
rect 42130 13356 42140 13412
rect 42196 13356 42588 13412
rect 42644 13356 42654 13412
rect 44594 13356 44604 13412
rect 44660 13356 45276 13412
rect 45332 13356 45342 13412
rect 46732 13356 47292 13412
rect 47348 13356 47358 13412
rect 52098 13356 52108 13412
rect 52164 13356 57820 13412
rect 57876 13356 59724 13412
rect 59780 13356 59790 13412
rect 64530 13356 64540 13412
rect 64596 13356 66668 13412
rect 66724 13356 67900 13412
rect 67956 13356 67966 13412
rect 10862 13300 10872 13356
rect 10928 13300 10976 13356
rect 11032 13300 11080 13356
rect 11136 13300 11146 13356
rect 30182 13300 30192 13356
rect 30248 13300 30296 13356
rect 30352 13300 30400 13356
rect 30456 13300 30466 13356
rect 49502 13300 49512 13356
rect 49568 13300 49616 13356
rect 49672 13300 49720 13356
rect 49776 13300 49786 13356
rect 68822 13300 68832 13356
rect 68888 13300 68936 13356
rect 68992 13300 69040 13356
rect 69096 13300 69106 13356
rect 24994 13244 25004 13300
rect 25060 13244 25340 13300
rect 25396 13244 25406 13300
rect 25676 13244 26012 13300
rect 26068 13244 26078 13300
rect 30604 13244 37268 13300
rect 41682 13244 41692 13300
rect 41748 13244 44268 13300
rect 44324 13244 44828 13300
rect 44884 13244 48860 13300
rect 48916 13244 48926 13300
rect 56018 13244 56028 13300
rect 56084 13244 58380 13300
rect 58436 13244 58446 13300
rect 25676 13188 25732 13244
rect 30604 13188 30660 13244
rect 15250 13132 15260 13188
rect 15316 13132 15708 13188
rect 15764 13132 15774 13188
rect 24322 13132 24332 13188
rect 24388 13132 25732 13188
rect 26012 13132 26796 13188
rect 26852 13132 26862 13188
rect 27346 13132 27356 13188
rect 27412 13132 30660 13188
rect 31602 13132 31612 13188
rect 31668 13132 33292 13188
rect 33348 13132 33358 13188
rect 35298 13132 35308 13188
rect 35364 13132 36316 13188
rect 36372 13132 36382 13188
rect 26012 13076 26068 13132
rect 37212 13076 37268 13244
rect 37762 13132 37772 13188
rect 37828 13132 38220 13188
rect 38276 13132 42252 13188
rect 42308 13132 44940 13188
rect 44996 13132 45006 13188
rect 46386 13132 46396 13188
rect 46452 13132 46844 13188
rect 46900 13132 46910 13188
rect 47730 13132 47740 13188
rect 47796 13132 53564 13188
rect 53620 13132 55244 13188
rect 55300 13132 55804 13188
rect 55860 13132 55870 13188
rect 66434 13132 66444 13188
rect 66500 13132 67228 13188
rect 67284 13132 67294 13188
rect 46396 13076 46452 13132
rect 2706 13020 2716 13076
rect 2772 13020 7868 13076
rect 7924 13020 7934 13076
rect 16258 13020 16268 13076
rect 16324 13020 16940 13076
rect 16996 13020 17006 13076
rect 18274 13020 18284 13076
rect 18340 13020 21532 13076
rect 21588 13020 21598 13076
rect 21746 13020 21756 13076
rect 21812 13020 24892 13076
rect 24948 13020 24958 13076
rect 25106 13020 25116 13076
rect 25172 13020 26068 13076
rect 26226 13020 26236 13076
rect 26292 13020 26460 13076
rect 26516 13020 26526 13076
rect 27570 13020 27580 13076
rect 27636 13020 28924 13076
rect 28980 13020 28990 13076
rect 37202 13020 37212 13076
rect 37268 13020 39116 13076
rect 39172 13020 39182 13076
rect 39330 13020 39340 13076
rect 39396 13020 46452 13076
rect 48636 13020 51660 13076
rect 51716 13020 51726 13076
rect 57026 13020 57036 13076
rect 57092 13020 57372 13076
rect 57428 13020 57438 13076
rect 62850 13020 62860 13076
rect 62916 13020 63756 13076
rect 63812 13020 66892 13076
rect 66948 13020 66958 13076
rect 3602 12908 3612 12964
rect 3668 12908 5740 12964
rect 5796 12908 5806 12964
rect 19506 12908 19516 12964
rect 19572 12908 22988 12964
rect 23044 12908 24500 12964
rect 25218 12908 25228 12964
rect 25284 12908 27468 12964
rect 27524 12908 27534 12964
rect 28690 12908 28700 12964
rect 28756 12908 29260 12964
rect 29316 12908 29326 12964
rect 32722 12908 32732 12964
rect 32788 12908 33740 12964
rect 33796 12908 33806 12964
rect 34626 12908 34636 12964
rect 34692 12908 35308 12964
rect 35364 12908 35374 12964
rect 39442 12908 39452 12964
rect 39508 12908 42364 12964
rect 42420 12908 42430 12964
rect 44146 12908 44156 12964
rect 44212 12908 45276 12964
rect 45332 12908 47068 12964
rect 47124 12908 47134 12964
rect 24444 12852 24500 12908
rect 28700 12852 28756 12908
rect 12338 12796 12348 12852
rect 12404 12796 13020 12852
rect 13076 12796 14028 12852
rect 14084 12796 14094 12852
rect 17826 12796 17836 12852
rect 17892 12796 18844 12852
rect 18900 12796 18910 12852
rect 20066 12796 20076 12852
rect 20132 12796 20300 12852
rect 20356 12796 20366 12852
rect 22642 12796 22652 12852
rect 22708 12796 24220 12852
rect 24276 12796 24286 12852
rect 24444 12796 28756 12852
rect 29026 12796 29036 12852
rect 29092 12796 41356 12852
rect 41412 12796 41422 12852
rect 46386 12796 46396 12852
rect 46452 12796 46956 12852
rect 47012 12796 47852 12852
rect 47908 12796 47918 12852
rect 48636 12740 48692 13020
rect 48962 12908 48972 12964
rect 49028 12908 51100 12964
rect 51156 12908 51166 12964
rect 52434 12908 52444 12964
rect 52500 12908 53452 12964
rect 53508 12908 55356 12964
rect 55412 12908 56924 12964
rect 56980 12908 56990 12964
rect 58370 12908 58380 12964
rect 58436 12908 65548 12964
rect 65604 12908 67452 12964
rect 67508 12908 67518 12964
rect 57026 12796 57036 12852
rect 57092 12796 57932 12852
rect 57988 12796 57998 12852
rect 59714 12796 59724 12852
rect 59780 12796 62188 12852
rect 15810 12684 15820 12740
rect 15876 12684 16156 12740
rect 16212 12684 16222 12740
rect 17266 12684 17276 12740
rect 17332 12684 19964 12740
rect 20020 12684 20030 12740
rect 20300 12684 21756 12740
rect 21812 12684 21822 12740
rect 23762 12684 23772 12740
rect 23828 12684 24108 12740
rect 24164 12684 24174 12740
rect 24434 12684 24444 12740
rect 24500 12684 25452 12740
rect 25508 12684 25518 12740
rect 31938 12684 31948 12740
rect 32004 12684 32956 12740
rect 33012 12684 33022 12740
rect 35634 12684 35644 12740
rect 35700 12684 35980 12740
rect 36036 12684 39732 12740
rect 40002 12684 40012 12740
rect 40068 12684 41132 12740
rect 41188 12684 41198 12740
rect 45602 12684 45612 12740
rect 45668 12684 46732 12740
rect 46788 12684 48636 12740
rect 48692 12684 48702 12740
rect 20300 12628 20356 12684
rect 16706 12572 16716 12628
rect 16772 12572 17948 12628
rect 18004 12572 20356 12628
rect 23650 12572 23660 12628
rect 23716 12572 24780 12628
rect 24836 12572 24846 12628
rect 31714 12572 31724 12628
rect 31780 12572 32732 12628
rect 32788 12572 32798 12628
rect 38098 12572 38108 12628
rect 38164 12572 39340 12628
rect 39396 12572 39406 12628
rect 20522 12516 20532 12572
rect 20588 12516 20636 12572
rect 20692 12516 20740 12572
rect 20796 12516 20806 12572
rect 16818 12460 16828 12516
rect 16884 12460 18284 12516
rect 18340 12460 18350 12516
rect 23202 12460 23212 12516
rect 23268 12460 24668 12516
rect 24724 12460 36428 12516
rect 36484 12460 38668 12516
rect 30818 12348 30828 12404
rect 30884 12348 33516 12404
rect 33572 12348 33582 12404
rect 33842 12348 33852 12404
rect 33908 12348 34524 12404
rect 34580 12348 36092 12404
rect 36148 12348 36158 12404
rect 38612 12292 38668 12460
rect 39676 12404 39732 12684
rect 62132 12628 62188 12796
rect 73892 12740 73948 12964
rect 74004 12908 74014 12964
rect 63970 12684 63980 12740
rect 64036 12684 64652 12740
rect 64708 12684 65548 12740
rect 65604 12684 65614 12740
rect 73266 12684 73276 12740
rect 73332 12684 73948 12740
rect 75618 12684 75628 12740
rect 75684 12684 76860 12740
rect 76916 12684 76926 12740
rect 50372 12572 58156 12628
rect 58212 12572 58222 12628
rect 62132 12572 63868 12628
rect 63924 12572 63934 12628
rect 73042 12572 73052 12628
rect 73108 12572 74172 12628
rect 74228 12572 74238 12628
rect 39842 12516 39852 12572
rect 39908 12516 39956 12572
rect 40012 12516 40060 12572
rect 40116 12516 40126 12572
rect 50372 12516 50428 12572
rect 59162 12516 59172 12572
rect 59228 12516 59276 12572
rect 59332 12516 59380 12572
rect 59436 12516 59446 12572
rect 78482 12516 78492 12572
rect 78548 12516 78596 12572
rect 78652 12516 78700 12572
rect 78756 12516 78766 12572
rect 42140 12460 50428 12516
rect 59612 12460 65100 12516
rect 65156 12460 65660 12516
rect 65716 12460 65726 12516
rect 42140 12404 42196 12460
rect 59612 12404 59668 12460
rect 39676 12348 39900 12404
rect 39956 12348 42196 12404
rect 42354 12348 42364 12404
rect 42420 12348 48972 12404
rect 49028 12348 49038 12404
rect 52882 12348 52892 12404
rect 52948 12348 57372 12404
rect 57428 12348 59052 12404
rect 59108 12348 59668 12404
rect 60386 12348 60396 12404
rect 60452 12348 61068 12404
rect 61124 12348 61134 12404
rect 61730 12348 61740 12404
rect 61796 12348 62188 12404
rect 62244 12348 62254 12404
rect 23874 12236 23884 12292
rect 23940 12236 27972 12292
rect 28130 12236 28140 12292
rect 28196 12236 28700 12292
rect 28756 12236 28766 12292
rect 31378 12236 31388 12292
rect 31444 12236 33292 12292
rect 33348 12236 33358 12292
rect 38612 12236 40348 12292
rect 40404 12236 41804 12292
rect 41860 12236 41870 12292
rect 44482 12236 44492 12292
rect 44548 12236 45500 12292
rect 45556 12236 46620 12292
rect 46676 12236 46686 12292
rect 57250 12236 57260 12292
rect 57316 12236 57932 12292
rect 57988 12236 58828 12292
rect 58884 12236 58894 12292
rect 59378 12236 59388 12292
rect 59444 12236 59836 12292
rect 59892 12236 59902 12292
rect 70802 12236 70812 12292
rect 70868 12236 72380 12292
rect 72436 12236 72446 12292
rect 27916 12180 27972 12236
rect 1810 12124 1820 12180
rect 1876 12124 5516 12180
rect 5572 12124 5582 12180
rect 12002 12124 12012 12180
rect 12068 12124 12684 12180
rect 12740 12124 12750 12180
rect 15698 12124 15708 12180
rect 15764 12124 16492 12180
rect 16548 12124 16558 12180
rect 20066 12124 20076 12180
rect 20132 12124 20142 12180
rect 24322 12124 24332 12180
rect 24388 12124 25676 12180
rect 25732 12124 25742 12180
rect 27916 12124 28588 12180
rect 28644 12124 28654 12180
rect 35074 12124 35084 12180
rect 35140 12124 37772 12180
rect 37828 12124 37838 12180
rect 43474 12124 43484 12180
rect 43540 12124 47628 12180
rect 47684 12124 47694 12180
rect 50372 12124 52332 12180
rect 52388 12124 52398 12180
rect 56354 12124 56364 12180
rect 56420 12124 58044 12180
rect 58100 12124 58110 12180
rect 58258 12124 58268 12180
rect 58324 12124 60396 12180
rect 60452 12124 60462 12180
rect 63858 12124 63868 12180
rect 63924 12124 66892 12180
rect 66948 12124 69244 12180
rect 69300 12124 69310 12180
rect 20076 12068 20132 12124
rect 50372 12068 50428 12124
rect 12898 12012 12908 12068
rect 12964 12012 15820 12068
rect 15876 12012 15886 12068
rect 16258 12012 16268 12068
rect 16324 12012 18620 12068
rect 18676 12012 19292 12068
rect 19348 12012 19358 12068
rect 20076 12012 20916 12068
rect 21746 12012 21756 12068
rect 21812 12012 22204 12068
rect 22260 12012 22270 12068
rect 25442 12012 25452 12068
rect 25508 12012 26236 12068
rect 26292 12012 26796 12068
rect 26852 12012 39004 12068
rect 39060 12012 41692 12068
rect 41748 12012 42812 12068
rect 42868 12012 43932 12068
rect 43988 12012 43998 12068
rect 50082 12012 50092 12068
rect 50148 12012 50428 12068
rect 56914 12012 56924 12068
rect 56980 12012 62412 12068
rect 62468 12012 63308 12068
rect 63364 12012 63374 12068
rect 20860 11956 20916 12012
rect 18834 11900 18844 11956
rect 18900 11900 19516 11956
rect 19572 11900 19582 11956
rect 20066 11900 20076 11956
rect 20132 11900 20142 11956
rect 20850 11900 20860 11956
rect 20916 11900 20926 11956
rect 24098 11900 24108 11956
rect 24164 11900 25676 11956
rect 25732 11900 26124 11956
rect 26180 11900 29036 11956
rect 29092 11900 29102 11956
rect 33058 11900 33068 11956
rect 33124 11900 38668 11956
rect 38724 11900 38734 11956
rect 43026 11900 43036 11956
rect 43092 11900 48748 11956
rect 48804 11900 53788 11956
rect 53844 11900 53854 11956
rect 54562 11900 54572 11956
rect 54628 11900 56700 11956
rect 56756 11900 56766 11956
rect 58034 11900 58044 11956
rect 58100 11900 64540 11956
rect 64596 11900 64606 11956
rect 20076 11844 20132 11900
rect 12674 11788 12684 11844
rect 12740 11788 13020 11844
rect 13076 11788 13086 11844
rect 13794 11788 13804 11844
rect 13860 11788 15148 11844
rect 15204 11788 15484 11844
rect 15540 11788 15550 11844
rect 18274 11788 18284 11844
rect 18340 11788 26572 11844
rect 26628 11788 26638 11844
rect 36194 11788 36204 11844
rect 36260 11788 44604 11844
rect 44660 11788 44670 11844
rect 54226 11788 54236 11844
rect 54292 11788 54908 11844
rect 54964 11788 54974 11844
rect 55122 11788 55132 11844
rect 55188 11788 57036 11844
rect 57092 11788 57102 11844
rect 10862 11732 10872 11788
rect 10928 11732 10976 11788
rect 11032 11732 11080 11788
rect 11136 11732 11146 11788
rect 30182 11732 30192 11788
rect 30248 11732 30296 11788
rect 30352 11732 30400 11788
rect 30456 11732 30466 11788
rect 49502 11732 49512 11788
rect 49568 11732 49616 11788
rect 49672 11732 49720 11788
rect 49776 11732 49786 11788
rect 68822 11732 68832 11788
rect 68888 11732 68936 11788
rect 68992 11732 69040 11788
rect 69096 11732 69106 11788
rect 18386 11676 18396 11732
rect 18452 11676 19740 11732
rect 19796 11676 19806 11732
rect 20962 11676 20972 11732
rect 21028 11676 21038 11732
rect 23650 11676 23660 11732
rect 23716 11676 24220 11732
rect 24276 11676 29092 11732
rect 33394 11676 33404 11732
rect 33460 11676 34188 11732
rect 34244 11676 34254 11732
rect 37314 11676 37324 11732
rect 37380 11676 38668 11732
rect 38724 11676 38734 11732
rect 42354 11676 42364 11732
rect 42420 11676 47180 11732
rect 47236 11676 47246 11732
rect 52098 11676 52108 11732
rect 52164 11676 65212 11732
rect 65268 11676 65278 11732
rect 65426 11676 65436 11732
rect 65492 11676 66780 11732
rect 66836 11676 67228 11732
rect 67284 11676 67294 11732
rect 17266 11564 17276 11620
rect 17332 11564 17612 11620
rect 17668 11564 19180 11620
rect 19236 11564 19246 11620
rect 20972 11508 21028 11676
rect 22194 11564 22204 11620
rect 22260 11564 23884 11620
rect 23940 11564 23950 11620
rect 24434 11564 24444 11620
rect 24500 11564 25340 11620
rect 25396 11564 28028 11620
rect 28084 11564 28094 11620
rect 29036 11508 29092 11676
rect 29250 11564 29260 11620
rect 29316 11564 76524 11620
rect 76580 11564 76590 11620
rect 4274 11452 4284 11508
rect 4340 11452 5068 11508
rect 5124 11452 5134 11508
rect 6962 11452 6972 11508
rect 7028 11452 8316 11508
rect 8372 11452 8382 11508
rect 20972 11452 21308 11508
rect 21364 11452 21374 11508
rect 21868 11452 25564 11508
rect 25620 11452 25630 11508
rect 25778 11452 25788 11508
rect 25844 11452 27244 11508
rect 27300 11452 27310 11508
rect 29036 11452 39004 11508
rect 39060 11452 40124 11508
rect 40180 11452 40796 11508
rect 40852 11452 42140 11508
rect 42196 11452 43148 11508
rect 43204 11452 43214 11508
rect 48514 11452 48524 11508
rect 48580 11452 50204 11508
rect 50260 11452 50270 11508
rect 59042 11452 59052 11508
rect 59108 11452 60732 11508
rect 60788 11452 60798 11508
rect 65202 11452 65212 11508
rect 65268 11452 68124 11508
rect 68180 11452 68190 11508
rect 21868 11396 21924 11452
rect 12114 11340 12124 11396
rect 12180 11340 12796 11396
rect 12852 11340 12862 11396
rect 16482 11340 16492 11396
rect 16548 11340 16828 11396
rect 16884 11340 16894 11396
rect 20850 11340 20860 11396
rect 20916 11340 21924 11396
rect 22754 11340 22764 11396
rect 22820 11340 23436 11396
rect 23492 11340 23502 11396
rect 23986 11340 23996 11396
rect 24052 11340 24892 11396
rect 24948 11340 24958 11396
rect 28130 11340 28140 11396
rect 28196 11340 29260 11396
rect 29316 11340 37996 11396
rect 38052 11340 43484 11396
rect 43540 11340 43820 11396
rect 43876 11340 44940 11396
rect 44996 11340 45006 11396
rect 49970 11340 49980 11396
rect 50036 11340 51548 11396
rect 51604 11340 53116 11396
rect 53172 11340 53182 11396
rect 75618 11340 75628 11396
rect 75684 11340 76748 11396
rect 76804 11340 76814 11396
rect 0 11284 800 11312
rect 28140 11284 28196 11340
rect 79200 11284 80000 11312
rect 0 11228 1932 11284
rect 1988 11228 1998 11284
rect 15474 11228 15484 11284
rect 15540 11228 16940 11284
rect 16996 11228 18620 11284
rect 18676 11228 18686 11284
rect 20402 11228 20412 11284
rect 20468 11228 22540 11284
rect 22596 11228 22606 11284
rect 23650 11228 23660 11284
rect 23716 11228 24108 11284
rect 24164 11228 24174 11284
rect 24546 11228 24556 11284
rect 24612 11228 25788 11284
rect 25844 11228 28196 11284
rect 30706 11228 30716 11284
rect 30772 11228 31724 11284
rect 31780 11228 31790 11284
rect 34178 11228 34188 11284
rect 34244 11228 37884 11284
rect 37940 11228 38220 11284
rect 38276 11228 38286 11284
rect 39330 11228 39340 11284
rect 39396 11228 41132 11284
rect 41188 11228 41804 11284
rect 41860 11228 41870 11284
rect 48178 11228 48188 11284
rect 48244 11228 50428 11284
rect 50484 11228 50494 11284
rect 52098 11228 52108 11284
rect 52164 11228 52780 11284
rect 52836 11228 52846 11284
rect 59490 11228 59500 11284
rect 59556 11228 60396 11284
rect 60452 11228 60462 11284
rect 70242 11228 70252 11284
rect 70308 11228 72604 11284
rect 72660 11228 72670 11284
rect 74620 11228 80000 11284
rect 0 11200 800 11228
rect 74620 11172 74676 11228
rect 79200 11200 80000 11228
rect 7746 11116 7756 11172
rect 7812 11116 8764 11172
rect 8820 11116 10444 11172
rect 10500 11116 10510 11172
rect 11778 11116 11788 11172
rect 11844 11116 14028 11172
rect 14084 11116 15148 11172
rect 16370 11116 16380 11172
rect 16436 11116 17500 11172
rect 17556 11116 17566 11172
rect 18050 11116 18060 11172
rect 18116 11116 21028 11172
rect 22866 11116 22876 11172
rect 22932 11116 24220 11172
rect 24276 11116 24286 11172
rect 26338 11116 26348 11172
rect 26404 11116 27804 11172
rect 27860 11116 27870 11172
rect 28466 11116 28476 11172
rect 28532 11116 30156 11172
rect 30212 11116 30222 11172
rect 32498 11116 32508 11172
rect 32564 11116 36428 11172
rect 36484 11116 37324 11172
rect 37380 11116 37390 11172
rect 39452 11116 41356 11172
rect 41412 11116 42476 11172
rect 42532 11116 42812 11172
rect 42868 11116 42878 11172
rect 45490 11116 45500 11172
rect 45556 11116 45948 11172
rect 46004 11116 46014 11172
rect 53890 11116 53900 11172
rect 53956 11116 54460 11172
rect 54516 11116 59388 11172
rect 59444 11116 61068 11172
rect 61124 11116 65436 11172
rect 65492 11116 65502 11172
rect 74610 11116 74620 11172
rect 74676 11116 74686 11172
rect 15092 10948 15148 11116
rect 20972 11060 21028 11116
rect 26348 11060 26404 11116
rect 39452 11060 39508 11116
rect 20972 11004 26404 11060
rect 28018 11004 28028 11060
rect 28084 11004 29708 11060
rect 29764 11004 36988 11060
rect 37044 11004 39452 11060
rect 39508 11004 39518 11060
rect 44594 11004 44604 11060
rect 44660 11004 48748 11060
rect 48804 11004 48814 11060
rect 56802 11004 56812 11060
rect 56868 11004 58716 11060
rect 58772 11004 58782 11060
rect 20522 10948 20532 11004
rect 20588 10948 20636 11004
rect 20692 10948 20740 11004
rect 20796 10948 20806 11004
rect 39842 10948 39852 11004
rect 39908 10948 39956 11004
rect 40012 10948 40060 11004
rect 40116 10948 40126 11004
rect 59162 10948 59172 11004
rect 59228 10948 59276 11004
rect 59332 10948 59380 11004
rect 59436 10948 59446 11004
rect 78482 10948 78492 11004
rect 78548 10948 78596 11004
rect 78652 10948 78700 11004
rect 78756 10948 78766 11004
rect 15092 10892 20356 10948
rect 22306 10892 22316 10948
rect 22372 10892 23548 10948
rect 23604 10892 23614 10948
rect 23986 10892 23996 10948
rect 24052 10892 24164 10948
rect 25442 10892 25452 10948
rect 25508 10892 25788 10948
rect 25844 10892 25854 10948
rect 40786 10892 40796 10948
rect 40852 10892 41356 10948
rect 41412 10892 42588 10948
rect 42644 10892 50092 10948
rect 50148 10892 50158 10948
rect 71250 10892 71260 10948
rect 71316 10892 72380 10948
rect 72436 10892 72446 10948
rect 3154 10780 3164 10836
rect 3220 10780 4732 10836
rect 4788 10780 4798 10836
rect 6178 10780 6188 10836
rect 6244 10780 8036 10836
rect 15922 10780 15932 10836
rect 15988 10780 17276 10836
rect 17332 10780 17342 10836
rect 7980 10724 8036 10780
rect 20300 10724 20356 10892
rect 21410 10780 21420 10836
rect 21476 10780 21756 10836
rect 21812 10780 21822 10836
rect 5170 10668 5180 10724
rect 5236 10668 5852 10724
rect 5908 10668 7532 10724
rect 7588 10668 7598 10724
rect 7970 10668 7980 10724
rect 8036 10668 9548 10724
rect 9604 10668 9614 10724
rect 11218 10668 11228 10724
rect 11284 10668 12012 10724
rect 12068 10668 19852 10724
rect 19908 10668 19918 10724
rect 20300 10668 22652 10724
rect 22708 10668 23660 10724
rect 23716 10668 23726 10724
rect 11228 10612 11284 10668
rect 24108 10612 24164 10892
rect 24546 10780 24556 10836
rect 24612 10780 24622 10836
rect 28578 10780 28588 10836
rect 28644 10780 76412 10836
rect 76468 10780 76972 10836
rect 77028 10780 77038 10836
rect 5618 10556 5628 10612
rect 5684 10556 6972 10612
rect 7028 10556 7038 10612
rect 7196 10556 11284 10612
rect 11778 10556 11788 10612
rect 11844 10556 12796 10612
rect 12852 10556 22204 10612
rect 22260 10556 22270 10612
rect 24098 10556 24108 10612
rect 24164 10556 24174 10612
rect 7196 10500 7252 10556
rect 24556 10500 24612 10780
rect 6626 10444 6636 10500
rect 6692 10444 7252 10500
rect 10098 10444 10108 10500
rect 10164 10444 10556 10500
rect 10612 10444 11340 10500
rect 11396 10444 11406 10500
rect 12898 10444 12908 10500
rect 12964 10444 15708 10500
rect 15764 10444 15774 10500
rect 17490 10444 17500 10500
rect 17556 10444 18508 10500
rect 18564 10444 19628 10500
rect 19684 10444 19694 10500
rect 19842 10444 19852 10500
rect 19908 10444 22764 10500
rect 22820 10444 24612 10500
rect 26852 10668 27468 10724
rect 27524 10668 28644 10724
rect 39330 10668 39340 10724
rect 39396 10668 40012 10724
rect 40068 10668 40078 10724
rect 55906 10668 55916 10724
rect 55972 10668 56924 10724
rect 56980 10668 56990 10724
rect 64978 10668 64988 10724
rect 65044 10668 67788 10724
rect 67844 10668 67854 10724
rect 68114 10668 68124 10724
rect 68180 10668 69356 10724
rect 69412 10668 69422 10724
rect 70130 10668 70140 10724
rect 70196 10668 70476 10724
rect 70532 10668 72604 10724
rect 72660 10668 72670 10724
rect 73378 10668 73388 10724
rect 73444 10668 74172 10724
rect 74228 10668 74238 10724
rect 4610 10332 4620 10388
rect 4676 10332 5068 10388
rect 5124 10332 5134 10388
rect 16034 10332 16044 10388
rect 16100 10332 21532 10388
rect 21588 10332 21598 10388
rect 23986 10332 23996 10388
rect 24052 10332 25340 10388
rect 25396 10332 25406 10388
rect 26852 10276 26908 10668
rect 28588 10612 28644 10668
rect 69356 10612 69412 10668
rect 28578 10556 28588 10612
rect 28644 10556 37660 10612
rect 37716 10556 43148 10612
rect 43204 10556 43214 10612
rect 43810 10556 43820 10612
rect 43876 10556 50652 10612
rect 50708 10556 50718 10612
rect 65986 10556 65996 10612
rect 66052 10556 66780 10612
rect 66836 10556 66846 10612
rect 69356 10556 71708 10612
rect 71764 10556 71774 10612
rect 43148 10500 43204 10556
rect 15474 10220 15484 10276
rect 15540 10220 15708 10276
rect 15764 10220 17388 10276
rect 17444 10220 17454 10276
rect 23762 10220 23772 10276
rect 23828 10220 25788 10276
rect 25844 10220 26908 10276
rect 32396 10444 38668 10500
rect 38724 10444 39676 10500
rect 39732 10444 39742 10500
rect 43148 10444 44268 10500
rect 44324 10444 44334 10500
rect 45490 10444 45500 10500
rect 45556 10444 53676 10500
rect 53732 10444 53742 10500
rect 63858 10444 63868 10500
rect 63924 10444 65660 10500
rect 65716 10444 65726 10500
rect 68562 10444 68572 10500
rect 68628 10444 69132 10500
rect 69188 10444 69916 10500
rect 69972 10444 69982 10500
rect 72706 10444 72716 10500
rect 72772 10444 75516 10500
rect 75572 10444 75582 10500
rect 10862 10164 10872 10220
rect 10928 10164 10976 10220
rect 11032 10164 11080 10220
rect 11136 10164 11146 10220
rect 30182 10164 30192 10220
rect 30248 10164 30296 10220
rect 30352 10164 30400 10220
rect 30456 10164 30466 10220
rect 11666 10108 11676 10164
rect 11732 10108 12012 10164
rect 12068 10108 12078 10164
rect 20076 10108 21196 10164
rect 21252 10108 21756 10164
rect 21812 10108 22876 10164
rect 22932 10108 22942 10164
rect 23314 10108 23324 10164
rect 23380 10108 24108 10164
rect 24164 10108 24174 10164
rect 24882 10108 24892 10164
rect 24948 10108 25564 10164
rect 25620 10108 25630 10164
rect 28242 10108 28252 10164
rect 28308 10108 30100 10164
rect 20076 10052 20132 10108
rect 30044 10052 30100 10108
rect 32396 10052 32452 10444
rect 38546 10332 38556 10388
rect 38612 10332 41580 10388
rect 41636 10332 41646 10388
rect 42354 10332 42364 10388
rect 42420 10332 43484 10388
rect 43540 10332 43550 10388
rect 47180 10332 76076 10388
rect 76132 10332 77644 10388
rect 77700 10332 77710 10388
rect 5058 9996 5068 10052
rect 5124 9996 6412 10052
rect 6468 9996 20132 10052
rect 20290 9996 20300 10052
rect 20356 9996 21308 10052
rect 21364 9996 21374 10052
rect 21522 9996 21532 10052
rect 21588 9996 25116 10052
rect 25172 9996 25182 10052
rect 30044 9996 30492 10052
rect 30548 9996 30558 10052
rect 32386 9996 32396 10052
rect 32452 9996 32462 10052
rect 37874 9996 37884 10052
rect 37940 9996 43036 10052
rect 43092 9996 43102 10052
rect 43250 9996 43260 10052
rect 43316 9996 45276 10052
rect 45332 9996 45342 10052
rect 47180 9940 47236 10332
rect 54338 10220 54348 10276
rect 54404 10220 55132 10276
rect 55188 10220 56812 10276
rect 56868 10220 56878 10276
rect 73378 10220 73388 10276
rect 73444 10220 74060 10276
rect 74116 10220 74126 10276
rect 49502 10164 49512 10220
rect 49568 10164 49616 10220
rect 49672 10164 49720 10220
rect 49776 10164 49786 10220
rect 68822 10164 68832 10220
rect 68888 10164 68936 10220
rect 68992 10164 69040 10220
rect 69096 10164 69106 10220
rect 72370 10108 72380 10164
rect 72436 10108 73612 10164
rect 73668 10108 73678 10164
rect 51314 9996 51324 10052
rect 51380 9996 53508 10052
rect 68898 9996 68908 10052
rect 68964 9996 69468 10052
rect 69524 9996 69534 10052
rect 72930 9996 72940 10052
rect 72996 9996 74284 10052
rect 74340 9996 74350 10052
rect 53452 9940 53508 9996
rect 73612 9940 73668 9996
rect 4722 9884 4732 9940
rect 4788 9884 6188 9940
rect 6244 9884 6254 9940
rect 14242 9884 14252 9940
rect 14308 9884 15372 9940
rect 15428 9884 15438 9940
rect 19730 9884 19740 9940
rect 19796 9884 19806 9940
rect 20738 9884 20748 9940
rect 20804 9884 21868 9940
rect 21924 9884 21934 9940
rect 26852 9884 47236 9940
rect 49298 9884 49308 9940
rect 49364 9884 51436 9940
rect 51492 9884 51502 9940
rect 53442 9884 53452 9940
rect 53508 9884 55804 9940
rect 55860 9884 55870 9940
rect 57922 9884 57932 9940
rect 57988 9884 61068 9940
rect 61124 9884 61134 9940
rect 69794 9884 69804 9940
rect 69860 9884 71372 9940
rect 71428 9884 71438 9940
rect 73602 9884 73612 9940
rect 73668 9884 73678 9940
rect 19740 9828 19796 9884
rect 26852 9828 26908 9884
rect 4162 9772 4172 9828
rect 4228 9772 4620 9828
rect 4676 9772 5740 9828
rect 5796 9772 11788 9828
rect 11844 9772 11854 9828
rect 13570 9772 13580 9828
rect 13636 9772 14476 9828
rect 14532 9772 14542 9828
rect 19740 9772 26908 9828
rect 34850 9772 34860 9828
rect 34916 9772 35868 9828
rect 35924 9772 35934 9828
rect 37314 9772 37324 9828
rect 37380 9772 47348 9828
rect 48738 9772 48748 9828
rect 48804 9772 50988 9828
rect 51044 9772 51054 9828
rect 51884 9772 53228 9828
rect 53284 9772 53294 9828
rect 68562 9772 68572 9828
rect 68628 9772 70700 9828
rect 70756 9772 70766 9828
rect 72034 9772 72044 9828
rect 72100 9772 72492 9828
rect 72548 9772 73500 9828
rect 73556 9772 73566 9828
rect 47292 9716 47348 9772
rect 51884 9716 51940 9772
rect 3154 9660 3164 9716
rect 3220 9660 3836 9716
rect 3892 9660 3902 9716
rect 17826 9660 17836 9716
rect 17892 9660 19628 9716
rect 19684 9660 22092 9716
rect 22148 9660 28476 9716
rect 28532 9660 28542 9716
rect 30482 9660 30492 9716
rect 30548 9660 31500 9716
rect 31556 9660 32396 9716
rect 32452 9660 32462 9716
rect 46162 9660 46172 9716
rect 46228 9660 47068 9716
rect 47124 9660 47134 9716
rect 47292 9660 51940 9716
rect 53116 9660 64988 9716
rect 65044 9660 65884 9716
rect 65940 9660 72940 9716
rect 72996 9660 73006 9716
rect 19852 9548 20636 9604
rect 20692 9548 20702 9604
rect 26852 9548 50428 9604
rect 51986 9548 51996 9604
rect 52052 9548 52892 9604
rect 52948 9548 52958 9604
rect 19852 9492 19908 9548
rect 26852 9492 26908 9548
rect 7858 9436 7868 9492
rect 7924 9436 10780 9492
rect 10836 9436 19852 9492
rect 19908 9436 19918 9492
rect 26450 9436 26460 9492
rect 26516 9436 26908 9492
rect 43026 9436 43036 9492
rect 43092 9436 47740 9492
rect 47796 9436 47806 9492
rect 20522 9380 20532 9436
rect 20588 9380 20636 9436
rect 20692 9380 20740 9436
rect 20796 9380 20806 9436
rect 39842 9380 39852 9436
rect 39908 9380 39956 9436
rect 40012 9380 40060 9436
rect 40116 9380 40126 9436
rect 50372 9380 50428 9548
rect 53116 9492 53172 9660
rect 50978 9436 50988 9492
rect 51044 9436 53172 9492
rect 53340 9548 76300 9604
rect 76356 9548 76366 9604
rect 53340 9380 53396 9548
rect 73490 9436 73500 9492
rect 73556 9436 74060 9492
rect 74116 9436 74126 9492
rect 59162 9380 59172 9436
rect 59228 9380 59276 9436
rect 59332 9380 59380 9436
rect 59436 9380 59446 9436
rect 78482 9380 78492 9436
rect 78548 9380 78596 9436
rect 78652 9380 78700 9436
rect 78756 9380 78766 9436
rect 10210 9324 10220 9380
rect 10276 9324 12348 9380
rect 12404 9324 13916 9380
rect 13972 9324 13982 9380
rect 50372 9324 53396 9380
rect 71026 9324 71036 9380
rect 71092 9324 72268 9380
rect 72324 9324 73276 9380
rect 73332 9324 73836 9380
rect 73892 9324 73902 9380
rect 4274 9212 4284 9268
rect 4340 9212 5292 9268
rect 5348 9212 34972 9268
rect 35028 9212 35038 9268
rect 48066 9212 48076 9268
rect 48132 9212 49644 9268
rect 49700 9212 49710 9268
rect 61282 9212 61292 9268
rect 61348 9212 63140 9268
rect 63084 9156 63140 9212
rect 5506 9100 5516 9156
rect 5572 9100 7084 9156
rect 7140 9100 8428 9156
rect 8484 9100 8494 9156
rect 10658 9100 10668 9156
rect 10724 9100 11452 9156
rect 11508 9100 12796 9156
rect 12852 9100 12862 9156
rect 13570 9100 13580 9156
rect 13636 9100 14028 9156
rect 14084 9100 20748 9156
rect 20804 9100 42812 9156
rect 42868 9100 42878 9156
rect 45938 9100 45948 9156
rect 46004 9100 47180 9156
rect 47236 9100 48860 9156
rect 48916 9100 48926 9156
rect 62132 9100 62524 9156
rect 62580 9100 62590 9156
rect 63074 9100 63084 9156
rect 63140 9100 63756 9156
rect 63812 9100 63822 9156
rect 18834 8988 18844 9044
rect 18900 8988 19964 9044
rect 20020 8988 20030 9044
rect 35634 8988 35644 9044
rect 35700 8988 36204 9044
rect 36260 8988 37212 9044
rect 37268 8988 37278 9044
rect 43474 8988 43484 9044
rect 43540 8988 47740 9044
rect 47796 8988 47806 9044
rect 48066 8988 48076 9044
rect 48132 8988 48972 9044
rect 49028 8988 49038 9044
rect 53218 8988 53228 9044
rect 53284 8988 54012 9044
rect 54068 8988 54078 9044
rect 47740 8932 47796 8988
rect 62132 8932 62188 9100
rect 62290 8988 62300 9044
rect 62356 8988 63980 9044
rect 64036 8988 64046 9044
rect 69234 8988 69244 9044
rect 69300 8988 69916 9044
rect 69972 8988 70364 9044
rect 70420 8988 70430 9044
rect 27346 8876 27356 8932
rect 27412 8876 29036 8932
rect 29092 8876 29102 8932
rect 47740 8876 49308 8932
rect 49364 8876 49374 8932
rect 50530 8876 50540 8932
rect 50596 8876 51100 8932
rect 51156 8876 51166 8932
rect 58370 8876 58380 8932
rect 58436 8876 60844 8932
rect 60900 8876 62188 8932
rect 66322 8876 66332 8932
rect 66388 8876 67900 8932
rect 67956 8876 67966 8932
rect 0 8820 800 8848
rect 79200 8820 80000 8848
rect 0 8764 1932 8820
rect 1988 8764 1998 8820
rect 7410 8764 7420 8820
rect 7476 8764 9996 8820
rect 10052 8764 20412 8820
rect 20468 8764 20478 8820
rect 77970 8764 77980 8820
rect 78036 8764 80000 8820
rect 0 8736 800 8764
rect 79200 8736 80000 8764
rect 18274 8652 18284 8708
rect 18340 8652 18956 8708
rect 19012 8652 19022 8708
rect 31164 8652 37548 8708
rect 37604 8652 37996 8708
rect 38052 8652 38062 8708
rect 10862 8596 10872 8652
rect 10928 8596 10976 8652
rect 11032 8596 11080 8652
rect 11136 8596 11146 8652
rect 30182 8596 30192 8652
rect 30248 8596 30296 8652
rect 30352 8596 30400 8652
rect 30456 8596 30466 8652
rect 12450 8540 12460 8596
rect 12516 8540 15148 8596
rect 16146 8540 16156 8596
rect 16212 8540 17276 8596
rect 17332 8540 17342 8596
rect 19058 8540 19068 8596
rect 19124 8540 19628 8596
rect 19684 8540 19694 8596
rect 15092 8484 15148 8540
rect 31164 8484 31220 8652
rect 49502 8596 49512 8652
rect 49568 8596 49616 8652
rect 49672 8596 49720 8652
rect 49776 8596 49786 8652
rect 68822 8596 68832 8652
rect 68888 8596 68936 8652
rect 68992 8596 69040 8652
rect 69096 8596 69106 8652
rect 31378 8540 31388 8596
rect 31444 8540 33180 8596
rect 33236 8540 34076 8596
rect 34132 8540 34972 8596
rect 35028 8540 35038 8596
rect 53666 8540 53676 8596
rect 53732 8540 59836 8596
rect 59892 8540 59902 8596
rect 60610 8540 60620 8596
rect 60676 8540 68460 8596
rect 68516 8540 68526 8596
rect 12562 8428 12572 8484
rect 12628 8428 13468 8484
rect 13524 8428 13534 8484
rect 15092 8428 31220 8484
rect 32946 8428 32956 8484
rect 33012 8428 37324 8484
rect 37380 8428 38332 8484
rect 38388 8428 38398 8484
rect 48850 8428 48860 8484
rect 48916 8428 69244 8484
rect 69300 8428 69310 8484
rect 15092 8316 36988 8372
rect 37044 8316 37054 8372
rect 37202 8316 37212 8372
rect 37268 8316 42588 8372
rect 42644 8316 42654 8372
rect 47282 8316 47292 8372
rect 47348 8316 48748 8372
rect 48804 8316 48814 8372
rect 51762 8316 51772 8372
rect 51828 8316 54236 8372
rect 54292 8316 54302 8372
rect 58146 8316 58156 8372
rect 58212 8316 59724 8372
rect 59780 8316 59790 8372
rect 63186 8316 63196 8372
rect 63252 8316 64316 8372
rect 64372 8316 64382 8372
rect 65650 8316 65660 8372
rect 65716 8316 67116 8372
rect 67172 8316 67182 8372
rect 71250 8316 71260 8372
rect 71316 8316 72156 8372
rect 72212 8316 72222 8372
rect 15092 8260 15148 8316
rect 10434 8204 10444 8260
rect 10500 8204 15148 8260
rect 19058 8204 19068 8260
rect 19124 8204 19516 8260
rect 19572 8204 19582 8260
rect 20066 8204 20076 8260
rect 20132 8204 21756 8260
rect 21812 8204 21822 8260
rect 21970 8204 21980 8260
rect 22036 8204 26124 8260
rect 26180 8204 26190 8260
rect 26786 8204 26796 8260
rect 26852 8204 26862 8260
rect 27458 8204 27468 8260
rect 27524 8204 28140 8260
rect 28196 8204 40908 8260
rect 40964 8204 40974 8260
rect 44034 8204 44044 8260
rect 44100 8204 56700 8260
rect 56756 8204 58380 8260
rect 58436 8204 58446 8260
rect 23874 8092 23884 8148
rect 23940 8092 24668 8148
rect 24724 8092 24734 8148
rect 26796 8036 26852 8204
rect 35634 8092 35644 8148
rect 35700 8092 37100 8148
rect 37156 8092 37166 8148
rect 40450 8092 40460 8148
rect 40516 8092 42364 8148
rect 42420 8092 42430 8148
rect 55122 8092 55132 8148
rect 55188 8092 55804 8148
rect 55860 8092 57148 8148
rect 57204 8092 58716 8148
rect 58772 8092 58782 8148
rect 63522 8092 63532 8148
rect 63588 8092 65548 8148
rect 65604 8092 65614 8148
rect 71474 8092 71484 8148
rect 71540 8092 72380 8148
rect 72436 8092 72446 8148
rect 3826 7980 3836 8036
rect 3892 7980 5628 8036
rect 5684 7980 5694 8036
rect 15922 7980 15932 8036
rect 15988 7980 17948 8036
rect 18004 7980 18014 8036
rect 25330 7980 25340 8036
rect 25396 7980 26012 8036
rect 26068 7980 26852 8036
rect 32732 7980 62188 8036
rect 32732 7924 32788 7980
rect 62132 7924 62188 7980
rect 25890 7868 25900 7924
rect 25956 7868 32788 7924
rect 38210 7868 38220 7924
rect 38276 7868 38780 7924
rect 38836 7868 38846 7924
rect 62132 7868 76972 7924
rect 77028 7868 77038 7924
rect 20522 7812 20532 7868
rect 20588 7812 20636 7868
rect 20692 7812 20740 7868
rect 20796 7812 20806 7868
rect 39842 7812 39852 7868
rect 39908 7812 39956 7868
rect 40012 7812 40060 7868
rect 40116 7812 40126 7868
rect 59162 7812 59172 7868
rect 59228 7812 59276 7868
rect 59332 7812 59380 7868
rect 59436 7812 59446 7868
rect 78482 7812 78492 7868
rect 78548 7812 78596 7868
rect 78652 7812 78700 7868
rect 78756 7812 78766 7868
rect 25900 7756 38668 7812
rect 43922 7756 43932 7812
rect 43988 7756 44604 7812
rect 44660 7756 44670 7812
rect 47394 7756 47404 7812
rect 47460 7756 52220 7812
rect 52276 7756 52286 7812
rect 2706 7644 2716 7700
rect 2772 7644 11340 7700
rect 11396 7644 11406 7700
rect 12114 7644 12124 7700
rect 12180 7644 13580 7700
rect 13636 7644 14252 7700
rect 14308 7644 17500 7700
rect 17556 7644 18732 7700
rect 18788 7644 18798 7700
rect 24210 7644 24220 7700
rect 24276 7644 25004 7700
rect 25060 7644 25340 7700
rect 25396 7644 25406 7700
rect 25900 7588 25956 7756
rect 38612 7700 38668 7756
rect 26114 7644 26124 7700
rect 26180 7644 26908 7700
rect 26964 7644 26974 7700
rect 38612 7644 48860 7700
rect 48916 7644 48926 7700
rect 69906 7644 69916 7700
rect 69972 7644 71148 7700
rect 71204 7644 73164 7700
rect 73220 7644 73230 7700
rect 8866 7532 8876 7588
rect 8932 7532 9660 7588
rect 9716 7532 9726 7588
rect 11106 7532 11116 7588
rect 11172 7532 11788 7588
rect 11844 7532 11854 7588
rect 19506 7532 19516 7588
rect 19572 7532 23996 7588
rect 24052 7532 25900 7588
rect 25956 7532 25966 7588
rect 40114 7532 40124 7588
rect 40180 7532 40796 7588
rect 40852 7532 41916 7588
rect 41972 7532 41982 7588
rect 42578 7532 42588 7588
rect 42644 7532 44044 7588
rect 44100 7532 44110 7588
rect 46834 7532 46844 7588
rect 46900 7532 65324 7588
rect 65380 7532 65390 7588
rect 13794 7420 13804 7476
rect 13860 7420 20188 7476
rect 20244 7420 20254 7476
rect 39442 7420 39452 7476
rect 39508 7420 41468 7476
rect 41524 7420 41534 7476
rect 56018 7420 56028 7476
rect 56084 7420 65660 7476
rect 65716 7420 65726 7476
rect 6066 7308 6076 7364
rect 6132 7308 7420 7364
rect 7476 7308 8652 7364
rect 8708 7308 12012 7364
rect 12068 7308 12078 7364
rect 33730 7308 33740 7364
rect 33796 7308 34412 7364
rect 34468 7308 37436 7364
rect 37492 7308 37502 7364
rect 50372 7308 69916 7364
rect 69972 7308 69982 7364
rect 71474 7308 71484 7364
rect 71540 7308 72268 7364
rect 72324 7308 72940 7364
rect 72996 7308 73276 7364
rect 73332 7308 73342 7364
rect 77186 7308 77196 7364
rect 77252 7308 77262 7364
rect 50372 7252 50428 7308
rect 77196 7252 77252 7308
rect 15138 7196 15148 7252
rect 15204 7196 34860 7252
rect 34916 7196 34926 7252
rect 42466 7196 42476 7252
rect 42532 7196 43260 7252
rect 43316 7196 45948 7252
rect 46004 7196 46014 7252
rect 48738 7196 48748 7252
rect 48804 7196 50428 7252
rect 68898 7196 68908 7252
rect 68964 7196 69692 7252
rect 69748 7196 69758 7252
rect 76962 7196 76972 7252
rect 77028 7196 77252 7252
rect 14018 7084 14028 7140
rect 14084 7084 27468 7140
rect 27524 7084 27534 7140
rect 38770 7084 38780 7140
rect 38836 7084 45612 7140
rect 45668 7084 45678 7140
rect 10862 7028 10872 7084
rect 10928 7028 10976 7084
rect 11032 7028 11080 7084
rect 11136 7028 11146 7084
rect 30182 7028 30192 7084
rect 30248 7028 30296 7084
rect 30352 7028 30400 7084
rect 30456 7028 30466 7084
rect 49502 7028 49512 7084
rect 49568 7028 49616 7084
rect 49672 7028 49720 7084
rect 49776 7028 49786 7084
rect 68822 7028 68832 7084
rect 68888 7028 68936 7084
rect 68992 7028 69040 7084
rect 69096 7028 69106 7084
rect 20178 6972 20188 7028
rect 20244 6972 22428 7028
rect 22484 6972 22494 7028
rect 31714 6972 31724 7028
rect 31780 6972 32620 7028
rect 32676 6972 40236 7028
rect 40292 6972 40302 7028
rect 41458 6972 41468 7028
rect 41524 6972 42028 7028
rect 42084 6972 42924 7028
rect 42980 6972 43932 7028
rect 43988 6972 43998 7028
rect 31724 6916 31780 6972
rect 9202 6860 9212 6916
rect 9268 6860 13132 6916
rect 13188 6860 13198 6916
rect 13356 6860 31780 6916
rect 34178 6860 34188 6916
rect 34244 6860 34748 6916
rect 34804 6860 35196 6916
rect 35252 6860 38108 6916
rect 38164 6860 38174 6916
rect 43362 6860 43372 6916
rect 43428 6860 48972 6916
rect 49028 6860 51772 6916
rect 51828 6860 51838 6916
rect 61954 6860 61964 6916
rect 62020 6860 63084 6916
rect 63140 6860 63150 6916
rect 13356 6804 13412 6860
rect 9762 6748 9772 6804
rect 9828 6748 13412 6804
rect 14354 6748 14364 6804
rect 14420 6748 16044 6804
rect 16100 6748 16110 6804
rect 20290 6748 20300 6804
rect 20356 6748 21308 6804
rect 21364 6748 21374 6804
rect 26898 6748 26908 6804
rect 26964 6748 29484 6804
rect 29540 6748 29550 6804
rect 36082 6748 36092 6804
rect 36148 6748 38444 6804
rect 38500 6748 38510 6804
rect 69682 6748 69692 6804
rect 69748 6748 71260 6804
rect 71316 6748 71326 6804
rect 4274 6636 4284 6692
rect 4340 6636 4844 6692
rect 4900 6636 38892 6692
rect 38948 6636 38958 6692
rect 43922 6636 43932 6692
rect 43988 6636 46620 6692
rect 46676 6636 46686 6692
rect 46844 6636 55468 6692
rect 55524 6636 56028 6692
rect 56084 6636 56094 6692
rect 57250 6636 57260 6692
rect 57316 6636 59164 6692
rect 59220 6636 59230 6692
rect 62962 6636 62972 6692
rect 63028 6636 64092 6692
rect 64148 6636 64158 6692
rect 65314 6636 65324 6692
rect 65380 6636 66220 6692
rect 66276 6636 69580 6692
rect 69636 6636 69646 6692
rect 70690 6636 70700 6692
rect 70756 6636 72156 6692
rect 72212 6636 72222 6692
rect 46844 6580 46900 6636
rect 2482 6524 2492 6580
rect 2548 6524 2558 6580
rect 19730 6524 19740 6580
rect 19796 6524 20412 6580
rect 20468 6524 20478 6580
rect 21634 6524 21644 6580
rect 21700 6524 36204 6580
rect 36260 6524 36270 6580
rect 45714 6524 45724 6580
rect 45780 6524 46900 6580
rect 49196 6524 50428 6580
rect 50484 6524 53508 6580
rect 53666 6524 53676 6580
rect 53732 6524 54348 6580
rect 54404 6524 54414 6580
rect 55234 6524 55244 6580
rect 55300 6524 55580 6580
rect 55636 6524 57372 6580
rect 57428 6524 58044 6580
rect 58100 6524 58110 6580
rect 62132 6524 65660 6580
rect 65716 6524 65726 6580
rect 69010 6524 69020 6580
rect 69076 6524 70476 6580
rect 70532 6524 71596 6580
rect 71652 6524 71662 6580
rect 0 6356 800 6384
rect 2492 6356 2548 6524
rect 49196 6468 49252 6524
rect 53452 6468 53508 6524
rect 62132 6468 62188 6524
rect 19170 6412 19180 6468
rect 19236 6412 21028 6468
rect 25330 6412 25340 6468
rect 25396 6412 27020 6468
rect 27076 6412 27468 6468
rect 27524 6412 27534 6468
rect 27906 6412 27916 6468
rect 27972 6412 29372 6468
rect 29428 6412 29438 6468
rect 35074 6412 35084 6468
rect 35140 6412 49196 6468
rect 49252 6412 49262 6468
rect 49420 6412 50876 6468
rect 50932 6412 50942 6468
rect 53452 6412 57148 6468
rect 57204 6412 57214 6468
rect 58258 6412 58268 6468
rect 58324 6412 59724 6468
rect 59780 6412 62188 6468
rect 68674 6412 68684 6468
rect 68740 6412 69356 6468
rect 69412 6412 69422 6468
rect 69794 6412 69804 6468
rect 69860 6412 70924 6468
rect 70980 6412 70990 6468
rect 0 6300 2548 6356
rect 0 6272 800 6300
rect 20522 6244 20532 6300
rect 20588 6244 20636 6300
rect 20692 6244 20740 6300
rect 20796 6244 20806 6300
rect 20972 6244 21028 6412
rect 49420 6356 49476 6412
rect 33282 6300 33292 6356
rect 33348 6300 35644 6356
rect 35700 6300 35710 6356
rect 44258 6300 44268 6356
rect 44324 6300 49476 6356
rect 50876 6356 50932 6412
rect 79200 6356 80000 6384
rect 50876 6300 55692 6356
rect 55748 6300 55758 6356
rect 70242 6300 70252 6356
rect 70308 6300 71708 6356
rect 71764 6300 71774 6356
rect 78876 6300 80000 6356
rect 39842 6244 39852 6300
rect 39908 6244 39956 6300
rect 40012 6244 40060 6300
rect 40116 6244 40126 6300
rect 59162 6244 59172 6300
rect 59228 6244 59276 6300
rect 59332 6244 59380 6300
rect 59436 6244 59446 6300
rect 78482 6244 78492 6300
rect 78548 6244 78596 6300
rect 78652 6244 78700 6300
rect 78756 6244 78766 6300
rect 20972 6188 35868 6244
rect 35924 6188 35934 6244
rect 42802 6188 42812 6244
rect 42868 6188 58268 6244
rect 58324 6188 58334 6244
rect 61730 6188 61740 6244
rect 61796 6188 63252 6244
rect 69570 6188 69580 6244
rect 69636 6188 70028 6244
rect 70084 6188 70588 6244
rect 70644 6188 71372 6244
rect 71428 6188 71438 6244
rect 8978 6076 8988 6132
rect 9044 6076 9996 6132
rect 10052 6076 10062 6132
rect 13122 6076 13132 6132
rect 13188 6076 14252 6132
rect 14308 6076 14318 6132
rect 15810 6076 15820 6132
rect 15876 6076 19740 6132
rect 19796 6076 19806 6132
rect 25106 6076 25116 6132
rect 25172 6076 25676 6132
rect 25732 6076 26012 6132
rect 26068 6076 26572 6132
rect 26628 6076 26638 6132
rect 36194 6076 36204 6132
rect 36260 6076 37100 6132
rect 37156 6076 37166 6132
rect 37426 6076 37436 6132
rect 37492 6076 37996 6132
rect 38052 6076 48748 6132
rect 48804 6076 48814 6132
rect 55346 6076 55356 6132
rect 55412 6076 56028 6132
rect 56084 6076 56588 6132
rect 56644 6076 56654 6132
rect 63196 6020 63252 6188
rect 78876 6132 78932 6300
rect 79200 6272 80000 6300
rect 70690 6076 70700 6132
rect 70756 6076 72940 6132
rect 72996 6076 74172 6132
rect 74228 6076 74238 6132
rect 77970 6076 77980 6132
rect 78036 6076 78932 6132
rect 11106 5964 11116 6020
rect 11172 5964 19964 6020
rect 20020 5964 20412 6020
rect 20468 5964 20478 6020
rect 26852 5964 35756 6020
rect 35812 5964 35822 6020
rect 48178 5964 48188 6020
rect 48244 5964 49532 6020
rect 49588 5964 49598 6020
rect 59938 5964 59948 6020
rect 60004 5964 62188 6020
rect 63186 5964 63196 6020
rect 63252 5964 63262 6020
rect 26852 5908 26908 5964
rect 62132 5908 62188 5964
rect 12674 5852 12684 5908
rect 12740 5852 13580 5908
rect 13636 5852 14588 5908
rect 14644 5852 15148 5908
rect 26338 5852 26348 5908
rect 26404 5852 26908 5908
rect 33618 5852 33628 5908
rect 33684 5852 34300 5908
rect 34356 5852 34366 5908
rect 38994 5852 39004 5908
rect 39060 5852 43036 5908
rect 43092 5852 43102 5908
rect 47842 5852 47852 5908
rect 47908 5852 48860 5908
rect 48916 5852 52668 5908
rect 52724 5852 52734 5908
rect 57474 5852 57484 5908
rect 57540 5852 60508 5908
rect 60564 5852 60574 5908
rect 62132 5852 65436 5908
rect 65492 5852 65884 5908
rect 65940 5852 68684 5908
rect 68740 5852 68750 5908
rect 15092 5796 15148 5852
rect 15092 5740 16716 5796
rect 16772 5740 16782 5796
rect 18386 5740 18396 5796
rect 18452 5740 19292 5796
rect 19348 5740 23548 5796
rect 23604 5740 24220 5796
rect 24276 5740 25004 5796
rect 25060 5740 25070 5796
rect 26674 5740 26684 5796
rect 26740 5740 28140 5796
rect 28196 5740 28206 5796
rect 45826 5740 45836 5796
rect 45892 5740 60620 5796
rect 60676 5740 60844 5796
rect 60900 5740 60910 5796
rect 68450 5740 68460 5796
rect 68516 5740 69356 5796
rect 69412 5740 69422 5796
rect 69906 5740 69916 5796
rect 69972 5740 70924 5796
rect 70980 5740 72268 5796
rect 72324 5740 72334 5796
rect 8978 5628 8988 5684
rect 9044 5628 11564 5684
rect 11620 5628 11630 5684
rect 14242 5628 14252 5684
rect 14308 5628 15148 5684
rect 15204 5628 15214 5684
rect 15698 5628 15708 5684
rect 15764 5628 17500 5684
rect 17556 5628 17566 5684
rect 20738 5628 20748 5684
rect 20804 5628 22428 5684
rect 22484 5628 22494 5684
rect 28466 5628 28476 5684
rect 28532 5628 29484 5684
rect 29540 5628 29550 5684
rect 61628 5628 70588 5684
rect 70644 5628 70654 5684
rect 26226 5516 26236 5572
rect 26292 5516 30100 5572
rect 10862 5460 10872 5516
rect 10928 5460 10976 5516
rect 11032 5460 11080 5516
rect 11136 5460 11146 5516
rect 14690 5404 14700 5460
rect 14756 5404 15036 5460
rect 15092 5404 27916 5460
rect 27972 5404 27982 5460
rect 30044 5348 30100 5516
rect 30182 5460 30192 5516
rect 30248 5460 30296 5516
rect 30352 5460 30400 5516
rect 30456 5460 30466 5516
rect 49502 5460 49512 5516
rect 49568 5460 49616 5516
rect 49672 5460 49720 5516
rect 49776 5460 49786 5516
rect 61628 5460 61684 5628
rect 68822 5460 68832 5516
rect 68888 5460 68936 5516
rect 68992 5460 69040 5516
rect 69096 5460 69106 5516
rect 59826 5404 59836 5460
rect 59892 5404 61628 5460
rect 61684 5404 61694 5460
rect 70802 5404 70812 5460
rect 70868 5404 72380 5460
rect 72436 5404 72446 5460
rect 30044 5292 36204 5348
rect 36260 5292 36652 5348
rect 36708 5292 36718 5348
rect 44818 5292 44828 5348
rect 44884 5292 45276 5348
rect 45332 5292 46508 5348
rect 46564 5292 47068 5348
rect 47124 5292 47134 5348
rect 55346 5292 55356 5348
rect 55412 5292 61404 5348
rect 61460 5292 61470 5348
rect 12898 5180 12908 5236
rect 12964 5180 13916 5236
rect 13972 5180 13982 5236
rect 14466 5180 14476 5236
rect 14532 5180 15148 5236
rect 17938 5180 17948 5236
rect 18004 5180 18956 5236
rect 19012 5180 19022 5236
rect 35634 5180 35644 5236
rect 35700 5180 37436 5236
rect 37492 5180 37502 5236
rect 45714 5180 45724 5236
rect 45780 5180 46620 5236
rect 46676 5180 46686 5236
rect 52994 5180 53004 5236
rect 53060 5180 56028 5236
rect 56084 5180 56094 5236
rect 57138 5180 57148 5236
rect 57204 5180 59388 5236
rect 59444 5180 59454 5236
rect 60722 5180 60732 5236
rect 60788 5180 64988 5236
rect 65044 5180 65660 5236
rect 65716 5180 65726 5236
rect 15092 5124 15148 5180
rect 59388 5124 59444 5180
rect 15092 5068 16268 5124
rect 16324 5068 16334 5124
rect 29698 5068 29708 5124
rect 29764 5068 31948 5124
rect 32004 5068 32014 5124
rect 35410 5068 35420 5124
rect 35476 5068 37100 5124
rect 37156 5068 37166 5124
rect 38210 5068 38220 5124
rect 38276 5068 38668 5124
rect 38724 5068 38734 5124
rect 42690 5068 42700 5124
rect 42756 5068 44940 5124
rect 44996 5068 45006 5124
rect 53554 5068 53564 5124
rect 53620 5068 54236 5124
rect 54292 5068 54302 5124
rect 55682 5068 55692 5124
rect 55748 5068 55916 5124
rect 55972 5068 55982 5124
rect 57810 5068 57820 5124
rect 57876 5068 57886 5124
rect 58146 5068 58156 5124
rect 58212 5068 58828 5124
rect 58884 5068 58894 5124
rect 59388 5068 61180 5124
rect 61236 5068 61246 5124
rect 61394 5068 61404 5124
rect 61460 5068 62972 5124
rect 63028 5068 63868 5124
rect 63924 5068 63934 5124
rect 65762 5068 65772 5124
rect 65828 5068 67228 5124
rect 67284 5068 67294 5124
rect 67890 5068 67900 5124
rect 67956 5068 69020 5124
rect 69076 5068 69086 5124
rect 57820 5012 57876 5068
rect 4386 4956 4396 5012
rect 4452 4956 10612 5012
rect 10770 4956 10780 5012
rect 10836 4956 12796 5012
rect 12852 4956 12862 5012
rect 23202 4956 23212 5012
rect 23268 4956 24556 5012
rect 24612 4956 24622 5012
rect 28690 4956 28700 5012
rect 28756 4956 30268 5012
rect 30324 4956 30334 5012
rect 31602 4956 31612 5012
rect 31668 4956 33292 5012
rect 33348 4956 33358 5012
rect 33516 4956 37772 5012
rect 37828 4956 37838 5012
rect 42354 4956 42364 5012
rect 42420 4956 46060 5012
rect 46116 4956 49868 5012
rect 49924 4956 49934 5012
rect 57820 4956 58716 5012
rect 58772 4956 59500 5012
rect 59556 4956 59566 5012
rect 63298 4956 63308 5012
rect 63364 4956 65548 5012
rect 65604 4956 65614 5012
rect 65986 4956 65996 5012
rect 66052 4956 66332 5012
rect 66388 4956 66398 5012
rect 67106 4956 67116 5012
rect 67172 4956 67676 5012
rect 67732 4956 67742 5012
rect 68562 4956 68572 5012
rect 68628 4956 70364 5012
rect 70420 4956 70430 5012
rect 10556 4900 10612 4956
rect 33516 4900 33572 4956
rect 9202 4844 9212 4900
rect 9268 4844 10332 4900
rect 10388 4844 10398 4900
rect 10556 4844 33572 4900
rect 35634 4844 35644 4900
rect 35700 4844 37660 4900
rect 37716 4844 37726 4900
rect 42914 4844 42924 4900
rect 42980 4844 44380 4900
rect 44436 4844 44446 4900
rect 49186 4844 49196 4900
rect 49252 4844 50652 4900
rect 50708 4844 50718 4900
rect 12450 4732 12460 4788
rect 12516 4732 13692 4788
rect 13748 4732 14476 4788
rect 14532 4732 18508 4788
rect 18564 4732 18574 4788
rect 40450 4732 40460 4788
rect 40516 4732 45052 4788
rect 45108 4732 45118 4788
rect 49410 4732 49420 4788
rect 49476 4732 50428 4788
rect 20522 4676 20532 4732
rect 20588 4676 20636 4732
rect 20692 4676 20740 4732
rect 20796 4676 20806 4732
rect 39842 4676 39852 4732
rect 39908 4676 39956 4732
rect 40012 4676 40060 4732
rect 40116 4676 40126 4732
rect 50372 4676 50428 4732
rect 59162 4676 59172 4732
rect 59228 4676 59276 4732
rect 59332 4676 59380 4732
rect 59436 4676 59446 4732
rect 78482 4676 78492 4732
rect 78548 4676 78596 4732
rect 78652 4676 78700 4732
rect 78756 4676 78766 4732
rect 23538 4620 23548 4676
rect 23604 4620 24444 4676
rect 24500 4620 27020 4676
rect 27076 4620 27804 4676
rect 27860 4620 27870 4676
rect 50372 4620 50652 4676
rect 50708 4620 55356 4676
rect 55412 4620 55422 4676
rect 16594 4508 16604 4564
rect 16660 4508 17612 4564
rect 17668 4508 17678 4564
rect 21746 4508 21756 4564
rect 21812 4508 23324 4564
rect 23380 4508 23390 4564
rect 26852 4508 71036 4564
rect 71092 4508 71102 4564
rect 14690 4396 14700 4452
rect 14756 4396 15372 4452
rect 15428 4396 15438 4452
rect 16706 4396 16716 4452
rect 16772 4396 25788 4452
rect 25844 4396 25854 4452
rect 26852 4340 26908 4508
rect 38658 4396 38668 4452
rect 38724 4396 49420 4452
rect 49476 4396 49486 4452
rect 56914 4396 56924 4452
rect 56980 4396 69692 4452
rect 69748 4396 69758 4452
rect 18722 4284 18732 4340
rect 18788 4284 19404 4340
rect 19460 4284 23884 4340
rect 23940 4284 25452 4340
rect 25508 4284 26908 4340
rect 28018 4284 28028 4340
rect 28084 4284 32284 4340
rect 32340 4284 32350 4340
rect 32498 4284 32508 4340
rect 32564 4284 33628 4340
rect 33684 4284 33694 4340
rect 40338 4284 40348 4340
rect 40404 4284 41020 4340
rect 41076 4284 41086 4340
rect 42018 4284 42028 4340
rect 42084 4284 42812 4340
rect 42868 4284 42878 4340
rect 47954 4284 47964 4340
rect 48020 4284 48860 4340
rect 48916 4284 48926 4340
rect 28028 4228 28084 4284
rect 42028 4228 42084 4284
rect 25778 4172 25788 4228
rect 25844 4172 28084 4228
rect 35298 4172 35308 4228
rect 35364 4172 42084 4228
rect 66322 4172 66332 4228
rect 66388 4172 68124 4228
rect 68180 4172 68190 4228
rect 1922 4060 1932 4116
rect 1988 4060 1998 4116
rect 5730 4060 5740 4116
rect 5796 4060 32788 4116
rect 36418 4060 36428 4116
rect 36484 4060 41916 4116
rect 41972 4060 41982 4116
rect 68226 4060 68236 4116
rect 68292 4060 69468 4116
rect 69524 4060 69534 4116
rect 0 3892 800 3920
rect 1932 3892 1988 4060
rect 32732 4004 32788 4060
rect 32732 3948 40236 4004
rect 40292 3948 40302 4004
rect 10862 3892 10872 3948
rect 10928 3892 10976 3948
rect 11032 3892 11080 3948
rect 11136 3892 11146 3948
rect 30182 3892 30192 3948
rect 30248 3892 30296 3948
rect 30352 3892 30400 3948
rect 30456 3892 30466 3948
rect 49502 3892 49512 3948
rect 49568 3892 49616 3948
rect 49672 3892 49720 3948
rect 49776 3892 49786 3948
rect 68822 3892 68832 3948
rect 68888 3892 68936 3948
rect 68992 3892 69040 3948
rect 69096 3892 69106 3948
rect 79200 3892 80000 3920
rect 0 3836 1988 3892
rect 77970 3836 77980 3892
rect 78036 3836 80000 3892
rect 0 3808 800 3836
rect 79200 3808 80000 3836
rect 4274 3724 4284 3780
rect 4340 3724 5180 3780
rect 5236 3724 38556 3780
rect 38612 3724 38622 3780
rect 42466 3724 42476 3780
rect 42532 3724 68684 3780
rect 68740 3724 68750 3780
rect 15092 3612 20188 3668
rect 20244 3612 20254 3668
rect 55794 3612 55804 3668
rect 55860 3612 57036 3668
rect 57092 3612 57102 3668
rect 62402 3612 62412 3668
rect 62468 3612 64764 3668
rect 64820 3612 64830 3668
rect 4274 3500 4284 3556
rect 4340 3500 5740 3556
rect 5796 3500 5806 3556
rect 15092 3444 15148 3612
rect 19730 3500 19740 3556
rect 19796 3500 20300 3556
rect 20356 3500 20972 3556
rect 21028 3500 21038 3556
rect 38612 3500 44716 3556
rect 44772 3500 44782 3556
rect 72146 3500 72156 3556
rect 72212 3500 72604 3556
rect 72660 3500 72670 3556
rect 38612 3444 38668 3500
rect 8194 3388 8204 3444
rect 8260 3388 15148 3444
rect 32498 3388 32508 3444
rect 32564 3388 38668 3444
rect 44482 3388 44492 3444
rect 44548 3388 47404 3444
rect 47460 3388 47470 3444
rect 48514 3388 48524 3444
rect 48580 3388 51212 3444
rect 51268 3388 51278 3444
rect 19618 3276 19628 3332
rect 19684 3276 77084 3332
rect 77140 3276 77150 3332
rect 20522 3108 20532 3164
rect 20588 3108 20636 3164
rect 20692 3108 20740 3164
rect 20796 3108 20806 3164
rect 39842 3108 39852 3164
rect 39908 3108 39956 3164
rect 40012 3108 40060 3164
rect 40116 3108 40126 3164
rect 59162 3108 59172 3164
rect 59228 3108 59276 3164
rect 59332 3108 59380 3164
rect 59436 3108 59446 3164
rect 78482 3108 78492 3164
rect 78548 3108 78596 3164
rect 78652 3108 78700 3164
rect 78756 3108 78766 3164
rect 11330 2940 11340 2996
rect 11396 2940 45388 2996
rect 45444 2940 45454 2996
rect 32274 2828 32284 2884
rect 32340 2828 67900 2884
rect 67956 2828 67966 2884
rect 15138 2716 15148 2772
rect 15204 2716 45948 2772
rect 46004 2716 46014 2772
rect 29362 2604 29372 2660
rect 29428 2604 69916 2660
rect 69972 2604 69982 2660
rect 24994 2492 25004 2548
rect 25060 2492 71484 2548
rect 71540 2492 71550 2548
rect 6962 2380 6972 2436
rect 7028 2380 35420 2436
rect 35476 2380 35486 2436
rect 1922 1484 1932 1540
rect 1988 1484 1998 1540
rect 0 1428 800 1456
rect 1932 1428 1988 1484
rect 79200 1428 80000 1456
rect 0 1372 1988 1428
rect 75506 1372 75516 1428
rect 75572 1372 80000 1428
rect 0 1344 800 1372
rect 79200 1344 80000 1372
<< via3 >>
rect 10872 36820 10928 36876
rect 10976 36820 11032 36876
rect 11080 36820 11136 36876
rect 30192 36820 30248 36876
rect 30296 36820 30352 36876
rect 30400 36820 30456 36876
rect 49512 36820 49568 36876
rect 49616 36820 49672 36876
rect 49720 36820 49776 36876
rect 68832 36820 68888 36876
rect 68936 36820 68992 36876
rect 69040 36820 69096 36876
rect 20532 36036 20588 36092
rect 20636 36036 20692 36092
rect 20740 36036 20796 36092
rect 39852 36036 39908 36092
rect 39956 36036 40012 36092
rect 40060 36036 40116 36092
rect 59172 36036 59228 36092
rect 59276 36036 59332 36092
rect 59380 36036 59436 36092
rect 78492 36036 78548 36092
rect 78596 36036 78652 36092
rect 78700 36036 78756 36092
rect 10872 35252 10928 35308
rect 10976 35252 11032 35308
rect 11080 35252 11136 35308
rect 30192 35252 30248 35308
rect 30296 35252 30352 35308
rect 30400 35252 30456 35308
rect 49512 35252 49568 35308
rect 49616 35252 49672 35308
rect 49720 35252 49776 35308
rect 68832 35252 68888 35308
rect 68936 35252 68992 35308
rect 69040 35252 69096 35308
rect 20532 34468 20588 34524
rect 20636 34468 20692 34524
rect 20740 34468 20796 34524
rect 39852 34468 39908 34524
rect 39956 34468 40012 34524
rect 40060 34468 40116 34524
rect 59172 34468 59228 34524
rect 59276 34468 59332 34524
rect 59380 34468 59436 34524
rect 78492 34468 78548 34524
rect 78596 34468 78652 34524
rect 78700 34468 78756 34524
rect 10872 33684 10928 33740
rect 10976 33684 11032 33740
rect 11080 33684 11136 33740
rect 30192 33684 30248 33740
rect 30296 33684 30352 33740
rect 30400 33684 30456 33740
rect 49512 33684 49568 33740
rect 49616 33684 49672 33740
rect 49720 33684 49776 33740
rect 68832 33684 68888 33740
rect 68936 33684 68992 33740
rect 69040 33684 69096 33740
rect 20532 32900 20588 32956
rect 20636 32900 20692 32956
rect 20740 32900 20796 32956
rect 39852 32900 39908 32956
rect 39956 32900 40012 32956
rect 40060 32900 40116 32956
rect 59172 32900 59228 32956
rect 59276 32900 59332 32956
rect 59380 32900 59436 32956
rect 78492 32900 78548 32956
rect 78596 32900 78652 32956
rect 78700 32900 78756 32956
rect 10872 32116 10928 32172
rect 10976 32116 11032 32172
rect 11080 32116 11136 32172
rect 30192 32116 30248 32172
rect 30296 32116 30352 32172
rect 30400 32116 30456 32172
rect 49512 32116 49568 32172
rect 49616 32116 49672 32172
rect 49720 32116 49776 32172
rect 68832 32116 68888 32172
rect 68936 32116 68992 32172
rect 69040 32116 69096 32172
rect 20532 31332 20588 31388
rect 20636 31332 20692 31388
rect 20740 31332 20796 31388
rect 39852 31332 39908 31388
rect 39956 31332 40012 31388
rect 40060 31332 40116 31388
rect 59172 31332 59228 31388
rect 59276 31332 59332 31388
rect 59380 31332 59436 31388
rect 78492 31332 78548 31388
rect 78596 31332 78652 31388
rect 78700 31332 78756 31388
rect 10872 30548 10928 30604
rect 10976 30548 11032 30604
rect 11080 30548 11136 30604
rect 30192 30548 30248 30604
rect 30296 30548 30352 30604
rect 30400 30548 30456 30604
rect 49512 30548 49568 30604
rect 49616 30548 49672 30604
rect 49720 30548 49776 30604
rect 68832 30548 68888 30604
rect 68936 30548 68992 30604
rect 69040 30548 69096 30604
rect 20532 29764 20588 29820
rect 20636 29764 20692 29820
rect 20740 29764 20796 29820
rect 39852 29764 39908 29820
rect 39956 29764 40012 29820
rect 40060 29764 40116 29820
rect 59172 29764 59228 29820
rect 59276 29764 59332 29820
rect 59380 29764 59436 29820
rect 78492 29764 78548 29820
rect 78596 29764 78652 29820
rect 78700 29764 78756 29820
rect 10872 28980 10928 29036
rect 10976 28980 11032 29036
rect 11080 28980 11136 29036
rect 30192 28980 30248 29036
rect 30296 28980 30352 29036
rect 30400 28980 30456 29036
rect 49512 28980 49568 29036
rect 49616 28980 49672 29036
rect 49720 28980 49776 29036
rect 68832 28980 68888 29036
rect 68936 28980 68992 29036
rect 69040 28980 69096 29036
rect 20532 28196 20588 28252
rect 20636 28196 20692 28252
rect 20740 28196 20796 28252
rect 39852 28196 39908 28252
rect 39956 28196 40012 28252
rect 40060 28196 40116 28252
rect 59172 28196 59228 28252
rect 59276 28196 59332 28252
rect 59380 28196 59436 28252
rect 78492 28196 78548 28252
rect 78596 28196 78652 28252
rect 78700 28196 78756 28252
rect 10872 27412 10928 27468
rect 10976 27412 11032 27468
rect 11080 27412 11136 27468
rect 30192 27412 30248 27468
rect 30296 27412 30352 27468
rect 30400 27412 30456 27468
rect 49512 27412 49568 27468
rect 49616 27412 49672 27468
rect 49720 27412 49776 27468
rect 68832 27412 68888 27468
rect 68936 27412 68992 27468
rect 69040 27412 69096 27468
rect 20532 26628 20588 26684
rect 20636 26628 20692 26684
rect 20740 26628 20796 26684
rect 39852 26628 39908 26684
rect 39956 26628 40012 26684
rect 40060 26628 40116 26684
rect 59172 26628 59228 26684
rect 59276 26628 59332 26684
rect 59380 26628 59436 26684
rect 78492 26628 78548 26684
rect 78596 26628 78652 26684
rect 78700 26628 78756 26684
rect 10872 25844 10928 25900
rect 10976 25844 11032 25900
rect 11080 25844 11136 25900
rect 30192 25844 30248 25900
rect 30296 25844 30352 25900
rect 30400 25844 30456 25900
rect 49512 25844 49568 25900
rect 49616 25844 49672 25900
rect 49720 25844 49776 25900
rect 68832 25844 68888 25900
rect 68936 25844 68992 25900
rect 69040 25844 69096 25900
rect 20532 25060 20588 25116
rect 20636 25060 20692 25116
rect 20740 25060 20796 25116
rect 39852 25060 39908 25116
rect 39956 25060 40012 25116
rect 40060 25060 40116 25116
rect 59172 25060 59228 25116
rect 59276 25060 59332 25116
rect 59380 25060 59436 25116
rect 78492 25060 78548 25116
rect 78596 25060 78652 25116
rect 78700 25060 78756 25116
rect 10872 24276 10928 24332
rect 10976 24276 11032 24332
rect 11080 24276 11136 24332
rect 30192 24276 30248 24332
rect 30296 24276 30352 24332
rect 30400 24276 30456 24332
rect 49512 24276 49568 24332
rect 49616 24276 49672 24332
rect 49720 24276 49776 24332
rect 68832 24276 68888 24332
rect 68936 24276 68992 24332
rect 69040 24276 69096 24332
rect 20532 23492 20588 23548
rect 20636 23492 20692 23548
rect 20740 23492 20796 23548
rect 39852 23492 39908 23548
rect 39956 23492 40012 23548
rect 40060 23492 40116 23548
rect 59172 23492 59228 23548
rect 59276 23492 59332 23548
rect 59380 23492 59436 23548
rect 78492 23492 78548 23548
rect 78596 23492 78652 23548
rect 78700 23492 78756 23548
rect 10872 22708 10928 22764
rect 10976 22708 11032 22764
rect 11080 22708 11136 22764
rect 30192 22708 30248 22764
rect 30296 22708 30352 22764
rect 30400 22708 30456 22764
rect 49512 22708 49568 22764
rect 49616 22708 49672 22764
rect 49720 22708 49776 22764
rect 68832 22708 68888 22764
rect 68936 22708 68992 22764
rect 69040 22708 69096 22764
rect 20532 21924 20588 21980
rect 20636 21924 20692 21980
rect 20740 21924 20796 21980
rect 39852 21924 39908 21980
rect 39956 21924 40012 21980
rect 40060 21924 40116 21980
rect 59172 21924 59228 21980
rect 59276 21924 59332 21980
rect 59380 21924 59436 21980
rect 78492 21924 78548 21980
rect 78596 21924 78652 21980
rect 78700 21924 78756 21980
rect 10872 21140 10928 21196
rect 10976 21140 11032 21196
rect 11080 21140 11136 21196
rect 30192 21140 30248 21196
rect 30296 21140 30352 21196
rect 30400 21140 30456 21196
rect 49512 21140 49568 21196
rect 49616 21140 49672 21196
rect 49720 21140 49776 21196
rect 68832 21140 68888 21196
rect 68936 21140 68992 21196
rect 69040 21140 69096 21196
rect 20532 20356 20588 20412
rect 20636 20356 20692 20412
rect 20740 20356 20796 20412
rect 39852 20356 39908 20412
rect 39956 20356 40012 20412
rect 40060 20356 40116 20412
rect 59172 20356 59228 20412
rect 59276 20356 59332 20412
rect 59380 20356 59436 20412
rect 78492 20356 78548 20412
rect 78596 20356 78652 20412
rect 78700 20356 78756 20412
rect 10872 19572 10928 19628
rect 10976 19572 11032 19628
rect 11080 19572 11136 19628
rect 30192 19572 30248 19628
rect 30296 19572 30352 19628
rect 30400 19572 30456 19628
rect 49512 19572 49568 19628
rect 49616 19572 49672 19628
rect 49720 19572 49776 19628
rect 68832 19572 68888 19628
rect 68936 19572 68992 19628
rect 69040 19572 69096 19628
rect 20532 18788 20588 18844
rect 20636 18788 20692 18844
rect 20740 18788 20796 18844
rect 39852 18788 39908 18844
rect 39956 18788 40012 18844
rect 40060 18788 40116 18844
rect 59172 18788 59228 18844
rect 59276 18788 59332 18844
rect 59380 18788 59436 18844
rect 78492 18788 78548 18844
rect 78596 18788 78652 18844
rect 78700 18788 78756 18844
rect 10872 18004 10928 18060
rect 10976 18004 11032 18060
rect 11080 18004 11136 18060
rect 30192 18004 30248 18060
rect 30296 18004 30352 18060
rect 30400 18004 30456 18060
rect 49512 18004 49568 18060
rect 49616 18004 49672 18060
rect 49720 18004 49776 18060
rect 68832 18004 68888 18060
rect 68936 18004 68992 18060
rect 69040 18004 69096 18060
rect 20532 17220 20588 17276
rect 20636 17220 20692 17276
rect 20740 17220 20796 17276
rect 39852 17220 39908 17276
rect 39956 17220 40012 17276
rect 40060 17220 40116 17276
rect 59172 17220 59228 17276
rect 59276 17220 59332 17276
rect 59380 17220 59436 17276
rect 78492 17220 78548 17276
rect 78596 17220 78652 17276
rect 78700 17220 78756 17276
rect 10872 16436 10928 16492
rect 10976 16436 11032 16492
rect 11080 16436 11136 16492
rect 30192 16436 30248 16492
rect 30296 16436 30352 16492
rect 30400 16436 30456 16492
rect 49512 16436 49568 16492
rect 49616 16436 49672 16492
rect 49720 16436 49776 16492
rect 68832 16436 68888 16492
rect 68936 16436 68992 16492
rect 69040 16436 69096 16492
rect 20532 15652 20588 15708
rect 20636 15652 20692 15708
rect 20740 15652 20796 15708
rect 39852 15652 39908 15708
rect 39956 15652 40012 15708
rect 40060 15652 40116 15708
rect 59172 15652 59228 15708
rect 59276 15652 59332 15708
rect 59380 15652 59436 15708
rect 78492 15652 78548 15708
rect 78596 15652 78652 15708
rect 78700 15652 78756 15708
rect 10872 14868 10928 14924
rect 10976 14868 11032 14924
rect 11080 14868 11136 14924
rect 30192 14868 30248 14924
rect 30296 14868 30352 14924
rect 30400 14868 30456 14924
rect 49512 14868 49568 14924
rect 49616 14868 49672 14924
rect 49720 14868 49776 14924
rect 68832 14868 68888 14924
rect 68936 14868 68992 14924
rect 69040 14868 69096 14924
rect 20532 14084 20588 14140
rect 20636 14084 20692 14140
rect 20740 14084 20796 14140
rect 39852 14084 39908 14140
rect 39956 14084 40012 14140
rect 40060 14084 40116 14140
rect 59172 14084 59228 14140
rect 59276 14084 59332 14140
rect 59380 14084 59436 14140
rect 78492 14084 78548 14140
rect 78596 14084 78652 14140
rect 78700 14084 78756 14140
rect 10872 13300 10928 13356
rect 10976 13300 11032 13356
rect 11080 13300 11136 13356
rect 30192 13300 30248 13356
rect 30296 13300 30352 13356
rect 30400 13300 30456 13356
rect 49512 13300 49568 13356
rect 49616 13300 49672 13356
rect 49720 13300 49776 13356
rect 68832 13300 68888 13356
rect 68936 13300 68992 13356
rect 69040 13300 69096 13356
rect 20532 12516 20588 12572
rect 20636 12516 20692 12572
rect 20740 12516 20796 12572
rect 39852 12516 39908 12572
rect 39956 12516 40012 12572
rect 40060 12516 40116 12572
rect 59172 12516 59228 12572
rect 59276 12516 59332 12572
rect 59380 12516 59436 12572
rect 78492 12516 78548 12572
rect 78596 12516 78652 12572
rect 78700 12516 78756 12572
rect 10872 11732 10928 11788
rect 10976 11732 11032 11788
rect 11080 11732 11136 11788
rect 30192 11732 30248 11788
rect 30296 11732 30352 11788
rect 30400 11732 30456 11788
rect 49512 11732 49568 11788
rect 49616 11732 49672 11788
rect 49720 11732 49776 11788
rect 68832 11732 68888 11788
rect 68936 11732 68992 11788
rect 69040 11732 69096 11788
rect 20532 10948 20588 11004
rect 20636 10948 20692 11004
rect 20740 10948 20796 11004
rect 39852 10948 39908 11004
rect 39956 10948 40012 11004
rect 40060 10948 40116 11004
rect 59172 10948 59228 11004
rect 59276 10948 59332 11004
rect 59380 10948 59436 11004
rect 78492 10948 78548 11004
rect 78596 10948 78652 11004
rect 78700 10948 78756 11004
rect 10872 10164 10928 10220
rect 10976 10164 11032 10220
rect 11080 10164 11136 10220
rect 30192 10164 30248 10220
rect 30296 10164 30352 10220
rect 30400 10164 30456 10220
rect 49512 10164 49568 10220
rect 49616 10164 49672 10220
rect 49720 10164 49776 10220
rect 68832 10164 68888 10220
rect 68936 10164 68992 10220
rect 69040 10164 69096 10220
rect 20532 9380 20588 9436
rect 20636 9380 20692 9436
rect 20740 9380 20796 9436
rect 39852 9380 39908 9436
rect 39956 9380 40012 9436
rect 40060 9380 40116 9436
rect 59172 9380 59228 9436
rect 59276 9380 59332 9436
rect 59380 9380 59436 9436
rect 78492 9380 78548 9436
rect 78596 9380 78652 9436
rect 78700 9380 78756 9436
rect 10872 8596 10928 8652
rect 10976 8596 11032 8652
rect 11080 8596 11136 8652
rect 30192 8596 30248 8652
rect 30296 8596 30352 8652
rect 30400 8596 30456 8652
rect 49512 8596 49568 8652
rect 49616 8596 49672 8652
rect 49720 8596 49776 8652
rect 68832 8596 68888 8652
rect 68936 8596 68992 8652
rect 69040 8596 69096 8652
rect 20532 7812 20588 7868
rect 20636 7812 20692 7868
rect 20740 7812 20796 7868
rect 39852 7812 39908 7868
rect 39956 7812 40012 7868
rect 40060 7812 40116 7868
rect 59172 7812 59228 7868
rect 59276 7812 59332 7868
rect 59380 7812 59436 7868
rect 78492 7812 78548 7868
rect 78596 7812 78652 7868
rect 78700 7812 78756 7868
rect 10872 7028 10928 7084
rect 10976 7028 11032 7084
rect 11080 7028 11136 7084
rect 30192 7028 30248 7084
rect 30296 7028 30352 7084
rect 30400 7028 30456 7084
rect 49512 7028 49568 7084
rect 49616 7028 49672 7084
rect 49720 7028 49776 7084
rect 68832 7028 68888 7084
rect 68936 7028 68992 7084
rect 69040 7028 69096 7084
rect 20532 6244 20588 6300
rect 20636 6244 20692 6300
rect 20740 6244 20796 6300
rect 39852 6244 39908 6300
rect 39956 6244 40012 6300
rect 40060 6244 40116 6300
rect 59172 6244 59228 6300
rect 59276 6244 59332 6300
rect 59380 6244 59436 6300
rect 78492 6244 78548 6300
rect 78596 6244 78652 6300
rect 78700 6244 78756 6300
rect 10872 5460 10928 5516
rect 10976 5460 11032 5516
rect 11080 5460 11136 5516
rect 30192 5460 30248 5516
rect 30296 5460 30352 5516
rect 30400 5460 30456 5516
rect 49512 5460 49568 5516
rect 49616 5460 49672 5516
rect 49720 5460 49776 5516
rect 68832 5460 68888 5516
rect 68936 5460 68992 5516
rect 69040 5460 69096 5516
rect 20532 4676 20588 4732
rect 20636 4676 20692 4732
rect 20740 4676 20796 4732
rect 39852 4676 39908 4732
rect 39956 4676 40012 4732
rect 40060 4676 40116 4732
rect 59172 4676 59228 4732
rect 59276 4676 59332 4732
rect 59380 4676 59436 4732
rect 78492 4676 78548 4732
rect 78596 4676 78652 4732
rect 78700 4676 78756 4732
rect 10872 3892 10928 3948
rect 10976 3892 11032 3948
rect 11080 3892 11136 3948
rect 30192 3892 30248 3948
rect 30296 3892 30352 3948
rect 30400 3892 30456 3948
rect 49512 3892 49568 3948
rect 49616 3892 49672 3948
rect 49720 3892 49776 3948
rect 68832 3892 68888 3948
rect 68936 3892 68992 3948
rect 69040 3892 69096 3948
rect 20532 3108 20588 3164
rect 20636 3108 20692 3164
rect 20740 3108 20796 3164
rect 39852 3108 39908 3164
rect 39956 3108 40012 3164
rect 40060 3108 40116 3164
rect 59172 3108 59228 3164
rect 59276 3108 59332 3164
rect 59380 3108 59436 3164
rect 78492 3108 78548 3164
rect 78596 3108 78652 3164
rect 78700 3108 78756 3164
<< metal4 >>
rect 10844 36876 11164 36908
rect 10844 36820 10872 36876
rect 10928 36820 10976 36876
rect 11032 36820 11080 36876
rect 11136 36820 11164 36876
rect 10844 35308 11164 36820
rect 10844 35252 10872 35308
rect 10928 35252 10976 35308
rect 11032 35252 11080 35308
rect 11136 35252 11164 35308
rect 10844 33740 11164 35252
rect 10844 33684 10872 33740
rect 10928 33684 10976 33740
rect 11032 33684 11080 33740
rect 11136 33684 11164 33740
rect 10844 32172 11164 33684
rect 10844 32116 10872 32172
rect 10928 32116 10976 32172
rect 11032 32116 11080 32172
rect 11136 32116 11164 32172
rect 10844 30604 11164 32116
rect 10844 30548 10872 30604
rect 10928 30548 10976 30604
rect 11032 30548 11080 30604
rect 11136 30548 11164 30604
rect 10844 29036 11164 30548
rect 10844 28980 10872 29036
rect 10928 28980 10976 29036
rect 11032 28980 11080 29036
rect 11136 28980 11164 29036
rect 10844 27468 11164 28980
rect 10844 27412 10872 27468
rect 10928 27412 10976 27468
rect 11032 27412 11080 27468
rect 11136 27412 11164 27468
rect 10844 25900 11164 27412
rect 10844 25844 10872 25900
rect 10928 25844 10976 25900
rect 11032 25844 11080 25900
rect 11136 25844 11164 25900
rect 10844 24332 11164 25844
rect 10844 24276 10872 24332
rect 10928 24276 10976 24332
rect 11032 24276 11080 24332
rect 11136 24276 11164 24332
rect 10844 22764 11164 24276
rect 10844 22708 10872 22764
rect 10928 22708 10976 22764
rect 11032 22708 11080 22764
rect 11136 22708 11164 22764
rect 10844 21196 11164 22708
rect 10844 21140 10872 21196
rect 10928 21140 10976 21196
rect 11032 21140 11080 21196
rect 11136 21140 11164 21196
rect 10844 19628 11164 21140
rect 10844 19572 10872 19628
rect 10928 19572 10976 19628
rect 11032 19572 11080 19628
rect 11136 19572 11164 19628
rect 10844 18060 11164 19572
rect 10844 18004 10872 18060
rect 10928 18004 10976 18060
rect 11032 18004 11080 18060
rect 11136 18004 11164 18060
rect 10844 16492 11164 18004
rect 10844 16436 10872 16492
rect 10928 16436 10976 16492
rect 11032 16436 11080 16492
rect 11136 16436 11164 16492
rect 10844 14924 11164 16436
rect 10844 14868 10872 14924
rect 10928 14868 10976 14924
rect 11032 14868 11080 14924
rect 11136 14868 11164 14924
rect 10844 13356 11164 14868
rect 10844 13300 10872 13356
rect 10928 13300 10976 13356
rect 11032 13300 11080 13356
rect 11136 13300 11164 13356
rect 10844 11788 11164 13300
rect 10844 11732 10872 11788
rect 10928 11732 10976 11788
rect 11032 11732 11080 11788
rect 11136 11732 11164 11788
rect 10844 10220 11164 11732
rect 10844 10164 10872 10220
rect 10928 10164 10976 10220
rect 11032 10164 11080 10220
rect 11136 10164 11164 10220
rect 10844 8652 11164 10164
rect 10844 8596 10872 8652
rect 10928 8596 10976 8652
rect 11032 8596 11080 8652
rect 11136 8596 11164 8652
rect 10844 7084 11164 8596
rect 10844 7028 10872 7084
rect 10928 7028 10976 7084
rect 11032 7028 11080 7084
rect 11136 7028 11164 7084
rect 10844 5516 11164 7028
rect 10844 5460 10872 5516
rect 10928 5460 10976 5516
rect 11032 5460 11080 5516
rect 11136 5460 11164 5516
rect 10844 3948 11164 5460
rect 10844 3892 10872 3948
rect 10928 3892 10976 3948
rect 11032 3892 11080 3948
rect 11136 3892 11164 3948
rect 10844 3076 11164 3892
rect 20504 36092 20824 36908
rect 20504 36036 20532 36092
rect 20588 36036 20636 36092
rect 20692 36036 20740 36092
rect 20796 36036 20824 36092
rect 20504 34524 20824 36036
rect 20504 34468 20532 34524
rect 20588 34468 20636 34524
rect 20692 34468 20740 34524
rect 20796 34468 20824 34524
rect 20504 32956 20824 34468
rect 20504 32900 20532 32956
rect 20588 32900 20636 32956
rect 20692 32900 20740 32956
rect 20796 32900 20824 32956
rect 20504 31388 20824 32900
rect 20504 31332 20532 31388
rect 20588 31332 20636 31388
rect 20692 31332 20740 31388
rect 20796 31332 20824 31388
rect 20504 29820 20824 31332
rect 20504 29764 20532 29820
rect 20588 29764 20636 29820
rect 20692 29764 20740 29820
rect 20796 29764 20824 29820
rect 20504 28252 20824 29764
rect 20504 28196 20532 28252
rect 20588 28196 20636 28252
rect 20692 28196 20740 28252
rect 20796 28196 20824 28252
rect 20504 26684 20824 28196
rect 20504 26628 20532 26684
rect 20588 26628 20636 26684
rect 20692 26628 20740 26684
rect 20796 26628 20824 26684
rect 20504 25116 20824 26628
rect 20504 25060 20532 25116
rect 20588 25060 20636 25116
rect 20692 25060 20740 25116
rect 20796 25060 20824 25116
rect 20504 23548 20824 25060
rect 20504 23492 20532 23548
rect 20588 23492 20636 23548
rect 20692 23492 20740 23548
rect 20796 23492 20824 23548
rect 20504 21980 20824 23492
rect 20504 21924 20532 21980
rect 20588 21924 20636 21980
rect 20692 21924 20740 21980
rect 20796 21924 20824 21980
rect 20504 20412 20824 21924
rect 20504 20356 20532 20412
rect 20588 20356 20636 20412
rect 20692 20356 20740 20412
rect 20796 20356 20824 20412
rect 20504 18844 20824 20356
rect 20504 18788 20532 18844
rect 20588 18788 20636 18844
rect 20692 18788 20740 18844
rect 20796 18788 20824 18844
rect 20504 17276 20824 18788
rect 20504 17220 20532 17276
rect 20588 17220 20636 17276
rect 20692 17220 20740 17276
rect 20796 17220 20824 17276
rect 20504 15708 20824 17220
rect 20504 15652 20532 15708
rect 20588 15652 20636 15708
rect 20692 15652 20740 15708
rect 20796 15652 20824 15708
rect 20504 14140 20824 15652
rect 20504 14084 20532 14140
rect 20588 14084 20636 14140
rect 20692 14084 20740 14140
rect 20796 14084 20824 14140
rect 20504 12572 20824 14084
rect 20504 12516 20532 12572
rect 20588 12516 20636 12572
rect 20692 12516 20740 12572
rect 20796 12516 20824 12572
rect 20504 11004 20824 12516
rect 20504 10948 20532 11004
rect 20588 10948 20636 11004
rect 20692 10948 20740 11004
rect 20796 10948 20824 11004
rect 20504 9436 20824 10948
rect 20504 9380 20532 9436
rect 20588 9380 20636 9436
rect 20692 9380 20740 9436
rect 20796 9380 20824 9436
rect 20504 7868 20824 9380
rect 20504 7812 20532 7868
rect 20588 7812 20636 7868
rect 20692 7812 20740 7868
rect 20796 7812 20824 7868
rect 20504 6300 20824 7812
rect 20504 6244 20532 6300
rect 20588 6244 20636 6300
rect 20692 6244 20740 6300
rect 20796 6244 20824 6300
rect 20504 4732 20824 6244
rect 20504 4676 20532 4732
rect 20588 4676 20636 4732
rect 20692 4676 20740 4732
rect 20796 4676 20824 4732
rect 20504 3164 20824 4676
rect 20504 3108 20532 3164
rect 20588 3108 20636 3164
rect 20692 3108 20740 3164
rect 20796 3108 20824 3164
rect 20504 3076 20824 3108
rect 30164 36876 30484 36908
rect 30164 36820 30192 36876
rect 30248 36820 30296 36876
rect 30352 36820 30400 36876
rect 30456 36820 30484 36876
rect 30164 35308 30484 36820
rect 30164 35252 30192 35308
rect 30248 35252 30296 35308
rect 30352 35252 30400 35308
rect 30456 35252 30484 35308
rect 30164 33740 30484 35252
rect 30164 33684 30192 33740
rect 30248 33684 30296 33740
rect 30352 33684 30400 33740
rect 30456 33684 30484 33740
rect 30164 32172 30484 33684
rect 30164 32116 30192 32172
rect 30248 32116 30296 32172
rect 30352 32116 30400 32172
rect 30456 32116 30484 32172
rect 30164 30604 30484 32116
rect 30164 30548 30192 30604
rect 30248 30548 30296 30604
rect 30352 30548 30400 30604
rect 30456 30548 30484 30604
rect 30164 29036 30484 30548
rect 30164 28980 30192 29036
rect 30248 28980 30296 29036
rect 30352 28980 30400 29036
rect 30456 28980 30484 29036
rect 30164 27468 30484 28980
rect 30164 27412 30192 27468
rect 30248 27412 30296 27468
rect 30352 27412 30400 27468
rect 30456 27412 30484 27468
rect 30164 25900 30484 27412
rect 30164 25844 30192 25900
rect 30248 25844 30296 25900
rect 30352 25844 30400 25900
rect 30456 25844 30484 25900
rect 30164 24332 30484 25844
rect 30164 24276 30192 24332
rect 30248 24276 30296 24332
rect 30352 24276 30400 24332
rect 30456 24276 30484 24332
rect 30164 22764 30484 24276
rect 30164 22708 30192 22764
rect 30248 22708 30296 22764
rect 30352 22708 30400 22764
rect 30456 22708 30484 22764
rect 30164 21196 30484 22708
rect 30164 21140 30192 21196
rect 30248 21140 30296 21196
rect 30352 21140 30400 21196
rect 30456 21140 30484 21196
rect 30164 19628 30484 21140
rect 30164 19572 30192 19628
rect 30248 19572 30296 19628
rect 30352 19572 30400 19628
rect 30456 19572 30484 19628
rect 30164 18060 30484 19572
rect 30164 18004 30192 18060
rect 30248 18004 30296 18060
rect 30352 18004 30400 18060
rect 30456 18004 30484 18060
rect 30164 16492 30484 18004
rect 30164 16436 30192 16492
rect 30248 16436 30296 16492
rect 30352 16436 30400 16492
rect 30456 16436 30484 16492
rect 30164 14924 30484 16436
rect 30164 14868 30192 14924
rect 30248 14868 30296 14924
rect 30352 14868 30400 14924
rect 30456 14868 30484 14924
rect 30164 13356 30484 14868
rect 30164 13300 30192 13356
rect 30248 13300 30296 13356
rect 30352 13300 30400 13356
rect 30456 13300 30484 13356
rect 30164 11788 30484 13300
rect 30164 11732 30192 11788
rect 30248 11732 30296 11788
rect 30352 11732 30400 11788
rect 30456 11732 30484 11788
rect 30164 10220 30484 11732
rect 30164 10164 30192 10220
rect 30248 10164 30296 10220
rect 30352 10164 30400 10220
rect 30456 10164 30484 10220
rect 30164 8652 30484 10164
rect 30164 8596 30192 8652
rect 30248 8596 30296 8652
rect 30352 8596 30400 8652
rect 30456 8596 30484 8652
rect 30164 7084 30484 8596
rect 30164 7028 30192 7084
rect 30248 7028 30296 7084
rect 30352 7028 30400 7084
rect 30456 7028 30484 7084
rect 30164 5516 30484 7028
rect 30164 5460 30192 5516
rect 30248 5460 30296 5516
rect 30352 5460 30400 5516
rect 30456 5460 30484 5516
rect 30164 3948 30484 5460
rect 30164 3892 30192 3948
rect 30248 3892 30296 3948
rect 30352 3892 30400 3948
rect 30456 3892 30484 3948
rect 30164 3076 30484 3892
rect 39824 36092 40144 36908
rect 39824 36036 39852 36092
rect 39908 36036 39956 36092
rect 40012 36036 40060 36092
rect 40116 36036 40144 36092
rect 39824 34524 40144 36036
rect 39824 34468 39852 34524
rect 39908 34468 39956 34524
rect 40012 34468 40060 34524
rect 40116 34468 40144 34524
rect 39824 32956 40144 34468
rect 39824 32900 39852 32956
rect 39908 32900 39956 32956
rect 40012 32900 40060 32956
rect 40116 32900 40144 32956
rect 39824 31388 40144 32900
rect 39824 31332 39852 31388
rect 39908 31332 39956 31388
rect 40012 31332 40060 31388
rect 40116 31332 40144 31388
rect 39824 29820 40144 31332
rect 39824 29764 39852 29820
rect 39908 29764 39956 29820
rect 40012 29764 40060 29820
rect 40116 29764 40144 29820
rect 39824 28252 40144 29764
rect 39824 28196 39852 28252
rect 39908 28196 39956 28252
rect 40012 28196 40060 28252
rect 40116 28196 40144 28252
rect 39824 26684 40144 28196
rect 39824 26628 39852 26684
rect 39908 26628 39956 26684
rect 40012 26628 40060 26684
rect 40116 26628 40144 26684
rect 39824 25116 40144 26628
rect 39824 25060 39852 25116
rect 39908 25060 39956 25116
rect 40012 25060 40060 25116
rect 40116 25060 40144 25116
rect 39824 23548 40144 25060
rect 39824 23492 39852 23548
rect 39908 23492 39956 23548
rect 40012 23492 40060 23548
rect 40116 23492 40144 23548
rect 39824 21980 40144 23492
rect 39824 21924 39852 21980
rect 39908 21924 39956 21980
rect 40012 21924 40060 21980
rect 40116 21924 40144 21980
rect 39824 20412 40144 21924
rect 39824 20356 39852 20412
rect 39908 20356 39956 20412
rect 40012 20356 40060 20412
rect 40116 20356 40144 20412
rect 39824 18844 40144 20356
rect 39824 18788 39852 18844
rect 39908 18788 39956 18844
rect 40012 18788 40060 18844
rect 40116 18788 40144 18844
rect 39824 17276 40144 18788
rect 39824 17220 39852 17276
rect 39908 17220 39956 17276
rect 40012 17220 40060 17276
rect 40116 17220 40144 17276
rect 39824 15708 40144 17220
rect 39824 15652 39852 15708
rect 39908 15652 39956 15708
rect 40012 15652 40060 15708
rect 40116 15652 40144 15708
rect 39824 14140 40144 15652
rect 39824 14084 39852 14140
rect 39908 14084 39956 14140
rect 40012 14084 40060 14140
rect 40116 14084 40144 14140
rect 39824 12572 40144 14084
rect 39824 12516 39852 12572
rect 39908 12516 39956 12572
rect 40012 12516 40060 12572
rect 40116 12516 40144 12572
rect 39824 11004 40144 12516
rect 39824 10948 39852 11004
rect 39908 10948 39956 11004
rect 40012 10948 40060 11004
rect 40116 10948 40144 11004
rect 39824 9436 40144 10948
rect 39824 9380 39852 9436
rect 39908 9380 39956 9436
rect 40012 9380 40060 9436
rect 40116 9380 40144 9436
rect 39824 7868 40144 9380
rect 39824 7812 39852 7868
rect 39908 7812 39956 7868
rect 40012 7812 40060 7868
rect 40116 7812 40144 7868
rect 39824 6300 40144 7812
rect 39824 6244 39852 6300
rect 39908 6244 39956 6300
rect 40012 6244 40060 6300
rect 40116 6244 40144 6300
rect 39824 4732 40144 6244
rect 39824 4676 39852 4732
rect 39908 4676 39956 4732
rect 40012 4676 40060 4732
rect 40116 4676 40144 4732
rect 39824 3164 40144 4676
rect 39824 3108 39852 3164
rect 39908 3108 39956 3164
rect 40012 3108 40060 3164
rect 40116 3108 40144 3164
rect 39824 3076 40144 3108
rect 49484 36876 49804 36908
rect 49484 36820 49512 36876
rect 49568 36820 49616 36876
rect 49672 36820 49720 36876
rect 49776 36820 49804 36876
rect 49484 35308 49804 36820
rect 49484 35252 49512 35308
rect 49568 35252 49616 35308
rect 49672 35252 49720 35308
rect 49776 35252 49804 35308
rect 49484 33740 49804 35252
rect 49484 33684 49512 33740
rect 49568 33684 49616 33740
rect 49672 33684 49720 33740
rect 49776 33684 49804 33740
rect 49484 32172 49804 33684
rect 49484 32116 49512 32172
rect 49568 32116 49616 32172
rect 49672 32116 49720 32172
rect 49776 32116 49804 32172
rect 49484 30604 49804 32116
rect 49484 30548 49512 30604
rect 49568 30548 49616 30604
rect 49672 30548 49720 30604
rect 49776 30548 49804 30604
rect 49484 29036 49804 30548
rect 49484 28980 49512 29036
rect 49568 28980 49616 29036
rect 49672 28980 49720 29036
rect 49776 28980 49804 29036
rect 49484 27468 49804 28980
rect 49484 27412 49512 27468
rect 49568 27412 49616 27468
rect 49672 27412 49720 27468
rect 49776 27412 49804 27468
rect 49484 25900 49804 27412
rect 49484 25844 49512 25900
rect 49568 25844 49616 25900
rect 49672 25844 49720 25900
rect 49776 25844 49804 25900
rect 49484 24332 49804 25844
rect 49484 24276 49512 24332
rect 49568 24276 49616 24332
rect 49672 24276 49720 24332
rect 49776 24276 49804 24332
rect 49484 22764 49804 24276
rect 49484 22708 49512 22764
rect 49568 22708 49616 22764
rect 49672 22708 49720 22764
rect 49776 22708 49804 22764
rect 49484 21196 49804 22708
rect 49484 21140 49512 21196
rect 49568 21140 49616 21196
rect 49672 21140 49720 21196
rect 49776 21140 49804 21196
rect 49484 19628 49804 21140
rect 49484 19572 49512 19628
rect 49568 19572 49616 19628
rect 49672 19572 49720 19628
rect 49776 19572 49804 19628
rect 49484 18060 49804 19572
rect 49484 18004 49512 18060
rect 49568 18004 49616 18060
rect 49672 18004 49720 18060
rect 49776 18004 49804 18060
rect 49484 16492 49804 18004
rect 49484 16436 49512 16492
rect 49568 16436 49616 16492
rect 49672 16436 49720 16492
rect 49776 16436 49804 16492
rect 49484 14924 49804 16436
rect 49484 14868 49512 14924
rect 49568 14868 49616 14924
rect 49672 14868 49720 14924
rect 49776 14868 49804 14924
rect 49484 13356 49804 14868
rect 49484 13300 49512 13356
rect 49568 13300 49616 13356
rect 49672 13300 49720 13356
rect 49776 13300 49804 13356
rect 49484 11788 49804 13300
rect 49484 11732 49512 11788
rect 49568 11732 49616 11788
rect 49672 11732 49720 11788
rect 49776 11732 49804 11788
rect 49484 10220 49804 11732
rect 49484 10164 49512 10220
rect 49568 10164 49616 10220
rect 49672 10164 49720 10220
rect 49776 10164 49804 10220
rect 49484 8652 49804 10164
rect 49484 8596 49512 8652
rect 49568 8596 49616 8652
rect 49672 8596 49720 8652
rect 49776 8596 49804 8652
rect 49484 7084 49804 8596
rect 49484 7028 49512 7084
rect 49568 7028 49616 7084
rect 49672 7028 49720 7084
rect 49776 7028 49804 7084
rect 49484 5516 49804 7028
rect 49484 5460 49512 5516
rect 49568 5460 49616 5516
rect 49672 5460 49720 5516
rect 49776 5460 49804 5516
rect 49484 3948 49804 5460
rect 49484 3892 49512 3948
rect 49568 3892 49616 3948
rect 49672 3892 49720 3948
rect 49776 3892 49804 3948
rect 49484 3076 49804 3892
rect 59144 36092 59464 36908
rect 59144 36036 59172 36092
rect 59228 36036 59276 36092
rect 59332 36036 59380 36092
rect 59436 36036 59464 36092
rect 59144 34524 59464 36036
rect 59144 34468 59172 34524
rect 59228 34468 59276 34524
rect 59332 34468 59380 34524
rect 59436 34468 59464 34524
rect 59144 32956 59464 34468
rect 59144 32900 59172 32956
rect 59228 32900 59276 32956
rect 59332 32900 59380 32956
rect 59436 32900 59464 32956
rect 59144 31388 59464 32900
rect 59144 31332 59172 31388
rect 59228 31332 59276 31388
rect 59332 31332 59380 31388
rect 59436 31332 59464 31388
rect 59144 29820 59464 31332
rect 59144 29764 59172 29820
rect 59228 29764 59276 29820
rect 59332 29764 59380 29820
rect 59436 29764 59464 29820
rect 59144 28252 59464 29764
rect 59144 28196 59172 28252
rect 59228 28196 59276 28252
rect 59332 28196 59380 28252
rect 59436 28196 59464 28252
rect 59144 26684 59464 28196
rect 59144 26628 59172 26684
rect 59228 26628 59276 26684
rect 59332 26628 59380 26684
rect 59436 26628 59464 26684
rect 59144 25116 59464 26628
rect 59144 25060 59172 25116
rect 59228 25060 59276 25116
rect 59332 25060 59380 25116
rect 59436 25060 59464 25116
rect 59144 23548 59464 25060
rect 59144 23492 59172 23548
rect 59228 23492 59276 23548
rect 59332 23492 59380 23548
rect 59436 23492 59464 23548
rect 59144 21980 59464 23492
rect 59144 21924 59172 21980
rect 59228 21924 59276 21980
rect 59332 21924 59380 21980
rect 59436 21924 59464 21980
rect 59144 20412 59464 21924
rect 59144 20356 59172 20412
rect 59228 20356 59276 20412
rect 59332 20356 59380 20412
rect 59436 20356 59464 20412
rect 59144 18844 59464 20356
rect 59144 18788 59172 18844
rect 59228 18788 59276 18844
rect 59332 18788 59380 18844
rect 59436 18788 59464 18844
rect 59144 17276 59464 18788
rect 59144 17220 59172 17276
rect 59228 17220 59276 17276
rect 59332 17220 59380 17276
rect 59436 17220 59464 17276
rect 59144 15708 59464 17220
rect 59144 15652 59172 15708
rect 59228 15652 59276 15708
rect 59332 15652 59380 15708
rect 59436 15652 59464 15708
rect 59144 14140 59464 15652
rect 59144 14084 59172 14140
rect 59228 14084 59276 14140
rect 59332 14084 59380 14140
rect 59436 14084 59464 14140
rect 59144 12572 59464 14084
rect 59144 12516 59172 12572
rect 59228 12516 59276 12572
rect 59332 12516 59380 12572
rect 59436 12516 59464 12572
rect 59144 11004 59464 12516
rect 59144 10948 59172 11004
rect 59228 10948 59276 11004
rect 59332 10948 59380 11004
rect 59436 10948 59464 11004
rect 59144 9436 59464 10948
rect 59144 9380 59172 9436
rect 59228 9380 59276 9436
rect 59332 9380 59380 9436
rect 59436 9380 59464 9436
rect 59144 7868 59464 9380
rect 59144 7812 59172 7868
rect 59228 7812 59276 7868
rect 59332 7812 59380 7868
rect 59436 7812 59464 7868
rect 59144 6300 59464 7812
rect 59144 6244 59172 6300
rect 59228 6244 59276 6300
rect 59332 6244 59380 6300
rect 59436 6244 59464 6300
rect 59144 4732 59464 6244
rect 59144 4676 59172 4732
rect 59228 4676 59276 4732
rect 59332 4676 59380 4732
rect 59436 4676 59464 4732
rect 59144 3164 59464 4676
rect 59144 3108 59172 3164
rect 59228 3108 59276 3164
rect 59332 3108 59380 3164
rect 59436 3108 59464 3164
rect 59144 3076 59464 3108
rect 68804 36876 69124 36908
rect 68804 36820 68832 36876
rect 68888 36820 68936 36876
rect 68992 36820 69040 36876
rect 69096 36820 69124 36876
rect 68804 35308 69124 36820
rect 68804 35252 68832 35308
rect 68888 35252 68936 35308
rect 68992 35252 69040 35308
rect 69096 35252 69124 35308
rect 68804 33740 69124 35252
rect 68804 33684 68832 33740
rect 68888 33684 68936 33740
rect 68992 33684 69040 33740
rect 69096 33684 69124 33740
rect 68804 32172 69124 33684
rect 68804 32116 68832 32172
rect 68888 32116 68936 32172
rect 68992 32116 69040 32172
rect 69096 32116 69124 32172
rect 68804 30604 69124 32116
rect 68804 30548 68832 30604
rect 68888 30548 68936 30604
rect 68992 30548 69040 30604
rect 69096 30548 69124 30604
rect 68804 29036 69124 30548
rect 68804 28980 68832 29036
rect 68888 28980 68936 29036
rect 68992 28980 69040 29036
rect 69096 28980 69124 29036
rect 68804 27468 69124 28980
rect 68804 27412 68832 27468
rect 68888 27412 68936 27468
rect 68992 27412 69040 27468
rect 69096 27412 69124 27468
rect 68804 25900 69124 27412
rect 68804 25844 68832 25900
rect 68888 25844 68936 25900
rect 68992 25844 69040 25900
rect 69096 25844 69124 25900
rect 68804 24332 69124 25844
rect 68804 24276 68832 24332
rect 68888 24276 68936 24332
rect 68992 24276 69040 24332
rect 69096 24276 69124 24332
rect 68804 22764 69124 24276
rect 68804 22708 68832 22764
rect 68888 22708 68936 22764
rect 68992 22708 69040 22764
rect 69096 22708 69124 22764
rect 68804 21196 69124 22708
rect 68804 21140 68832 21196
rect 68888 21140 68936 21196
rect 68992 21140 69040 21196
rect 69096 21140 69124 21196
rect 68804 19628 69124 21140
rect 68804 19572 68832 19628
rect 68888 19572 68936 19628
rect 68992 19572 69040 19628
rect 69096 19572 69124 19628
rect 68804 18060 69124 19572
rect 68804 18004 68832 18060
rect 68888 18004 68936 18060
rect 68992 18004 69040 18060
rect 69096 18004 69124 18060
rect 68804 16492 69124 18004
rect 68804 16436 68832 16492
rect 68888 16436 68936 16492
rect 68992 16436 69040 16492
rect 69096 16436 69124 16492
rect 68804 14924 69124 16436
rect 68804 14868 68832 14924
rect 68888 14868 68936 14924
rect 68992 14868 69040 14924
rect 69096 14868 69124 14924
rect 68804 13356 69124 14868
rect 68804 13300 68832 13356
rect 68888 13300 68936 13356
rect 68992 13300 69040 13356
rect 69096 13300 69124 13356
rect 68804 11788 69124 13300
rect 68804 11732 68832 11788
rect 68888 11732 68936 11788
rect 68992 11732 69040 11788
rect 69096 11732 69124 11788
rect 68804 10220 69124 11732
rect 68804 10164 68832 10220
rect 68888 10164 68936 10220
rect 68992 10164 69040 10220
rect 69096 10164 69124 10220
rect 68804 8652 69124 10164
rect 68804 8596 68832 8652
rect 68888 8596 68936 8652
rect 68992 8596 69040 8652
rect 69096 8596 69124 8652
rect 68804 7084 69124 8596
rect 68804 7028 68832 7084
rect 68888 7028 68936 7084
rect 68992 7028 69040 7084
rect 69096 7028 69124 7084
rect 68804 5516 69124 7028
rect 68804 5460 68832 5516
rect 68888 5460 68936 5516
rect 68992 5460 69040 5516
rect 69096 5460 69124 5516
rect 68804 3948 69124 5460
rect 68804 3892 68832 3948
rect 68888 3892 68936 3948
rect 68992 3892 69040 3948
rect 69096 3892 69124 3948
rect 68804 3076 69124 3892
rect 78464 36092 78784 36908
rect 78464 36036 78492 36092
rect 78548 36036 78596 36092
rect 78652 36036 78700 36092
rect 78756 36036 78784 36092
rect 78464 34524 78784 36036
rect 78464 34468 78492 34524
rect 78548 34468 78596 34524
rect 78652 34468 78700 34524
rect 78756 34468 78784 34524
rect 78464 32956 78784 34468
rect 78464 32900 78492 32956
rect 78548 32900 78596 32956
rect 78652 32900 78700 32956
rect 78756 32900 78784 32956
rect 78464 31388 78784 32900
rect 78464 31332 78492 31388
rect 78548 31332 78596 31388
rect 78652 31332 78700 31388
rect 78756 31332 78784 31388
rect 78464 29820 78784 31332
rect 78464 29764 78492 29820
rect 78548 29764 78596 29820
rect 78652 29764 78700 29820
rect 78756 29764 78784 29820
rect 78464 28252 78784 29764
rect 78464 28196 78492 28252
rect 78548 28196 78596 28252
rect 78652 28196 78700 28252
rect 78756 28196 78784 28252
rect 78464 26684 78784 28196
rect 78464 26628 78492 26684
rect 78548 26628 78596 26684
rect 78652 26628 78700 26684
rect 78756 26628 78784 26684
rect 78464 25116 78784 26628
rect 78464 25060 78492 25116
rect 78548 25060 78596 25116
rect 78652 25060 78700 25116
rect 78756 25060 78784 25116
rect 78464 23548 78784 25060
rect 78464 23492 78492 23548
rect 78548 23492 78596 23548
rect 78652 23492 78700 23548
rect 78756 23492 78784 23548
rect 78464 21980 78784 23492
rect 78464 21924 78492 21980
rect 78548 21924 78596 21980
rect 78652 21924 78700 21980
rect 78756 21924 78784 21980
rect 78464 20412 78784 21924
rect 78464 20356 78492 20412
rect 78548 20356 78596 20412
rect 78652 20356 78700 20412
rect 78756 20356 78784 20412
rect 78464 18844 78784 20356
rect 78464 18788 78492 18844
rect 78548 18788 78596 18844
rect 78652 18788 78700 18844
rect 78756 18788 78784 18844
rect 78464 17276 78784 18788
rect 78464 17220 78492 17276
rect 78548 17220 78596 17276
rect 78652 17220 78700 17276
rect 78756 17220 78784 17276
rect 78464 15708 78784 17220
rect 78464 15652 78492 15708
rect 78548 15652 78596 15708
rect 78652 15652 78700 15708
rect 78756 15652 78784 15708
rect 78464 14140 78784 15652
rect 78464 14084 78492 14140
rect 78548 14084 78596 14140
rect 78652 14084 78700 14140
rect 78756 14084 78784 14140
rect 78464 12572 78784 14084
rect 78464 12516 78492 12572
rect 78548 12516 78596 12572
rect 78652 12516 78700 12572
rect 78756 12516 78784 12572
rect 78464 11004 78784 12516
rect 78464 10948 78492 11004
rect 78548 10948 78596 11004
rect 78652 10948 78700 11004
rect 78756 10948 78784 11004
rect 78464 9436 78784 10948
rect 78464 9380 78492 9436
rect 78548 9380 78596 9436
rect 78652 9380 78700 9436
rect 78756 9380 78784 9436
rect 78464 7868 78784 9380
rect 78464 7812 78492 7868
rect 78548 7812 78596 7868
rect 78652 7812 78700 7868
rect 78756 7812 78784 7868
rect 78464 6300 78784 7812
rect 78464 6244 78492 6300
rect 78548 6244 78596 6300
rect 78652 6244 78700 6300
rect 78756 6244 78784 6300
rect 78464 4732 78784 6244
rect 78464 4676 78492 4732
rect 78548 4676 78596 4732
rect 78652 4676 78700 4732
rect 78756 4676 78784 4732
rect 78464 3164 78784 4676
rect 78464 3108 78492 3164
rect 78548 3108 78596 3164
rect 78652 3108 78700 3164
rect 78756 3108 78784 3164
rect 78464 3076 78784 3108
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1045_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27216 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1046_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1047_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 33040 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1048_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 34496 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1049_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37184 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1050_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16576 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1051_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 32032 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1052_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25872 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1053_
timestamp 1698175906
transform 1 0 29232 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1054_
timestamp 1698175906
transform 1 0 33376 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1055_
timestamp 1698175906
transform -1 0 43232 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1056_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1057_
timestamp 1698175906
transform 1 0 36400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1058_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 30912 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1059_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27664 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1060_
timestamp 1698175906
transform 1 0 36960 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1061_
timestamp 1698175906
transform 1 0 37072 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1062_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 34944 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1063_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 32368 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1064_
timestamp 1698175906
transform -1 0 27216 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1065_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1066_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 33600 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1067_
timestamp 1698175906
transform 1 0 41664 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1068_
timestamp 1698175906
transform 1 0 40432 0 1 17248
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1069_
timestamp 1698175906
transform -1 0 35168 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1070_
timestamp 1698175906
transform -1 0 37072 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1071_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 40432 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1072_
timestamp 1698175906
transform -1 0 27440 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1073_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 36624 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1074_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 43344 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1075_
timestamp 1698175906
transform -1 0 21840 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1076_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 36400 0 1 17248
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1077_
timestamp 1698175906
transform -1 0 29008 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1078_
timestamp 1698175906
transform -1 0 24528 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1079_
timestamp 1698175906
transform -1 0 16800 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1080_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 10976
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1081_
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1082_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 35392 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1083_
timestamp 1698175906
transform -1 0 36400 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1084_
timestamp 1698175906
transform -1 0 41328 0 1 18816
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1085_
timestamp 1698175906
transform -1 0 38080 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1086_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 35168 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1087_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 28336 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1088_
timestamp 1698175906
transform -1 0 14896 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1089_
timestamp 1698175906
transform -1 0 37296 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1090_
timestamp 1698175906
transform -1 0 40208 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1091_
timestamp 1698175906
transform 1 0 33936 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1092_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 34160 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1093_
timestamp 1698175906
transform -1 0 34496 0 1 17248
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1094_
timestamp 1698175906
transform -1 0 30576 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1095_
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1096_
timestamp 1698175906
transform -1 0 14448 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1097_
timestamp 1698175906
transform 1 0 11648 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1098_
timestamp 1698175906
transform 1 0 24416 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1099_
timestamp 1698175906
transform -1 0 29904 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14784 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12208 0 -1 12544
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1102_
timestamp 1698175906
transform -1 0 28112 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1103_
timestamp 1698175906
transform 1 0 17920 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1104_
timestamp 1698175906
transform -1 0 20384 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1105_
timestamp 1698175906
transform 1 0 17136 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18704 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1108_
timestamp 1698175906
transform -1 0 77952 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1109_
timestamp 1698175906
transform 1 0 53760 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1110_
timestamp 1698175906
transform 1 0 52752 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1111_
timestamp 1698175906
transform 1 0 55328 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1112_
timestamp 1698175906
transform 1 0 54320 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1113_
timestamp 1698175906
transform 1 0 54880 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1114_
timestamp 1698175906
transform -1 0 25424 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1115_
timestamp 1698175906
transform 1 0 52864 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1116_
timestamp 1698175906
transform 1 0 53424 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1117_
timestamp 1698175906
transform 1 0 52864 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1118_
timestamp 1698175906
transform 1 0 53424 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1119_
timestamp 1698175906
transform 1 0 56448 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1120_
timestamp 1698175906
transform -1 0 28448 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16688 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1122_
timestamp 1698175906
transform -1 0 56224 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1123_
timestamp 1698175906
transform -1 0 14000 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1124_
timestamp 1698175906
transform 1 0 54208 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1125_
timestamp 1698175906
transform -1 0 12768 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1126_
timestamp 1698175906
transform 1 0 54320 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1127_
timestamp 1698175906
transform -1 0 12432 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _1128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11536 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1129_
timestamp 1698175906
transform 1 0 56448 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1130_
timestamp 1698175906
transform 1 0 56448 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1131_
timestamp 1698175906
transform -1 0 20832 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1132_
timestamp 1698175906
transform -1 0 60032 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1133_
timestamp 1698175906
transform -1 0 19488 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1134_
timestamp 1698175906
transform -1 0 18256 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15568 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1136_
timestamp 1698175906
transform 1 0 25760 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1137_
timestamp 1698175906
transform -1 0 27216 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1138_
timestamp 1698175906
transform -1 0 27328 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1139_
timestamp 1698175906
transform 1 0 30240 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28672 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1141_
timestamp 1698175906
transform -1 0 26432 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1142_
timestamp 1698175906
transform -1 0 19824 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1143_
timestamp 1698175906
transform 1 0 14784 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1144_
timestamp 1698175906
transform 1 0 26432 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28784 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1146_
timestamp 1698175906
transform -1 0 29232 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1147_
timestamp 1698175906
transform -1 0 24640 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1148_
timestamp 1698175906
transform 1 0 27664 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1149_
timestamp 1698175906
transform 1 0 29792 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1150_
timestamp 1698175906
transform -1 0 30688 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1151_
timestamp 1698175906
transform 1 0 50960 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1152_
timestamp 1698175906
transform 1 0 16352 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27328 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1154_
timestamp 1698175906
transform 1 0 29120 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1155_
timestamp 1698175906
transform -1 0 19488 0 -1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1156_
timestamp 1698175906
transform 1 0 33936 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1157_
timestamp 1698175906
transform 1 0 25536 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1158_
timestamp 1698175906
transform 1 0 28112 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1159_
timestamp 1698175906
transform -1 0 27664 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1160_
timestamp 1698175906
transform 1 0 27328 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1161_
timestamp 1698175906
transform -1 0 29568 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1162_
timestamp 1698175906
transform -1 0 19936 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1163_
timestamp 1698175906
transform -1 0 27328 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17024 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1165_
timestamp 1698175906
transform 1 0 17808 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1166_
timestamp 1698175906
transform 1 0 18928 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1167_
timestamp 1698175906
transform -1 0 19376 0 -1 25088
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1169_
timestamp 1698175906
transform 1 0 27552 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1170_
timestamp 1698175906
transform 1 0 24864 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1171_
timestamp 1698175906
transform 1 0 26320 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1172_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28560 0 -1 12544
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1173_
timestamp 1698175906
transform -1 0 28784 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1174_
timestamp 1698175906
transform 1 0 21280 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1175_
timestamp 1698175906
transform -1 0 23856 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1176_
timestamp 1698175906
transform 1 0 22624 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1177_
timestamp 1698175906
transform 1 0 25200 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1178_
timestamp 1698175906
transform -1 0 28336 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 35056 0 -1 17248
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1180_
timestamp 1698175906
transform 1 0 27440 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1181_
timestamp 1698175906
transform 1 0 24304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_1  _1182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25200 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1183_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26544 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1184_
timestamp 1698175906
transform 1 0 28560 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1185_
timestamp 1698175906
transform -1 0 77280 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1186_
timestamp 1698175906
transform 1 0 40768 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1187_
timestamp 1698175906
transform 1 0 38528 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1188_
timestamp 1698175906
transform -1 0 24864 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1189_
timestamp 1698175906
transform -1 0 37968 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1190_
timestamp 1698175906
transform -1 0 37520 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1191_
timestamp 1698175906
transform -1 0 38528 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _1192_
timestamp 1698175906
transform -1 0 28560 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1193_
timestamp 1698175906
transform 1 0 35952 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1194_
timestamp 1698175906
transform 1 0 39648 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1195_
timestamp 1698175906
transform 1 0 23856 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1196_
timestamp 1698175906
transform -1 0 26208 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1197_
timestamp 1698175906
transform 1 0 21728 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1198_
timestamp 1698175906
transform 1 0 22624 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1199_
timestamp 1698175906
transform -1 0 28784 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1200_
timestamp 1698175906
transform -1 0 36288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1201_
timestamp 1698175906
transform -1 0 29232 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1202_
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1203_
timestamp 1698175906
transform 1 0 22512 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1204_
timestamp 1698175906
transform 1 0 27664 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1205_
timestamp 1698175906
transform 1 0 27216 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1206_
timestamp 1698175906
transform 1 0 21840 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1207_
timestamp 1698175906
transform -1 0 22848 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1208_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19600 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1209_
timestamp 1698175906
transform -1 0 21952 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1210_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 1 25088
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1211_
timestamp 1698175906
transform -1 0 3248 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1212_
timestamp 1698175906
transform -1 0 15904 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1213_
timestamp 1698175906
transform -1 0 27328 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1214_
timestamp 1698175906
transform 1 0 15568 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1215_
timestamp 1698175906
transform 1 0 17024 0 1 15680
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1216_
timestamp 1698175906
transform 1 0 11760 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1217_
timestamp 1698175906
transform 1 0 10192 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1218_
timestamp 1698175906
transform -1 0 33824 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1219_
timestamp 1698175906
transform 1 0 37296 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1220_
timestamp 1698175906
transform -1 0 31472 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1221_
timestamp 1698175906
transform -1 0 12320 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1222_
timestamp 1698175906
transform 1 0 11088 0 -1 15680
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1223_
timestamp 1698175906
transform -1 0 18592 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1224_
timestamp 1698175906
transform -1 0 18032 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1225_
timestamp 1698175906
transform -1 0 19152 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1226_
timestamp 1698175906
transform 1 0 18032 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1227_
timestamp 1698175906
transform -1 0 77280 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1228_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23520 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1229_
timestamp 1698175906
transform -1 0 21952 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1230_
timestamp 1698175906
transform -1 0 26544 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1231_
timestamp 1698175906
transform 1 0 15568 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _1232_
timestamp 1698175906
transform 1 0 10192 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1233_
timestamp 1698175906
transform 1 0 16576 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1234_
timestamp 1698175906
transform 1 0 15904 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1235_
timestamp 1698175906
transform 1 0 16128 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1236_
timestamp 1698175906
transform 1 0 28896 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1237_
timestamp 1698175906
transform -1 0 19600 0 -1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1238_
timestamp 1698175906
transform 1 0 34608 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1239_
timestamp 1698175906
transform -1 0 27216 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1240_
timestamp 1698175906
transform -1 0 20384 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1241_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18480 0 1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1242_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19488 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1243_
timestamp 1698175906
transform 1 0 27664 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1244_
timestamp 1698175906
transform 1 0 19376 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1245_
timestamp 1698175906
transform 1 0 19936 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1246_
timestamp 1698175906
transform 1 0 18144 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1247_
timestamp 1698175906
transform 1 0 27328 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1248_
timestamp 1698175906
transform -1 0 27888 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1249_
timestamp 1698175906
transform 1 0 17472 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1250_
timestamp 1698175906
transform 1 0 17584 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1251_
timestamp 1698175906
transform 1 0 18256 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1252_
timestamp 1698175906
transform -1 0 20944 0 1 31360
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1253_
timestamp 1698175906
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1254_
timestamp 1698175906
transform -1 0 35392 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1255_
timestamp 1698175906
transform 1 0 15680 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1256_
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1257_
timestamp 1698175906
transform 1 0 10752 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1258_
timestamp 1698175906
transform 1 0 9856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1259_
timestamp 1698175906
transform -1 0 12432 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1260_
timestamp 1698175906
transform 1 0 11088 0 -1 18816
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1261_
timestamp 1698175906
transform -1 0 19264 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1262_
timestamp 1698175906
transform -1 0 17136 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1263_
timestamp 1698175906
transform -1 0 19152 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1264_
timestamp 1698175906
transform 1 0 17136 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1265_
timestamp 1698175906
transform -1 0 77280 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1266_
timestamp 1698175906
transform 1 0 14000 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1267_
timestamp 1698175906
transform 1 0 16576 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _1268_
timestamp 1698175906
transform 1 0 10304 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1269_
timestamp 1698175906
transform 1 0 16464 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1270_
timestamp 1698175906
transform -1 0 16128 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1271_
timestamp 1698175906
transform -1 0 15792 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1272_
timestamp 1698175906
transform -1 0 14000 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1273_
timestamp 1698175906
transform 1 0 16464 0 1 18816
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1274_
timestamp 1698175906
transform -1 0 27328 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1275_
timestamp 1698175906
transform -1 0 16128 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1276_
timestamp 1698175906
transform 1 0 12992 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1277_
timestamp 1698175906
transform 1 0 13552 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1278_
timestamp 1698175906
transform -1 0 16352 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1279_
timestamp 1698175906
transform 1 0 13776 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1280_
timestamp 1698175906
transform -1 0 18480 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1281_
timestamp 1698175906
transform -1 0 16128 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1282_
timestamp 1698175906
transform -1 0 21616 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1283_
timestamp 1698175906
transform -1 0 20944 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1284_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20832 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1285_
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1286_
timestamp 1698175906
transform 1 0 11872 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1287_
timestamp 1698175906
transform -1 0 14784 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1288_
timestamp 1698175906
transform 1 0 12096 0 -1 10976
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1289_
timestamp 1698175906
transform -1 0 21952 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1290_
timestamp 1698175906
transform 1 0 19824 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1291_
timestamp 1698175906
transform 1 0 20720 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1292_
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1293_
timestamp 1698175906
transform -1 0 77280 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1294_
timestamp 1698175906
transform -1 0 29232 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1295_
timestamp 1698175906
transform 1 0 26992 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1296_
timestamp 1698175906
transform 1 0 24976 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _1297_
timestamp 1698175906
transform -1 0 24976 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1298_
timestamp 1698175906
transform 1 0 22400 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1299_
timestamp 1698175906
transform 1 0 23744 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1300_
timestamp 1698175906
transform 1 0 24416 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1301_
timestamp 1698175906
transform -1 0 22960 0 -1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1302_
timestamp 1698175906
transform -1 0 28336 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1303_
timestamp 1698175906
transform -1 0 27328 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1304_
timestamp 1698175906
transform 1 0 25312 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1305_
timestamp 1698175906
transform -1 0 26320 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1306_
timestamp 1698175906
transform 1 0 15120 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1307_
timestamp 1698175906
transform -1 0 16912 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1308_
timestamp 1698175906
transform -1 0 18256 0 1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1309_
timestamp 1698175906
transform 1 0 24080 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1310_
timestamp 1698175906
transform 1 0 23184 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1311_
timestamp 1698175906
transform -1 0 24864 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1312_
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1313_
timestamp 1698175906
transform 1 0 25312 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1314_
timestamp 1698175906
transform 1 0 25200 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1315_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 29008 0 -1 31360
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1316_
timestamp 1698175906
transform -1 0 23744 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1317_
timestamp 1698175906
transform 1 0 21280 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1318_
timestamp 1698175906
transform 1 0 22400 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1319_
timestamp 1698175906
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1320_
timestamp 1698175906
transform 1 0 9856 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1321_
timestamp 1698175906
transform -1 0 12656 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1322_
timestamp 1698175906
transform 1 0 11200 0 -1 20384
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1323_
timestamp 1698175906
transform -1 0 20384 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1324_
timestamp 1698175906
transform -1 0 20608 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1325_
timestamp 1698175906
transform 1 0 20608 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1326_
timestamp 1698175906
transform 1 0 22736 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1327_
timestamp 1698175906
transform -1 0 77392 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1328_
timestamp 1698175906
transform -1 0 22176 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _1329_
timestamp 1698175906
transform 1 0 10192 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1330_
timestamp 1698175906
transform 1 0 18032 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1331_
timestamp 1698175906
transform 1 0 19040 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1332_
timestamp 1698175906
transform 1 0 20384 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1333_
timestamp 1698175906
transform -1 0 22064 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1334_
timestamp 1698175906
transform -1 0 24416 0 -1 18816
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1335_
timestamp 1698175906
transform -1 0 26768 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1336_
timestamp 1698175906
transform -1 0 21280 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1337_
timestamp 1698175906
transform 1 0 20160 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1338_
timestamp 1698175906
transform 1 0 21504 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1339_
timestamp 1698175906
transform -1 0 24080 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1340_
timestamp 1698175906
transform 1 0 21728 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1341_
timestamp 1698175906
transform -1 0 24864 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1342_
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1343_
timestamp 1698175906
transform -1 0 32144 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1344_
timestamp 1698175906
transform 1 0 31920 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1345_
timestamp 1698175906
transform -1 0 32368 0 -1 14112
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1346_
timestamp 1698175906
transform 1 0 31584 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1347_
timestamp 1698175906
transform -1 0 31584 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1348_
timestamp 1698175906
transform -1 0 32368 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1349_
timestamp 1698175906
transform 1 0 30128 0 1 14112
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1350_
timestamp 1698175906
transform 1 0 33824 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1351_
timestamp 1698175906
transform 1 0 33488 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1352_
timestamp 1698175906
transform -1 0 33488 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1353_
timestamp 1698175906
transform 1 0 32368 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1354_
timestamp 1698175906
transform -1 0 77280 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1355_
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1356_
timestamp 1698175906
transform 1 0 34832 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1357_
timestamp 1698175906
transform 1 0 32032 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1358_
timestamp 1698175906
transform -1 0 33824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1359_
timestamp 1698175906
transform 1 0 33152 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1360_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 34832 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1361_
timestamp 1698175906
transform -1 0 34608 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1362_
timestamp 1698175906
transform 1 0 30912 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1363_
timestamp 1698175906
transform 1 0 30576 0 -1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1364_
timestamp 1698175906
transform -1 0 30688 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1365_
timestamp 1698175906
transform 1 0 29120 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1366_
timestamp 1698175906
transform 1 0 29680 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1367_
timestamp 1698175906
transform -1 0 23632 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1368_
timestamp 1698175906
transform -1 0 24976 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1369_
timestamp 1698175906
transform -1 0 25200 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1370_
timestamp 1698175906
transform 1 0 26096 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1371_
timestamp 1698175906
transform 1 0 29568 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1372_
timestamp 1698175906
transform -1 0 33824 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1373_
timestamp 1698175906
transform -1 0 31808 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1374_
timestamp 1698175906
transform 1 0 31920 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1375_
timestamp 1698175906
transform 1 0 34720 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1376_
timestamp 1698175906
transform -1 0 32144 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1377_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 34720 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1378_
timestamp 1698175906
transform -1 0 34384 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1379_
timestamp 1698175906
transform -1 0 32368 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1380_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 42784 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1381_
timestamp 1698175906
transform 1 0 52528 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1382_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 38192 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1383_
timestamp 1698175906
transform 1 0 51520 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1384_
timestamp 1698175906
transform 1 0 37744 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1385_
timestamp 1698175906
transform 1 0 51184 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1386_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 50176 0 -1 12544
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1387_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1388_
timestamp 1698175906
transform 1 0 39424 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1389_
timestamp 1698175906
transform 1 0 48608 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1390_
timestamp 1698175906
transform 1 0 40656 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1391_
timestamp 1698175906
transform 1 0 47488 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1392_
timestamp 1698175906
transform 1 0 39872 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1393_
timestamp 1698175906
transform 1 0 39200 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_4  _1394_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 44016 0 1 12544
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1395_
timestamp 1698175906
transform 1 0 46480 0 1 14112
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1396_
timestamp 1698175906
transform 1 0 48608 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1397_
timestamp 1698175906
transform 1 0 30912 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1398_
timestamp 1698175906
transform 1 0 33040 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1399_
timestamp 1698175906
transform -1 0 49616 0 1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _1400_
timestamp 1698175906
transform 1 0 40992 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1401_
timestamp 1698175906
transform 1 0 41104 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1402_
timestamp 1698175906
transform -1 0 44016 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1403_
timestamp 1698175906
transform -1 0 42336 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1404_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 36624 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1405_
timestamp 1698175906
transform -1 0 36960 0 -1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1406_
timestamp 1698175906
transform 1 0 31808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1407_
timestamp 1698175906
transform -1 0 34832 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1408_
timestamp 1698175906
transform -1 0 33936 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1409_
timestamp 1698175906
transform -1 0 35504 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1410_
timestamp 1698175906
transform 1 0 31024 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1411_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 30128 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1412_
timestamp 1698175906
transform 1 0 32032 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1413_
timestamp 1698175906
transform 1 0 29232 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1414_
timestamp 1698175906
transform 1 0 33264 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1415_
timestamp 1698175906
transform 1 0 32144 0 1 26656
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1416_
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1417_
timestamp 1698175906
transform 1 0 39536 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1418_
timestamp 1698175906
transform 1 0 50848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1419_
timestamp 1698175906
transform 1 0 37072 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1420_
timestamp 1698175906
transform 1 0 50960 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1421_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 60704 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1422_
timestamp 1698175906
transform 1 0 56560 0 -1 14112
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1423_
timestamp 1698175906
transform -1 0 59472 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1424_
timestamp 1698175906
transform 1 0 58352 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1425_
timestamp 1698175906
transform 1 0 46592 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1426_
timestamp 1698175906
transform 1 0 57792 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1427_
timestamp 1698175906
transform 1 0 56448 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1428_
timestamp 1698175906
transform -1 0 60032 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1429_
timestamp 1698175906
transform 1 0 55440 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1430_
timestamp 1698175906
transform 1 0 54544 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1431_
timestamp 1698175906
transform 1 0 57680 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1432_
timestamp 1698175906
transform 1 0 54992 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1433_
timestamp 1698175906
transform -1 0 57232 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1434_
timestamp 1698175906
transform 1 0 57120 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1435_
timestamp 1698175906
transform 1 0 55104 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1436_
timestamp 1698175906
transform 1 0 56448 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1437_
timestamp 1698175906
transform -1 0 59024 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1438_
timestamp 1698175906
transform -1 0 50288 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1439_
timestamp 1698175906
transform 1 0 30912 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1440_
timestamp 1698175906
transform 1 0 35168 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1441_
timestamp 1698175906
transform -1 0 35280 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1442_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1443_
timestamp 1698175906
transform 1 0 18592 0 1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1444_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 33600 0 1 29792
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1445_
timestamp 1698175906
transform -1 0 31920 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1446_
timestamp 1698175906
transform -1 0 35168 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1447_
timestamp 1698175906
transform -1 0 35056 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1448_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 30464 0 1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1449_
timestamp 1698175906
transform -1 0 32592 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1450_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 34496 0 1 32928
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1451_
timestamp 1698175906
transform -1 0 32704 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1452_
timestamp 1698175906
transform -1 0 31696 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1453_
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1454_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 31248 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1455_
timestamp 1698175906
transform 1 0 33152 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1456_
timestamp 1698175906
transform -1 0 67984 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1457_
timestamp 1698175906
transform -1 0 69552 0 -1 14112
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1458_
timestamp 1698175906
transform 1 0 65408 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1459_
timestamp 1698175906
transform 1 0 65072 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1460_
timestamp 1698175906
transform 1 0 44800 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1461_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 67200 0 1 12544
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1462_
timestamp 1698175906
transform -1 0 64064 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1463_
timestamp 1698175906
transform 1 0 63728 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1464_
timestamp 1698175906
transform 1 0 64624 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1465_
timestamp 1698175906
transform 1 0 46704 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1466_
timestamp 1698175906
transform 1 0 31248 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1467_
timestamp 1698175906
transform -1 0 30576 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1468_
timestamp 1698175906
transform -1 0 30576 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1469_
timestamp 1698175906
transform -1 0 29568 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1470_
timestamp 1698175906
transform -1 0 31584 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1471_
timestamp 1698175906
transform -1 0 30688 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1472_
timestamp 1698175906
transform 1 0 30240 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1473_
timestamp 1698175906
transform 1 0 29344 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1474_
timestamp 1698175906
transform -1 0 29680 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1475_
timestamp 1698175906
transform 1 0 28000 0 -1 32928
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1476_
timestamp 1698175906
transform -1 0 4144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1477_
timestamp 1698175906
transform 1 0 56448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1478_
timestamp 1698175906
transform 1 0 52528 0 1 15680
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1479_
timestamp 1698175906
transform 1 0 54432 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1480_
timestamp 1698175906
transform 1 0 54656 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1481_
timestamp 1698175906
transform 1 0 49840 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1482_
timestamp 1698175906
transform -1 0 59584 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1483_
timestamp 1698175906
transform 1 0 55216 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1484_
timestamp 1698175906
transform -1 0 57344 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1485_
timestamp 1698175906
transform -1 0 58576 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1486_
timestamp 1698175906
transform -1 0 58240 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1487_
timestamp 1698175906
transform -1 0 54656 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1488_
timestamp 1698175906
transform -1 0 40544 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1489_
timestamp 1698175906
transform 1 0 39760 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1490_
timestamp 1698175906
transform -1 0 39424 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1491_
timestamp 1698175906
transform -1 0 38080 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1492_
timestamp 1698175906
transform 1 0 27776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1493_
timestamp 1698175906
transform -1 0 32704 0 -1 34496
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1494_
timestamp 1698175906
transform 1 0 30240 0 1 34496
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1495_
timestamp 1698175906
transform -1 0 37408 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1496_
timestamp 1698175906
transform -1 0 36624 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1497_
timestamp 1698175906
transform 1 0 35840 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1498_
timestamp 1698175906
transform 1 0 36400 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1499_
timestamp 1698175906
transform 1 0 37744 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1500_
timestamp 1698175906
transform 1 0 48608 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1501_
timestamp 1698175906
transform 1 0 46816 0 1 12544
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1502_
timestamp 1698175906
transform -1 0 48384 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1503_
timestamp 1698175906
transform -1 0 51520 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1504_
timestamp 1698175906
transform 1 0 37632 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1505_
timestamp 1698175906
transform 1 0 40880 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1506_
timestamp 1698175906
transform 1 0 27328 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _1507_
timestamp 1698175906
transform 1 0 42112 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1508_
timestamp 1698175906
transform -1 0 43456 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1509_
timestamp 1698175906
transform -1 0 44240 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1510_
timestamp 1698175906
transform -1 0 44240 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1511_
timestamp 1698175906
transform 1 0 42112 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1512_
timestamp 1698175906
transform -1 0 40544 0 -1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1513_
timestamp 1698175906
transform 1 0 38752 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1514_
timestamp 1698175906
transform -1 0 39760 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1515_
timestamp 1698175906
transform 1 0 37408 0 1 32928
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1516_
timestamp 1698175906
transform 1 0 39760 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1517_
timestamp 1698175906
transform -1 0 42224 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1518_
timestamp 1698175906
transform 1 0 29568 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1519_
timestamp 1698175906
transform -1 0 40544 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1520_
timestamp 1698175906
transform 1 0 38192 0 1 31360
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1521_
timestamp 1698175906
transform 1 0 68208 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1522_
timestamp 1698175906
transform 1 0 68208 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1523_
timestamp 1698175906
transform -1 0 70224 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1524_
timestamp 1698175906
transform 1 0 68208 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1525_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 66640 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1526_
timestamp 1698175906
transform 1 0 66416 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1527_
timestamp 1698175906
transform 1 0 66640 0 -1 26656
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1528_
timestamp 1698175906
transform 1 0 69104 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1529_
timestamp 1698175906
transform 1 0 65520 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1530_
timestamp 1698175906
transform 1 0 68208 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1531_
timestamp 1698175906
transform -1 0 71120 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1532_
timestamp 1698175906
transform 1 0 60032 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1533_
timestamp 1698175906
transform 1 0 61488 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1534_
timestamp 1698175906
transform 1 0 62048 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1535_
timestamp 1698175906
transform 1 0 66528 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1536_
timestamp 1698175906
transform 1 0 66416 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1537_
timestamp 1698175906
transform -1 0 67984 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1538_
timestamp 1698175906
transform 1 0 67424 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1539_
timestamp 1698175906
transform 1 0 68208 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1540_
timestamp 1698175906
transform -1 0 69328 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1541_
timestamp 1698175906
transform 1 0 65296 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1542_
timestamp 1698175906
transform -1 0 65632 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1543_
timestamp 1698175906
transform 1 0 65744 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1544_
timestamp 1698175906
transform 1 0 65968 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1545_
timestamp 1698175906
transform -1 0 66640 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1546_
timestamp 1698175906
transform -1 0 67984 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1547_
timestamp 1698175906
transform -1 0 63504 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1548_
timestamp 1698175906
transform -1 0 37408 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1549_
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1550_
timestamp 1698175906
transform -1 0 41664 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1551_
timestamp 1698175906
transform -1 0 40096 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1552_
timestamp 1698175906
transform 1 0 33824 0 -1 34496
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1553_
timestamp 1698175906
transform 1 0 42336 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1554_
timestamp 1698175906
transform -1 0 43120 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1555_
timestamp 1698175906
transform 1 0 37296 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1556_
timestamp 1698175906
transform 1 0 35840 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1557_
timestamp 1698175906
transform 1 0 35728 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1558_
timestamp 1698175906
transform -1 0 37632 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1559_
timestamp 1698175906
transform -1 0 39536 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1560_
timestamp 1698175906
transform -1 0 36624 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1561_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 36064 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1562_
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1563_
timestamp 1698175906
transform 1 0 72128 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1564_
timestamp 1698175906
transform 1 0 70336 0 1 25088
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1565_
timestamp 1698175906
transform 1 0 72128 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1566_
timestamp 1698175906
transform -1 0 74032 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1567_
timestamp 1698175906
transform -1 0 43008 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1568_
timestamp 1698175906
transform -1 0 41664 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1569_
timestamp 1698175906
transform 1 0 72128 0 -1 25088
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1570_
timestamp 1698175906
transform -1 0 71792 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1571_
timestamp 1698175906
transform -1 0 72912 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1572_
timestamp 1698175906
transform -1 0 70784 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1573_
timestamp 1698175906
transform -1 0 63616 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1574_
timestamp 1698175906
transform -1 0 62832 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1575_
timestamp 1698175906
transform -1 0 42112 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1576_
timestamp 1698175906
transform -1 0 41104 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1577_
timestamp 1698175906
transform -1 0 38752 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1578_
timestamp 1698175906
transform -1 0 38416 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1579_
timestamp 1698175906
transform 1 0 37632 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1580_
timestamp 1698175906
transform 1 0 38752 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1581_
timestamp 1698175906
transform 1 0 38416 0 1 29792
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1582_
timestamp 1698175906
transform 1 0 70112 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1583_
timestamp 1698175906
transform 1 0 70112 0 1 21952
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1584_
timestamp 1698175906
transform 1 0 70112 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1585_
timestamp 1698175906
transform -1 0 73920 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1586_
timestamp 1698175906
transform 1 0 39648 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1587_
timestamp 1698175906
transform -1 0 40432 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1588_
timestamp 1698175906
transform -1 0 43456 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1589_
timestamp 1698175906
transform -1 0 71792 0 1 23520
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1590_
timestamp 1698175906
transform -1 0 73136 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1591_
timestamp 1698175906
transform -1 0 70112 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1592_
timestamp 1698175906
transform -1 0 69104 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1593_
timestamp 1698175906
transform -1 0 63504 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1594_
timestamp 1698175906
transform -1 0 62608 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1595_
timestamp 1698175906
transform -1 0 43008 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1596_
timestamp 1698175906
transform -1 0 39984 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1597_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 38416 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1598_
timestamp 1698175906
transform 1 0 37296 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1599_
timestamp 1698175906
transform -1 0 38416 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1600_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 38416 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1601_
timestamp 1698175906
transform 1 0 37744 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1602_
timestamp 1698175906
transform -1 0 43904 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1603_
timestamp 1698175906
transform -1 0 41664 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1604_
timestamp 1698175906
transform 1 0 39536 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1605_
timestamp 1698175906
transform 1 0 39536 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1606_
timestamp 1698175906
transform -1 0 40544 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1607_
timestamp 1698175906
transform 1 0 70112 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1608_
timestamp 1698175906
transform 1 0 69664 0 1 17248
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1609_
timestamp 1698175906
transform -1 0 71904 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1610_
timestamp 1698175906
transform 1 0 72128 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1611_
timestamp 1698175906
transform -1 0 39312 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1612_
timestamp 1698175906
transform -1 0 71008 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1613_
timestamp 1698175906
transform -1 0 70112 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1614_
timestamp 1698175906
transform 1 0 69440 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1615_
timestamp 1698175906
transform -1 0 67424 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1616_
timestamp 1698175906
transform -1 0 70224 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1617_
timestamp 1698175906
transform 1 0 65072 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1618_
timestamp 1698175906
transform -1 0 65520 0 1 21952
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1619_
timestamp 1698175906
transform -1 0 43120 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1620_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 40544 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1621_
timestamp 1698175906
transform 1 0 38976 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1622_
timestamp 1698175906
transform -1 0 38640 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1623_
timestamp 1698175906
transform -1 0 41664 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1624_
timestamp 1698175906
transform -1 0 39088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1625_
timestamp 1698175906
transform 1 0 40208 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1626_
timestamp 1698175906
transform 1 0 38640 0 1 23520
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1627_
timestamp 1698175906
transform -1 0 17248 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1628_
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1629_
timestamp 1698175906
transform -1 0 28112 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1630_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26880 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1631_
timestamp 1698175906
transform 1 0 29344 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1632_
timestamp 1698175906
transform -1 0 31584 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1633_
timestamp 1698175906
transform 1 0 15792 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1634_
timestamp 1698175906
transform -1 0 20272 0 1 23520
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1635_
timestamp 1698175906
transform -1 0 14000 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1636_
timestamp 1698175906
transform -1 0 44240 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1637_
timestamp 1698175906
transform -1 0 43904 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1638_
timestamp 1698175906
transform 1 0 39984 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1639_
timestamp 1698175906
transform 1 0 42336 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1640_
timestamp 1698175906
transform 1 0 43904 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1641_
timestamp 1698175906
transform 1 0 44464 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1642_
timestamp 1698175906
transform -1 0 74592 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1643_
timestamp 1698175906
transform 1 0 17360 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1644_
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1645_
timestamp 1698175906
transform -1 0 24752 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1646_
timestamp 1698175906
transform 1 0 49616 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1647_
timestamp 1698175906
transform 1 0 17360 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1648_
timestamp 1698175906
transform 1 0 43568 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1649_
timestamp 1698175906
transform -1 0 24528 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1650_
timestamp 1698175906
transform 1 0 23632 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1651_
timestamp 1698175906
transform -1 0 25872 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1652_
timestamp 1698175906
transform 1 0 23072 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1653_
timestamp 1698175906
transform 1 0 21504 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1654_
timestamp 1698175906
transform 1 0 49168 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1655_
timestamp 1698175906
transform -1 0 13776 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1656_
timestamp 1698175906
transform -1 0 27216 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1657_
timestamp 1698175906
transform 1 0 46032 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1658_
timestamp 1698175906
transform 1 0 17472 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1659_
timestamp 1698175906
transform 1 0 17248 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1660_
timestamp 1698175906
transform 1 0 45696 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1661_
timestamp 1698175906
transform 1 0 49952 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1662_
timestamp 1698175906
transform -1 0 18928 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1663_
timestamp 1698175906
transform -1 0 14224 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1664_
timestamp 1698175906
transform -1 0 7392 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1665_
timestamp 1698175906
transform -1 0 36400 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1666_
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1667_
timestamp 1698175906
transform -1 0 3808 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1668_
timestamp 1698175906
transform -1 0 16352 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1669_
timestamp 1698175906
transform 1 0 14224 0 -1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1670_
timestamp 1698175906
transform 1 0 15232 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1671_
timestamp 1698175906
transform 1 0 14672 0 1 25088
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1672_
timestamp 1698175906
transform -1 0 6048 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1673_
timestamp 1698175906
transform -1 0 6160 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1674_
timestamp 1698175906
transform -1 0 6160 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1675_
timestamp 1698175906
transform -1 0 20944 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1676_
timestamp 1698175906
transform 1 0 28560 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1677_
timestamp 1698175906
transform -1 0 27104 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1678_
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1679_
timestamp 1698175906
transform -1 0 20384 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1680_
timestamp 1698175906
transform -1 0 8064 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1681_
timestamp 1698175906
transform 1 0 4480 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1682_
timestamp 1698175906
transform -1 0 3360 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1683_
timestamp 1698175906
transform -1 0 27664 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1684_
timestamp 1698175906
transform -1 0 23744 0 -1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1685_
timestamp 1698175906
transform 1 0 21952 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1686_
timestamp 1698175906
transform 1 0 20048 0 -1 25088
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1687_
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1688_
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1689_
timestamp 1698175906
transform -1 0 8512 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1690_
timestamp 1698175906
transform 1 0 43680 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1691_
timestamp 1698175906
transform -1 0 46704 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1692_
timestamp 1698175906
transform -1 0 44464 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1693_
timestamp 1698175906
transform -1 0 31360 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1694_
timestamp 1698175906
transform 1 0 31360 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1695_
timestamp 1698175906
transform -1 0 35280 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1696_
timestamp 1698175906
transform -1 0 66080 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1697_
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1698_
timestamp 1698175906
transform 1 0 35392 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1699_
timestamp 1698175906
transform 1 0 45248 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1700_
timestamp 1698175906
transform -1 0 48832 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1701_
timestamp 1698175906
transform -1 0 45696 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1702_
timestamp 1698175906
transform -1 0 44800 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1703_
timestamp 1698175906
transform -1 0 42896 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1704_
timestamp 1698175906
transform 1 0 44688 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1705_
timestamp 1698175906
transform 1 0 42448 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1706_
timestamp 1698175906
transform 1 0 46480 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1707_
timestamp 1698175906
transform 1 0 48608 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1708_
timestamp 1698175906
transform 1 0 48608 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1709_
timestamp 1698175906
transform 1 0 47488 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1710_
timestamp 1698175906
transform 1 0 48720 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1711_
timestamp 1698175906
transform 1 0 50288 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1712_
timestamp 1698175906
transform -1 0 47712 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1713_
timestamp 1698175906
transform -1 0 48384 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1714_
timestamp 1698175906
transform 1 0 48608 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1715_
timestamp 1698175906
transform -1 0 56112 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1716_
timestamp 1698175906
transform 1 0 54096 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1717_
timestamp 1698175906
transform -1 0 53872 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1718_
timestamp 1698175906
transform -1 0 49952 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1719_
timestamp 1698175906
transform -1 0 48272 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1720_
timestamp 1698175906
transform -1 0 45696 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1721_
timestamp 1698175906
transform 1 0 44800 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1722_
timestamp 1698175906
transform -1 0 64064 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1723_
timestamp 1698175906
transform -1 0 66864 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1724_
timestamp 1698175906
transform -1 0 66752 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1725_
timestamp 1698175906
transform 1 0 51632 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1726_
timestamp 1698175906
transform 1 0 50848 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1727_
timestamp 1698175906
transform 1 0 53760 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1728_
timestamp 1698175906
transform 1 0 51520 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1729_
timestamp 1698175906
transform -1 0 55216 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1730_
timestamp 1698175906
transform -1 0 55216 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1731_
timestamp 1698175906
transform 1 0 51520 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1732_
timestamp 1698175906
transform 1 0 51632 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1733_
timestamp 1698175906
transform 1 0 52528 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1734_
timestamp 1698175906
transform 1 0 60704 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1735_
timestamp 1698175906
transform 1 0 46256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1736_
timestamp 1698175906
transform 1 0 64288 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1737_
timestamp 1698175906
transform 1 0 63504 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1738_
timestamp 1698175906
transform 1 0 50064 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1739_
timestamp 1698175906
transform 1 0 55216 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1740_
timestamp 1698175906
transform -1 0 55664 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1741_
timestamp 1698175906
transform -1 0 55888 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1742_
timestamp 1698175906
transform -1 0 51632 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1743_
timestamp 1698175906
transform 1 0 50624 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1744_
timestamp 1698175906
transform -1 0 49952 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1745_
timestamp 1698175906
transform 1 0 45136 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1746_
timestamp 1698175906
transform -1 0 45696 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1747_
timestamp 1698175906
transform -1 0 60928 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1748_
timestamp 1698175906
transform 1 0 55664 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1749_
timestamp 1698175906
transform 1 0 58800 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1750_
timestamp 1698175906
transform 1 0 61600 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1751_
timestamp 1698175906
transform -1 0 59248 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1752_
timestamp 1698175906
transform 1 0 59584 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1753_
timestamp 1698175906
transform -1 0 68880 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1754_
timestamp 1698175906
transform 1 0 66192 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1755_
timestamp 1698175906
transform 1 0 64848 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1756_
timestamp 1698175906
transform 1 0 59248 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1757_
timestamp 1698175906
transform -1 0 58576 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1758_
timestamp 1698175906
transform 1 0 57904 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1759_
timestamp 1698175906
transform -1 0 58240 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1760_
timestamp 1698175906
transform 1 0 57232 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1761_
timestamp 1698175906
transform 1 0 59360 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1762_
timestamp 1698175906
transform -1 0 72800 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1763_
timestamp 1698175906
transform 1 0 70224 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1764_
timestamp 1698175906
transform 1 0 69552 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1698175906
transform -1 0 61488 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1766_
timestamp 1698175906
transform 1 0 57568 0 -1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1767_
timestamp 1698175906
transform 1 0 59360 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1768_
timestamp 1698175906
transform 1 0 60368 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1769_
timestamp 1698175906
transform -1 0 74704 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1770_
timestamp 1698175906
transform 1 0 73360 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1771_
timestamp 1698175906
transform 1 0 73920 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1772_
timestamp 1698175906
transform -1 0 57456 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1773_
timestamp 1698175906
transform -1 0 57904 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1774_
timestamp 1698175906
transform 1 0 50960 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1775_
timestamp 1698175906
transform 1 0 50736 0 -1 20384
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1776_
timestamp 1698175906
transform 1 0 71568 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1777_
timestamp 1698175906
transform 1 0 72352 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1778_
timestamp 1698175906
transform -1 0 73696 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1779_
timestamp 1698175906
transform -1 0 42672 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1780_
timestamp 1698175906
transform 1 0 40880 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1781_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 42672 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1782_
timestamp 1698175906
transform -1 0 42336 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1783_
timestamp 1698175906
transform 1 0 11536 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1784_
timestamp 1698175906
transform -1 0 11312 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1785_
timestamp 1698175906
transform 1 0 26208 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1786_
timestamp 1698175906
transform 1 0 26432 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1787_
timestamp 1698175906
transform 1 0 7504 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1788_
timestamp 1698175906
transform -1 0 7840 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1789_
timestamp 1698175906
transform 1 0 5600 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1790_
timestamp 1698175906
transform -1 0 5152 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1791_
timestamp 1698175906
transform -1 0 42336 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1792_
timestamp 1698175906
transform 1 0 7504 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1793_
timestamp 1698175906
transform 1 0 7280 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1794_
timestamp 1698175906
transform 1 0 7504 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1795_
timestamp 1698175906
transform -1 0 8288 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1796_
timestamp 1698175906
transform 1 0 30800 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1797_
timestamp 1698175906
transform -1 0 31024 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1798_
timestamp 1698175906
transform 1 0 38864 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1799_
timestamp 1698175906
transform 1 0 39424 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1800_
timestamp 1698175906
transform -1 0 62160 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1801_
timestamp 1698175906
transform 1 0 54544 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1802_
timestamp 1698175906
transform -1 0 55328 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1803_
timestamp 1698175906
transform 1 0 61488 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1804_
timestamp 1698175906
transform -1 0 62496 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1805_
timestamp 1698175906
transform 1 0 52528 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1806_
timestamp 1698175906
transform -1 0 51520 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1807_
timestamp 1698175906
transform -1 0 52304 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1808_
timestamp 1698175906
transform -1 0 53200 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1809_
timestamp 1698175906
transform 1 0 76048 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1810_
timestamp 1698175906
transform 1 0 76048 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1811_
timestamp 1698175906
transform -1 0 76720 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1812_
timestamp 1698175906
transform 1 0 74144 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1813_
timestamp 1698175906
transform 1 0 74592 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1814_
timestamp 1698175906
transform -1 0 78288 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1815_
timestamp 1698175906
transform -1 0 78400 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1816_
timestamp 1698175906
transform 1 0 75376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1817_
timestamp 1698175906
transform -1 0 77504 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1818_
timestamp 1698175906
transform 1 0 76048 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1819_
timestamp 1698175906
transform -1 0 14448 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1820_
timestamp 1698175906
transform 1 0 42000 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1821_
timestamp 1698175906
transform 1 0 14672 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1822_
timestamp 1698175906
transform -1 0 45136 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1823_
timestamp 1698175906
transform -1 0 16464 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1824_
timestamp 1698175906
transform -1 0 46928 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1825_
timestamp 1698175906
transform 1 0 47376 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1826_
timestamp 1698175906
transform -1 0 43568 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1827_
timestamp 1698175906
transform -1 0 23968 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1828_
timestamp 1698175906
transform -1 0 24640 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1829_
timestamp 1698175906
transform 1 0 18928 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1830_
timestamp 1698175906
transform 1 0 42560 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1831_
timestamp 1698175906
transform 1 0 18368 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1832_
timestamp 1698175906
transform -1 0 13776 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1833_
timestamp 1698175906
transform -1 0 15680 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1834_
timestamp 1698175906
transform 1 0 14000 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1835_
timestamp 1698175906
transform -1 0 12880 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1836_
timestamp 1698175906
transform -1 0 25872 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1837_
timestamp 1698175906
transform -1 0 25984 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1838_
timestamp 1698175906
transform 1 0 25200 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1839_
timestamp 1698175906
transform -1 0 20944 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1840_
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1841_
timestamp 1698175906
transform -1 0 20720 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1842_
timestamp 1698175906
transform 1 0 42112 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1698175906
transform 1 0 42224 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1844_
timestamp 1698175906
transform -1 0 24864 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1845_
timestamp 1698175906
transform 1 0 17584 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1846_
timestamp 1698175906
transform -1 0 38080 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1847_
timestamp 1698175906
transform -1 0 37744 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1848_
timestamp 1698175906
transform 1 0 31696 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1849_
timestamp 1698175906
transform -1 0 37856 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1850_
timestamp 1698175906
transform -1 0 37072 0 -1 26656
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1851_
timestamp 1698175906
transform 1 0 45360 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1852_
timestamp 1698175906
transform -1 0 44688 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1853_
timestamp 1698175906
transform 1 0 42784 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1854_
timestamp 1698175906
transform -1 0 45360 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1855_
timestamp 1698175906
transform 1 0 42784 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1856_
timestamp 1698175906
transform 1 0 56560 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1857_
timestamp 1698175906
transform 1 0 44240 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1858_
timestamp 1698175906
transform 1 0 44800 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1859_
timestamp 1698175906
transform 1 0 44800 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1860_
timestamp 1698175906
transform -1 0 46592 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1861_
timestamp 1698175906
transform 1 0 44688 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1862_
timestamp 1698175906
transform 1 0 47152 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1863_
timestamp 1698175906
transform -1 0 46816 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1864_
timestamp 1698175906
transform 1 0 43456 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1865_
timestamp 1698175906
transform 1 0 44688 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1866_
timestamp 1698175906
transform 1 0 57456 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1867_
timestamp 1698175906
transform 1 0 48496 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1868_
timestamp 1698175906
transform 1 0 49168 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1869_
timestamp 1698175906
transform 1 0 48720 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1870_
timestamp 1698175906
transform -1 0 47040 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1871_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 47040 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1872_
timestamp 1698175906
transform -1 0 51184 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1873_
timestamp 1698175906
transform -1 0 51296 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1874_
timestamp 1698175906
transform -1 0 50400 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1875_
timestamp 1698175906
transform 1 0 47600 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1876_
timestamp 1698175906
transform -1 0 50288 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1877_
timestamp 1698175906
transform -1 0 49616 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1878_
timestamp 1698175906
transform 1 0 45696 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1879_
timestamp 1698175906
transform -1 0 47600 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1880_
timestamp 1698175906
transform 1 0 43456 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1881_
timestamp 1698175906
transform 1 0 43568 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1882_
timestamp 1698175906
transform 1 0 44240 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1883_
timestamp 1698175906
transform 1 0 50512 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1884_
timestamp 1698175906
transform 1 0 48048 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1885_
timestamp 1698175906
transform -1 0 49504 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1886_
timestamp 1698175906
transform 1 0 49504 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1887_
timestamp 1698175906
transform 1 0 49728 0 1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1888_
timestamp 1698175906
transform -1 0 52416 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1889_
timestamp 1698175906
transform -1 0 52192 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1890_
timestamp 1698175906
transform 1 0 50512 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1891_
timestamp 1698175906
transform 1 0 52752 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1892_
timestamp 1698175906
transform 1 0 53424 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1893_
timestamp 1698175906
transform 1 0 53648 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1894_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 51632 0 -1 28224
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1895_
timestamp 1698175906
transform 1 0 52528 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1896_
timestamp 1698175906
transform -1 0 52304 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1897_
timestamp 1698175906
transform 1 0 46144 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1898_
timestamp 1698175906
transform -1 0 55440 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1899_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 53984 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1900_
timestamp 1698175906
transform 1 0 55552 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1901_
timestamp 1698175906
transform 1 0 60816 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1902_
timestamp 1698175906
transform -1 0 61600 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1903_
timestamp 1698175906
transform 1 0 62384 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1904_
timestamp 1698175906
transform 1 0 60368 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1905_
timestamp 1698175906
transform 1 0 61152 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1906_
timestamp 1698175906
transform -1 0 59472 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1907_
timestamp 1698175906
transform -1 0 57568 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1908_
timestamp 1698175906
transform 1 0 59472 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1909_
timestamp 1698175906
transform -1 0 62832 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1910_
timestamp 1698175906
transform -1 0 62384 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1911_
timestamp 1698175906
transform 1 0 57792 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1912_
timestamp 1698175906
transform 1 0 58688 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1913_
timestamp 1698175906
transform -1 0 57792 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1914_
timestamp 1698175906
transform 1 0 59472 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1915_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 60144 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1916_
timestamp 1698175906
transform 1 0 59584 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1917_
timestamp 1698175906
transform -1 0 60144 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1918_
timestamp 1698175906
transform -1 0 59136 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1919_
timestamp 1698175906
transform 1 0 58352 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1920_
timestamp 1698175906
transform 1 0 59360 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1921_
timestamp 1698175906
transform 1 0 59136 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1922_
timestamp 1698175906
transform 1 0 58912 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1923_
timestamp 1698175906
transform 1 0 60480 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1924_
timestamp 1698175906
transform 1 0 50848 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1925_
timestamp 1698175906
transform -1 0 59360 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1926_
timestamp 1698175906
transform 1 0 57680 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1927_
timestamp 1698175906
transform -1 0 58016 0 1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1928_
timestamp 1698175906
transform 1 0 52304 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1929_
timestamp 1698175906
transform 1 0 53200 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1930_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 41328 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1931_
timestamp 1698175906
transform 1 0 42336 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1932_
timestamp 1698175906
transform -1 0 24304 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1933_
timestamp 1698175906
transform -1 0 41664 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1934_
timestamp 1698175906
transform 1 0 27440 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1935_
timestamp 1698175906
transform -1 0 17808 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1936_
timestamp 1698175906
transform 1 0 15120 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1937_
timestamp 1698175906
transform -1 0 26544 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1938_
timestamp 1698175906
transform -1 0 24640 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1939_
timestamp 1698175906
transform 1 0 23296 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1940_
timestamp 1698175906
transform -1 0 15456 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1941_
timestamp 1698175906
transform -1 0 14896 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1942_
timestamp 1698175906
transform -1 0 16576 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1943_
timestamp 1698175906
transform 1 0 14448 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1944_
timestamp 1698175906
transform -1 0 20944 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1945_
timestamp 1698175906
transform 1 0 19488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1946_
timestamp 1698175906
transform -1 0 22736 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1947_
timestamp 1698175906
transform 1 0 21504 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1948_
timestamp 1698175906
transform -1 0 31696 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1949_
timestamp 1698175906
transform 1 0 30352 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1950_
timestamp 1698175906
transform 1 0 38864 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1951_
timestamp 1698175906
transform -1 0 39648 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1952_
timestamp 1698175906
transform 1 0 65072 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1953_
timestamp 1698175906
transform 1 0 58128 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1954_
timestamp 1698175906
transform 1 0 57456 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1955_
timestamp 1698175906
transform -1 0 66304 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1956_
timestamp 1698175906
transform -1 0 66976 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1957_
timestamp 1698175906
transform 1 0 53536 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1958_
timestamp 1698175906
transform -1 0 53984 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1959_
timestamp 1698175906
transform 1 0 52528 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1960_
timestamp 1698175906
transform -1 0 52304 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1961_
timestamp 1698175906
transform 1 0 74256 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1962_
timestamp 1698175906
transform 1 0 76048 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1963_
timestamp 1698175906
transform 1 0 75152 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1964_
timestamp 1698175906
transform 1 0 74144 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1965_
timestamp 1698175906
transform 1 0 74032 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1966_
timestamp 1698175906
transform 1 0 76048 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1967_
timestamp 1698175906
transform -1 0 74928 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1968_
timestamp 1698175906
transform -1 0 78288 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1969_
timestamp 1698175906
transform -1 0 75824 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1970_
timestamp 1698175906
transform -1 0 77840 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1971_
timestamp 1698175906
transform 1 0 43680 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1972_
timestamp 1698175906
transform -1 0 47264 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1973_
timestamp 1698175906
transform 1 0 70896 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1974_
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1975_
timestamp 1698175906
transform -1 0 15904 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1976_
timestamp 1698175906
transform 1 0 22176 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1977_
timestamp 1698175906
transform -1 0 20944 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1978_
timestamp 1698175906
transform -1 0 38304 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1979_
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1980_
timestamp 1698175906
transform -1 0 3696 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1981_
timestamp 1698175906
transform 1 0 5488 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1982_
timestamp 1698175906
transform -1 0 3920 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1983_
timestamp 1698175906
transform 1 0 6384 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1984_
timestamp 1698175906
transform -1 0 6720 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1985_
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1986_
timestamp 1698175906
transform -1 0 10080 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1987_
timestamp 1698175906
transform -1 0 66416 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1988_
timestamp 1698175906
transform 1 0 34048 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1989_
timestamp 1698175906
transform -1 0 33824 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1990_
timestamp 1698175906
transform 1 0 40768 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1991_
timestamp 1698175906
transform -1 0 40544 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1992_
timestamp 1698175906
transform -1 0 59472 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1993_
timestamp 1698175906
transform 1 0 57120 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1994_
timestamp 1698175906
transform -1 0 66976 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1995_
timestamp 1698175906
transform -1 0 66864 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1996_
timestamp 1698175906
transform 1 0 47488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1997_
timestamp 1698175906
transform 1 0 63616 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1998_
timestamp 1698175906
transform 1 0 62608 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1999_
timestamp 1698175906
transform 1 0 47600 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2000_
timestamp 1698175906
transform 1 0 47712 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2001_
timestamp 1698175906
transform -1 0 68096 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2002_
timestamp 1698175906
transform -1 0 67872 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2003_
timestamp 1698175906
transform -1 0 71904 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2004_
timestamp 1698175906
transform -1 0 71792 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2005_
timestamp 1698175906
transform -1 0 75152 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2006_
timestamp 1698175906
transform 1 0 75152 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2007_
timestamp 1698175906
transform 1 0 72128 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2008_
timestamp 1698175906
transform 1 0 72128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2009_
timestamp 1698175906
transform 1 0 43456 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2010_
timestamp 1698175906
transform -1 0 46256 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2011_
timestamp 1698175906
transform 1 0 70336 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2012_
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2013_
timestamp 1698175906
transform -1 0 13328 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2014_
timestamp 1698175906
transform -1 0 28784 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2015_
timestamp 1698175906
transform -1 0 29680 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2016_
timestamp 1698175906
transform -1 0 10304 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2017_
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2018_
timestamp 1698175906
transform -1 0 3920 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2019_
timestamp 1698175906
transform 1 0 3472 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2020_
timestamp 1698175906
transform -1 0 3360 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2021_
timestamp 1698175906
transform 1 0 3584 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2022_
timestamp 1698175906
transform -1 0 3360 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2023_
timestamp 1698175906
transform 1 0 7504 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2024_
timestamp 1698175906
transform 1 0 6832 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2025_
timestamp 1698175906
transform -1 0 61936 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2026_
timestamp 1698175906
transform 1 0 33040 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2027_
timestamp 1698175906
transform -1 0 31808 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2028_
timestamp 1698175906
transform 1 0 48384 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2029_
timestamp 1698175906
transform 1 0 47712 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2030_
timestamp 1698175906
transform -1 0 58464 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2031_
timestamp 1698175906
transform -1 0 59136 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2032_
timestamp 1698175906
transform 1 0 62384 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2033_
timestamp 1698175906
transform 1 0 62496 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2034_
timestamp 1698175906
transform 1 0 47264 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2035_
timestamp 1698175906
transform 1 0 61824 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2036_
timestamp 1698175906
transform 1 0 61152 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2037_
timestamp 1698175906
transform -1 0 48384 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2038_
timestamp 1698175906
transform -1 0 49280 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2039_
timestamp 1698175906
transform 1 0 65968 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2040_
timestamp 1698175906
transform -1 0 65968 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2041_
timestamp 1698175906
transform -1 0 74032 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2042_
timestamp 1698175906
transform -1 0 71568 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2043_
timestamp 1698175906
transform 1 0 72128 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2044_
timestamp 1698175906
transform -1 0 71008 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2045_
timestamp 1698175906
transform -1 0 72688 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2046_
timestamp 1698175906
transform 1 0 69888 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2047_
timestamp 1698175906
transform 1 0 42672 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2048_
timestamp 1698175906
transform 1 0 44688 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2049_
timestamp 1698175906
transform 1 0 12992 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2050_
timestamp 1698175906
transform 1 0 11312 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2051_
timestamp 1698175906
transform 1 0 8736 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2052_
timestamp 1698175906
transform 1 0 26656 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2053_
timestamp 1698175906
transform -1 0 26656 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2054_
timestamp 1698175906
transform -1 0 9184 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2055_
timestamp 1698175906
transform 1 0 5040 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2056_
timestamp 1698175906
transform -1 0 4592 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2057_
timestamp 1698175906
transform 1 0 3584 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2058_
timestamp 1698175906
transform -1 0 3360 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2059_
timestamp 1698175906
transform -1 0 6384 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2060_
timestamp 1698175906
transform -1 0 6160 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2061_
timestamp 1698175906
transform 1 0 8848 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2062_
timestamp 1698175906
transform -1 0 7392 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2063_
timestamp 1698175906
transform 1 0 60704 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2064_
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2065_
timestamp 1698175906
transform 1 0 35168 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2066_
timestamp 1698175906
transform 1 0 48608 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2067_
timestamp 1698175906
transform 1 0 47712 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2068_
timestamp 1698175906
transform 1 0 53984 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2069_
timestamp 1698175906
transform -1 0 53872 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2070_
timestamp 1698175906
transform 1 0 61936 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2071_
timestamp 1698175906
transform -1 0 62272 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2072_
timestamp 1698175906
transform 1 0 44800 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2073_
timestamp 1698175906
transform 1 0 60928 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2074_
timestamp 1698175906
transform 1 0 60256 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2075_
timestamp 1698175906
transform 1 0 44688 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2076_
timestamp 1698175906
transform 1 0 44688 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2077_
timestamp 1698175906
transform 1 0 66080 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2078_
timestamp 1698175906
transform -1 0 66080 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2079_
timestamp 1698175906
transform 1 0 69888 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2080_
timestamp 1698175906
transform -1 0 70336 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2081_
timestamp 1698175906
transform 1 0 69776 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2082_
timestamp 1698175906
transform 1 0 69552 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2083_
timestamp 1698175906
transform 1 0 67424 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2084_
timestamp 1698175906
transform 1 0 68208 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2085_
timestamp 1698175906
transform 1 0 43344 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _2086_
timestamp 1698175906
transform -1 0 46592 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2087_
timestamp 1698175906
transform 1 0 68656 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2088_
timestamp 1698175906
transform 1 0 17696 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2089_
timestamp 1698175906
transform -1 0 16128 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2090_
timestamp 1698175906
transform 1 0 23184 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2091_
timestamp 1698175906
transform -1 0 23520 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2092_
timestamp 1698175906
transform 1 0 12208 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2093_
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2094_
timestamp 1698175906
transform -1 0 8960 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2095_
timestamp 1698175906
transform 1 0 11424 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2096_
timestamp 1698175906
transform -1 0 11872 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2097_
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2098_
timestamp 1698175906
transform 1 0 8400 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2099_
timestamp 1698175906
transform 1 0 13664 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2100_
timestamp 1698175906
transform -1 0 11872 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2101_
timestamp 1698175906
transform -1 0 37856 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2102_
timestamp 1698175906
transform 1 0 34272 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2103_
timestamp 1698175906
transform -1 0 34496 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2104_
timestamp 1698175906
transform 1 0 42672 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2105_
timestamp 1698175906
transform 1 0 43120 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2106_
timestamp 1698175906
transform 1 0 57568 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2107_
timestamp 1698175906
transform -1 0 58016 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2108_
timestamp 1698175906
transform 1 0 61712 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2109_
timestamp 1698175906
transform -1 0 62272 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2110_
timestamp 1698175906
transform 1 0 46816 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2111_
timestamp 1698175906
transform 1 0 58016 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2112_
timestamp 1698175906
transform 1 0 57792 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2113_
timestamp 1698175906
transform 1 0 47376 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2114_
timestamp 1698175906
transform -1 0 47376 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2115_
timestamp 1698175906
transform 1 0 64624 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2116_
timestamp 1698175906
transform 1 0 63392 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2117_
timestamp 1698175906
transform 1 0 66192 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2118_
timestamp 1698175906
transform 1 0 66304 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2119_
timestamp 1698175906
transform -1 0 71904 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2120_
timestamp 1698175906
transform 1 0 72128 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2121_
timestamp 1698175906
transform -1 0 70112 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2122_
timestamp 1698175906
transform 1 0 68992 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2124_
timestamp 1698175906
transform 1 0 21280 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2125_
timestamp 1698175906
transform 1 0 2016 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2126_
timestamp 1698175906
transform 1 0 2016 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2127_
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2128_
timestamp 1698175906
transform 1 0 6944 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2129_
timestamp 1698175906
transform -1 0 37520 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 43456 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2131_
timestamp 1698175906
transform 1 0 52192 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2132_
timestamp 1698175906
transform 1 0 64848 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2133_
timestamp 1698175906
transform 1 0 64176 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2134_
timestamp 1698175906
transform 1 0 44240 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2135_
timestamp 1698175906
transform 1 0 64624 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2136_
timestamp 1698175906
transform 1 0 70000 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2137_
timestamp 1698175906
transform -1 0 77840 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2138_
timestamp 1698175906
transform 1 0 72464 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2139_
timestamp 1698175906
transform 1 0 9632 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2140_
timestamp 1698175906
transform 1 0 25984 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2141_
timestamp 1698175906
transform 1 0 5936 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2142_
timestamp 1698175906
transform 1 0 2688 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2143_
timestamp 1698175906
transform -1 0 9184 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2144_
timestamp 1698175906
transform 1 0 5936 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2145_
timestamp 1698175906
transform 1 0 29456 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2146_
timestamp 1698175906
transform 1 0 38752 0 1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2147_
timestamp 1698175906
transform 1 0 53872 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2148_
timestamp 1698175906
transform 1 0 60704 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2149_
timestamp 1698175906
transform 1 0 49840 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2150_
timestamp 1698175906
transform -1 0 53536 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2151_
timestamp 1698175906
transform 1 0 75152 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2152_
timestamp 1698175906
transform 1 0 74032 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2153_
timestamp 1698175906
transform 1 0 74928 0 -1 21952
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2154_
timestamp 1698175906
transform -1 0 78064 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2155_
timestamp 1698175906
transform 1 0 13552 0 -1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2156_
timestamp 1698175906
transform 1 0 21280 0 1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2157_
timestamp 1698175906
transform 1 0 10080 0 -1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2158_
timestamp 1698175906
transform 1 0 10752 0 -1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2159_
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2160_
timestamp 1698175906
transform 1 0 19152 0 -1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2161_
timestamp 1698175906
transform -1 0 45248 0 -1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2162_
timestamp 1698175906
transform -1 0 61264 0 -1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2163_
timestamp 1698175906
transform 1 0 49056 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2164_
timestamp 1698175906
transform 1 0 44912 0 -1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2165_
timestamp 1698175906
transform 1 0 51184 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2166_
timestamp 1698175906
transform 1 0 51408 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2167_
timestamp 1698175906
transform 1 0 60592 0 -1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2168_
timestamp 1698175906
transform 1 0 60368 0 1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2169_
timestamp 1698175906
transform 1 0 60592 0 -1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2170_
timestamp 1698175906
transform 1 0 54208 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2171_
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2172_
timestamp 1698175906
transform -1 0 25200 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2173_
timestamp 1698175906
transform -1 0 15456 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2174_
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2175_
timestamp 1698175906
transform 1 0 18592 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2176_
timestamp 1698175906
transform -1 0 23296 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2177_
timestamp 1698175906
transform 1 0 29456 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2178_
timestamp 1698175906
transform 1 0 38192 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2179_
timestamp 1698175906
transform 1 0 57680 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2180_
timestamp 1698175906
transform 1 0 64736 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2181_
timestamp 1698175906
transform 1 0 52528 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2182_
timestamp 1698175906
transform 1 0 50736 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2183_
timestamp 1698175906
transform 1 0 74704 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2184_
timestamp 1698175906
transform 1 0 74704 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2185_
timestamp 1698175906
transform 1 0 73360 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2186_
timestamp 1698175906
transform -1 0 78400 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2187_
timestamp 1698175906
transform 1 0 13776 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2188_
timestamp 1698175906
transform 1 0 19712 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2189_
timestamp 1698175906
transform 1 0 1792 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2190_
timestamp 1698175906
transform 1 0 2240 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2191_
timestamp 1698175906
transform 1 0 5376 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2192_
timestamp 1698175906
transform 1 0 8288 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2193_
timestamp 1698175906
transform 1 0 31808 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2194_
timestamp 1698175906
transform 1 0 38752 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2195_
timestamp 1698175906
transform 1 0 57232 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2196_
timestamp 1698175906
transform 1 0 65072 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2197_
timestamp 1698175906
transform -1 0 64064 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2198_
timestamp 1698175906
transform 1 0 47376 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2199_
timestamp 1698175906
transform 1 0 65520 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2200_
timestamp 1698175906
transform 1 0 69888 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2201_
timestamp 1698175906
transform -1 0 78064 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2202_
timestamp 1698175906
transform 1 0 70560 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2203_
timestamp 1698175906
transform 1 0 9856 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2204_
timestamp 1698175906
transform -1 0 29792 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2205_
timestamp 1698175906
transform 1 0 2016 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2206_
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2207_
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2208_
timestamp 1698175906
transform 1 0 6496 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2209_
timestamp 1698175906
transform 1 0 29456 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2210_
timestamp 1698175906
transform 1 0 48608 0 -1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2211_
timestamp 1698175906
transform 1 0 56448 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2212_
timestamp 1698175906
transform -1 0 65072 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2213_
timestamp 1698175906
transform -1 0 64064 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2214_
timestamp 1698175906
transform 1 0 46368 0 1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2215_
timestamp 1698175906
transform 1 0 64400 0 1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2216_
timestamp 1698175906
transform 1 0 70336 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2217_
timestamp 1698175906
transform 1 0 69440 0 1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2218_
timestamp 1698175906
transform 1 0 69328 0 1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2219_
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2220_
timestamp 1698175906
transform 1 0 25424 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2221_
timestamp 1698175906
transform 1 0 1792 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2222_
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2223_
timestamp 1698175906
transform 1 0 2912 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2224_
timestamp 1698175906
transform 1 0 5600 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2225_
timestamp 1698175906
transform -1 0 38640 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2226_
timestamp 1698175906
transform 1 0 47600 0 1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2227_
timestamp 1698175906
transform 1 0 52080 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2228_
timestamp 1698175906
transform 1 0 60480 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2229_
timestamp 1698175906
transform 1 0 60368 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2230_
timestamp 1698175906
transform -1 0 46368 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2231_
timestamp 1698175906
transform 1 0 64512 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2232_
timestamp 1698175906
transform 1 0 68880 0 1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2233_
timestamp 1698175906
transform -1 0 72016 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2234_
timestamp 1698175906
transform -1 0 70336 0 -1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2235_
timestamp 1698175906
transform 1 0 14448 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2236_
timestamp 1698175906
transform 1 0 21840 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2237_
timestamp 1698175906
transform 1 0 7168 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2238_
timestamp 1698175906
transform 1 0 9856 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2239_
timestamp 1698175906
transform -1 0 10528 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2240_
timestamp 1698175906
transform 1 0 10416 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2241_
timestamp 1698175906
transform 1 0 32816 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2242_
timestamp 1698175906
transform 1 0 42896 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2243_
timestamp 1698175906
transform 1 0 56672 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2244_
timestamp 1698175906
transform 1 0 60928 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2245_
timestamp 1698175906
transform -1 0 60144 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2246_
timestamp 1698175906
transform 1 0 45136 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2247_
timestamp 1698175906
transform 1 0 63168 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2248_
timestamp 1698175906
transform 1 0 65856 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2249_
timestamp 1698175906
transform -1 0 74256 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2250_
timestamp 1698175906
transform 1 0 68320 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1045__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26096 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__A1
timestamp 1698175906
transform -1 0 28784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__A3
timestamp 1698175906
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__I
timestamp 1698175906
transform 1 0 25200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__A1
timestamp 1698175906
transform 1 0 25536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__A2
timestamp 1698175906
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__I
timestamp 1698175906
transform 1 0 43904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1058__I
timestamp 1698175906
transform 1 0 31584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A3
timestamp 1698175906
transform 1 0 26992 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__I
timestamp 1698175906
transform 1 0 27440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__B
timestamp 1698175906
transform 1 0 34272 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__I
timestamp 1698175906
transform 1 0 42336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1068__A1
timestamp 1698175906
transform 1 0 40208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__A1
timestamp 1698175906
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__I
timestamp 1698175906
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__A1
timestamp 1698175906
transform 1 0 39648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__B
timestamp 1698175906
transform -1 0 39424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__A2
timestamp 1698175906
transform -1 0 31360 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__I
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__I
timestamp 1698175906
transform 1 0 38752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__A1
timestamp 1698175906
transform -1 0 32256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__I
timestamp 1698175906
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__I
timestamp 1698175906
transform 1 0 25536 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__A3
timestamp 1698175906
transform 1 0 15008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__A2
timestamp 1698175906
transform 1 0 18032 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__I
timestamp 1698175906
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__I
timestamp 1698175906
transform -1 0 76160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1109__I
timestamp 1698175906
transform 1 0 55104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1110__I
timestamp 1698175906
transform -1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__I
timestamp 1698175906
transform 1 0 54096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__I
timestamp 1698175906
transform 1 0 25648 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__I
timestamp 1698175906
transform -1 0 52864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__I
timestamp 1698175906
transform 1 0 52640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1118__I
timestamp 1698175906
transform 1 0 53200 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__I
timestamp 1698175906
transform -1 0 27776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__B1
timestamp 1698175906
transform 1 0 16912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1123__I
timestamp 1698175906
transform 1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__I
timestamp 1698175906
transform -1 0 12432 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__I
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1131__I
timestamp 1698175906
transform 1 0 21056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__I
timestamp 1698175906
transform 1 0 19712 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__I
timestamp 1698175906
transform 1 0 24640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__A1
timestamp 1698175906
transform 1 0 25648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1144__I
timestamp 1698175906
transform 1 0 25760 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1145__A1
timestamp 1698175906
transform -1 0 25760 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1148__A1
timestamp 1698175906
transform 1 0 26544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1151__I
timestamp 1698175906
transform 1 0 50736 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__A2
timestamp 1698175906
transform -1 0 16576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__B
timestamp 1698175906
transform 1 0 19488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__I
timestamp 1698175906
transform 1 0 35392 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1161__A1
timestamp 1698175906
transform 1 0 30240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1161__A2
timestamp 1698175906
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__A2
timestamp 1698175906
transform 1 0 16800 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__A1
timestamp 1698175906
transform 1 0 19824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1167__A1
timestamp 1698175906
transform -1 0 19712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1171__A3
timestamp 1698175906
transform 1 0 26096 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__A2
timestamp 1698175906
transform 1 0 26320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1173__A3
timestamp 1698175906
transform 1 0 29008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1174__I
timestamp 1698175906
transform 1 0 22176 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__A2
timestamp 1698175906
transform 1 0 26880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__B1
timestamp 1698175906
transform 1 0 27104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1185__I
timestamp 1698175906
transform -1 0 76608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1186__I
timestamp 1698175906
transform 1 0 41664 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__I
timestamp 1698175906
transform 1 0 39200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1188__A2
timestamp 1698175906
transform -1 0 23856 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1188__B1
timestamp 1698175906
transform -1 0 26096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1189__I
timestamp 1698175906
transform 1 0 37520 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1190__I
timestamp 1698175906
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1191__I
timestamp 1698175906
transform -1 0 37968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__A2
timestamp 1698175906
transform 1 0 28560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__B1
timestamp 1698175906
transform 1 0 29680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__C1
timestamp 1698175906
transform 1 0 29232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__I
timestamp 1698175906
transform 1 0 36624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1194__I
timestamp 1698175906
transform -1 0 40096 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1195__A2
timestamp 1698175906
transform 1 0 23184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1195__B1
timestamp 1698175906
transform 1 0 23632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1197__A1
timestamp 1698175906
transform -1 0 23520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1197__A2
timestamp 1698175906
transform 1 0 23744 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__B
timestamp 1698175906
transform 1 0 29232 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1201__A1
timestamp 1698175906
transform -1 0 30016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1201__A2
timestamp 1698175906
transform -1 0 28000 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1209__A2
timestamp 1698175906
transform 1 0 22176 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__B1
timestamp 1698175906
transform -1 0 26096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1211__I
timestamp 1698175906
transform 1 0 3248 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1221__A2
timestamp 1698175906
transform 1 0 12320 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1221__A3
timestamp 1698175906
transform 1 0 13552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__A2
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__I
timestamp 1698175906
transform -1 0 76608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1230__I
timestamp 1698175906
transform -1 0 26992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1231__B1
timestamp 1698175906
transform 1 0 16800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__A1
timestamp 1698175906
transform -1 0 27440 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1245__A1
timestamp 1698175906
transform 1 0 20720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1247__A2
timestamp 1698175906
transform 1 0 27440 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1250__A1
timestamp 1698175906
transform -1 0 17920 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__A1
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__A2
timestamp 1698175906
transform -1 0 14448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1259__A2
timestamp 1698175906
transform -1 0 10976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1259__A3
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__A2
timestamp 1698175906
transform 1 0 15344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1261__A1
timestamp 1698175906
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1261__A2
timestamp 1698175906
transform 1 0 19824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1265__I
timestamp 1698175906
transform 1 0 76384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__A1
timestamp 1698175906
transform 1 0 18256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__B1
timestamp 1698175906
transform 1 0 17808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1269__A1
timestamp 1698175906
transform 1 0 16240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1274__A1
timestamp 1698175906
transform -1 0 28672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A1
timestamp 1698175906
transform 1 0 19040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__B2
timestamp 1698175906
transform 1 0 19712 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1281__A1
timestamp 1698175906
transform 1 0 16800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1283__A1
timestamp 1698175906
transform -1 0 20160 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1285__I
timestamp 1698175906
transform -1 0 12208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__I
timestamp 1698175906
transform 1 0 11200 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1287__A1
timestamp 1698175906
transform -1 0 11872 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1287__A2
timestamp 1698175906
transform 1 0 15456 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1287__A3
timestamp 1698175906
transform -1 0 15008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1288__A2
timestamp 1698175906
transform -1 0 17472 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1289__A1
timestamp 1698175906
transform -1 0 21168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1293__I
timestamp 1698175906
transform 1 0 76384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__A2
timestamp 1698175906
transform 1 0 29232 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A1
timestamp 1698175906
transform -1 0 24976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A2
timestamp 1698175906
transform -1 0 26208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__B1
timestamp 1698175906
transform 1 0 26768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__A1
timestamp 1698175906
transform 1 0 22176 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__A2
timestamp 1698175906
transform -1 0 25872 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__B1
timestamp 1698175906
transform -1 0 25424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__B2
timestamp 1698175906
transform 1 0 22624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__C1
timestamp 1698175906
transform 1 0 25424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__C2
timestamp 1698175906
transform 1 0 22736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1298__A1
timestamp 1698175906
transform 1 0 21728 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1298__A2
timestamp 1698175906
transform -1 0 23296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1298__B1
timestamp 1698175906
transform -1 0 23744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1301__B
timestamp 1698175906
transform 1 0 22960 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1302__A1
timestamp 1698175906
transform -1 0 28784 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1302__A2
timestamp 1698175906
transform 1 0 29008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1303__A1
timestamp 1698175906
transform 1 0 26768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1312__A1
timestamp 1698175906
transform 1 0 23968 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__A1
timestamp 1698175906
transform -1 0 21616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__A2
timestamp 1698175906
transform 1 0 22064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1318__A3
timestamp 1698175906
transform -1 0 23184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1321__A2
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1321__A3
timestamp 1698175906
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1322__A2
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1322__B1
timestamp 1698175906
transform 1 0 17920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1323__A1
timestamp 1698175906
transform 1 0 19600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1323__A2
timestamp 1698175906
transform 1 0 20384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1324__A2
timestamp 1698175906
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1324__A3
timestamp 1698175906
transform -1 0 20832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1327__I
timestamp 1698175906
transform 1 0 77616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1328__A1
timestamp 1698175906
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1328__B1
timestamp 1698175906
transform -1 0 22176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1330__A1
timestamp 1698175906
transform 1 0 17808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1341__A1
timestamp 1698175906
transform 1 0 25424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1341__B2
timestamp 1698175906
transform -1 0 26768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__A1
timestamp 1698175906
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1344__A2
timestamp 1698175906
transform 1 0 31696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__A2
timestamp 1698175906
transform 1 0 32032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__A3
timestamp 1698175906
transform 1 0 29456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1348__A3
timestamp 1698175906
transform -1 0 30912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__A2
timestamp 1698175906
transform -1 0 30128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__B1
timestamp 1698175906
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A2
timestamp 1698175906
transform 1 0 34496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A3
timestamp 1698175906
transform 1 0 34272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1354__I
timestamp 1698175906
transform 1 0 76384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1356__A2
timestamp 1698175906
transform 1 0 36064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1356__B1
timestamp 1698175906
transform 1 0 35616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__A2
timestamp 1698175906
transform -1 0 33264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__B1
timestamp 1698175906
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__A2
timestamp 1698175906
transform 1 0 34832 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__A2
timestamp 1698175906
transform -1 0 34608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__B1
timestamp 1698175906
transform 1 0 34160 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1361__A1
timestamp 1698175906
transform 1 0 33488 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1361__A2
timestamp 1698175906
transform 1 0 31024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__A1
timestamp 1698175906
transform 1 0 30688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__I
timestamp 1698175906
transform -1 0 34720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1377__B2
timestamp 1698175906
transform 1 0 33376 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1383__I
timestamp 1698175906
transform 1 0 53312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__I
timestamp 1698175906
transform 1 0 50960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__A2
timestamp 1698175906
transform -1 0 55888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__B1
timestamp 1698175906
transform -1 0 56896 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__B2
timestamp 1698175906
transform -1 0 50176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__C1
timestamp 1698175906
transform -1 0 56112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1388__A1
timestamp 1698175906
transform 1 0 42000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1389__I
timestamp 1698175906
transform -1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__A2
timestamp 1698175906
transform -1 0 37296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__B1
timestamp 1698175906
transform 1 0 37072 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__B2
timestamp 1698175906
transform 1 0 44912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1395__A1
timestamp 1698175906
transform 1 0 52976 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1395__A2
timestamp 1698175906
transform 1 0 52080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1395__B1
timestamp 1698175906
transform 1 0 52864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1397__A1
timestamp 1698175906
transform 1 0 30688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__B
timestamp 1698175906
transform -1 0 46928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__A2
timestamp 1698175906
transform 1 0 38976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__B1
timestamp 1698175906
transform -1 0 41216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__C1
timestamp 1698175906
transform 1 0 39424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__C2
timestamp 1698175906
transform 1 0 42560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1401__A1
timestamp 1698175906
transform 1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1401__A2
timestamp 1698175906
transform 1 0 40320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1401__B1
timestamp 1698175906
transform -1 0 42784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__A2
timestamp 1698175906
transform 1 0 44240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__B1
timestamp 1698175906
transform -1 0 43680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__I0
timestamp 1698175906
transform -1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__I1
timestamp 1698175906
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__S
timestamp 1698175906
transform 1 0 35728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1416__I
timestamp 1698175906
transform 1 0 2016 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1421__A2
timestamp 1698175906
transform -1 0 60816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1421__B1
timestamp 1698175906
transform -1 0 61152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1422__A2
timestamp 1698175906
transform 1 0 54432 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1422__B1
timestamp 1698175906
transform 1 0 55328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1422__C1
timestamp 1698175906
transform 1 0 54880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__A2
timestamp 1698175906
transform 1 0 59696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__B1
timestamp 1698175906
transform -1 0 57456 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1425__I
timestamp 1698175906
transform 1 0 46368 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1426__I
timestamp 1698175906
transform 1 0 59360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1427__I
timestamp 1698175906
transform 1 0 58016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__I
timestamp 1698175906
transform 1 0 56224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1430__I
timestamp 1698175906
transform 1 0 54320 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__B1
timestamp 1698175906
transform -1 0 57456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1432__I
timestamp 1698175906
transform 1 0 54768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1433__B
timestamp 1698175906
transform -1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1434__I
timestamp 1698175906
transform 1 0 58912 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1435__I
timestamp 1698175906
transform 1 0 55776 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__A1
timestamp 1698175906
transform 1 0 48160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__B
timestamp 1698175906
transform -1 0 50512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1440__A2
timestamp 1698175906
transform -1 0 35392 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__A1
timestamp 1698175906
transform -1 0 35504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1450__A1
timestamp 1698175906
transform 1 0 34720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__A2
timestamp 1698175906
transform -1 0 31248 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__B2
timestamp 1698175906
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A2
timestamp 1698175906
transform 1 0 68208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__B1
timestamp 1698175906
transform 1 0 63840 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A2
timestamp 1698175906
transform 1 0 63504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__B1
timestamp 1698175906
transform 1 0 64176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__C1
timestamp 1698175906
transform 1 0 62832 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1458__A2
timestamp 1698175906
transform 1 0 63840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1458__B1
timestamp 1698175906
transform -1 0 65184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1460__I
timestamp 1698175906
transform 1 0 45696 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__C1
timestamp 1698175906
transform 1 0 64512 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1465__I1
timestamp 1698175906
transform 1 0 48384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__I0
timestamp 1698175906
transform 1 0 30576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__I1
timestamp 1698175906
transform -1 0 33152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__A2
timestamp 1698175906
transform -1 0 28336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__A2
timestamp 1698175906
transform 1 0 29456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1473__B
timestamp 1698175906
transform -1 0 28112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A1
timestamp 1698175906
transform 1 0 27328 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A2
timestamp 1698175906
transform 1 0 34272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__B2
timestamp 1698175906
transform -1 0 28000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1476__I
timestamp 1698175906
transform 1 0 4368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__A2
timestamp 1698175906
transform 1 0 58464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__B1
timestamp 1698175906
transform 1 0 56000 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__B1
timestamp 1698175906
transform 1 0 52528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__C1
timestamp 1698175906
transform -1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1479__A2
timestamp 1698175906
transform -1 0 54432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1481__I
timestamp 1698175906
transform -1 0 49840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1483__B1
timestamp 1698175906
transform -1 0 56224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__B
timestamp 1698175906
transform 1 0 56672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A2
timestamp 1698175906
transform -1 0 39088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__A1
timestamp 1698175906
transform 1 0 41104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__A1
timestamp 1698175906
transform -1 0 40096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__A1
timestamp 1698175906
transform -1 0 35840 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1498__A2
timestamp 1698175906
transform -1 0 36400 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1498__B2
timestamp 1698175906
transform 1 0 35728 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__B1
timestamp 1698175906
transform -1 0 46816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__C1
timestamp 1698175906
transform 1 0 45920 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__A2
timestamp 1698175906
transform 1 0 46368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__A1
timestamp 1698175906
transform 1 0 41440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__A2
timestamp 1698175906
transform 1 0 43232 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__A2
timestamp 1698175906
transform 1 0 40768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__B1
timestamp 1698175906
transform 1 0 43904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__C1
timestamp 1698175906
transform 1 0 42784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1698175906
transform 1 0 42112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__B1
timestamp 1698175906
transform -1 0 42672 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1509__A2
timestamp 1698175906
transform -1 0 43232 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1509__B1
timestamp 1698175906
transform 1 0 44912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__I0
timestamp 1698175906
transform 1 0 41664 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__S
timestamp 1698175906
transform -1 0 41440 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__B2
timestamp 1698175906
transform 1 0 40992 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__I
timestamp 1698175906
transform -1 0 67984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__I
timestamp 1698175906
transform 1 0 68544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__I
timestamp 1698175906
transform 1 0 68656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__I
timestamp 1698175906
transform 1 0 65520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__I
timestamp 1698175906
transform -1 0 65072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1528__I
timestamp 1698175906
transform 1 0 69104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__I
timestamp 1698175906
transform -1 0 65520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__I
timestamp 1698175906
transform 1 0 60592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1539__I
timestamp 1698175906
transform -1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1542__B
timestamp 1698175906
transform 1 0 64512 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1554__A2
timestamp 1698175906
transform -1 0 43568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A2
timestamp 1698175906
transform 1 0 37072 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1558__A1
timestamp 1698175906
transform 1 0 35616 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__A2
timestamp 1698175906
transform -1 0 40880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__A2
timestamp 1698175906
transform 1 0 35840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1567__A2
timestamp 1698175906
transform 1 0 43232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__A2
timestamp 1698175906
transform 1 0 42336 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A2
timestamp 1698175906
transform -1 0 41328 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A2
timestamp 1698175906
transform -1 0 41776 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__B2
timestamp 1698175906
transform -1 0 38192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A2
timestamp 1698175906
transform 1 0 44128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1595__A2
timestamp 1698175906
transform 1 0 43232 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__B
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A2
timestamp 1698175906
transform -1 0 41888 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1604__A2
timestamp 1698175906
transform -1 0 40992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1604__B2
timestamp 1698175906
transform 1 0 38192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__A1
timestamp 1698175906
transform 1 0 75152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__C2
timestamp 1698175906
transform 1 0 69552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A1
timestamp 1698175906
transform -1 0 69664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__A1
timestamp 1698175906
transform 1 0 67648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1619__A2
timestamp 1698175906
transform 1 0 43344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__A1
timestamp 1698175906
transform 1 0 41888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__A1
timestamp 1698175906
transform 1 0 41888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__B
timestamp 1698175906
transform 1 0 40992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A1
timestamp 1698175906
transform 1 0 38304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A2
timestamp 1698175906
transform -1 0 39312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__I
timestamp 1698175906
transform 1 0 18928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__A2
timestamp 1698175906
transform -1 0 28112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A1
timestamp 1698175906
transform -1 0 26432 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__I
timestamp 1698175906
transform -1 0 30912 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__A1
timestamp 1698175906
transform 1 0 15008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1635__I
timestamp 1698175906
transform 1 0 14224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__I
timestamp 1698175906
transform 1 0 44912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__A1
timestamp 1698175906
transform 1 0 43232 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__I
timestamp 1698175906
transform -1 0 73696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__S
timestamp 1698175906
transform -1 0 19488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__I
timestamp 1698175906
transform 1 0 49392 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__I
timestamp 1698175906
transform 1 0 43792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__A1
timestamp 1698175906
transform 1 0 22400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__A2
timestamp 1698175906
transform -1 0 23520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__B1
timestamp 1698175906
transform -1 0 23072 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__B2
timestamp 1698175906
transform 1 0 24192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A1
timestamp 1698175906
transform 1 0 25088 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A2
timestamp 1698175906
transform -1 0 23632 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__I
timestamp 1698175906
transform 1 0 24976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__S
timestamp 1698175906
transform -1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__I
timestamp 1698175906
transform 1 0 50288 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__A2
timestamp 1698175906
transform 1 0 14000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A1
timestamp 1698175906
transform -1 0 25872 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__I
timestamp 1698175906
transform 1 0 45024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A1
timestamp 1698175906
transform 1 0 18256 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__A1
timestamp 1698175906
transform -1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__I
timestamp 1698175906
transform 1 0 45472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A1
timestamp 1698175906
transform 1 0 19376 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A2
timestamp 1698175906
transform 1 0 20272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__B2
timestamp 1698175906
transform 1 0 19824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__I
timestamp 1698175906
transform 1 0 35952 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__S
timestamp 1698175906
transform 1 0 7168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A3
timestamp 1698175906
transform 1 0 15344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A1
timestamp 1698175906
transform 1 0 14672 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A1
timestamp 1698175906
transform 1 0 16576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__I1
timestamp 1698175906
transform 1 0 6384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__S
timestamp 1698175906
transform 1 0 6832 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__A2
timestamp 1698175906
transform 1 0 21392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__A1
timestamp 1698175906
transform -1 0 29904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__A3
timestamp 1698175906
transform 1 0 26320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__A4
timestamp 1698175906
transform 1 0 25872 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A1
timestamp 1698175906
transform -1 0 26880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A2
timestamp 1698175906
transform -1 0 27328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A1
timestamp 1698175906
transform -1 0 27328 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A2
timestamp 1698175906
transform -1 0 26880 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__B2
timestamp 1698175906
transform -1 0 27328 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A2
timestamp 1698175906
transform -1 0 20608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__I1
timestamp 1698175906
transform 1 0 6384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__S
timestamp 1698175906
transform -1 0 7056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A1
timestamp 1698175906
transform -1 0 26432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A2
timestamp 1698175906
transform 1 0 27104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A1
timestamp 1698175906
transform -1 0 25984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A1
timestamp 1698175906
transform -1 0 22960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__I
timestamp 1698175906
transform -1 0 10304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__I1
timestamp 1698175906
transform 1 0 12096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__S
timestamp 1698175906
transform -1 0 11312 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A1
timestamp 1698175906
transform 1 0 43008 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A2
timestamp 1698175906
transform 1 0 43456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A3
timestamp 1698175906
transform 1 0 43456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A1
timestamp 1698175906
transform -1 0 46928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__A1
timestamp 1698175906
transform 1 0 30240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__B1
timestamp 1698175906
transform -1 0 32032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__B2
timestamp 1698175906
transform 1 0 32256 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A2
timestamp 1698175906
transform 1 0 31136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__I
timestamp 1698175906
transform 1 0 34384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__I
timestamp 1698175906
transform 1 0 64960 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__S
timestamp 1698175906
transform 1 0 38752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__A1
timestamp 1698175906
transform 1 0 44912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__A2
timestamp 1698175906
transform 1 0 42560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__A3
timestamp 1698175906
transform -1 0 44240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__A4
timestamp 1698175906
transform 1 0 46928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__A1
timestamp 1698175906
transform -1 0 44688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__A2
timestamp 1698175906
transform -1 0 46816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__B2
timestamp 1698175906
transform 1 0 45920 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__A1
timestamp 1698175906
transform -1 0 43680 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__A2
timestamp 1698175906
transform 1 0 42784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__I
timestamp 1698175906
transform 1 0 42896 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__I1
timestamp 1698175906
transform 1 0 47040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__S
timestamp 1698175906
transform 1 0 46592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__I
timestamp 1698175906
transform 1 0 47152 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__A1
timestamp 1698175906
transform 1 0 49392 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__A1
timestamp 1698175906
transform 1 0 47600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__A2
timestamp 1698175906
transform 1 0 48832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__I
timestamp 1698175906
transform 1 0 55216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__S
timestamp 1698175906
transform 1 0 56000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__A1
timestamp 1698175906
transform 1 0 45920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__A2
timestamp 1698175906
transform -1 0 45920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__B2
timestamp 1698175906
transform 1 0 45248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__A1
timestamp 1698175906
transform 1 0 44800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__A2
timestamp 1698175906
transform -1 0 44576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__I
timestamp 1698175906
transform -1 0 63392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__S
timestamp 1698175906
transform 1 0 67088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__A1
timestamp 1698175906
transform 1 0 51408 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__I
timestamp 1698175906
transform -1 0 50848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__A1
timestamp 1698175906
transform -1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__S
timestamp 1698175906
transform 1 0 63840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__A1
timestamp 1698175906
transform 1 0 49840 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__A1
timestamp 1698175906
transform -1 0 50960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__S
timestamp 1698175906
transform -1 0 47936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A1
timestamp 1698175906
transform 1 0 61712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A2
timestamp 1698175906
transform 1 0 62160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__A1
timestamp 1698175906
transform -1 0 58464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__I
timestamp 1698175906
transform -1 0 68208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__S
timestamp 1698175906
transform 1 0 65968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A1
timestamp 1698175906
transform 1 0 59248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A2
timestamp 1698175906
transform 1 0 60592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__A1
timestamp 1698175906
transform 1 0 58800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__I
timestamp 1698175906
transform 1 0 71904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__S
timestamp 1698175906
transform 1 0 69328 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__A1
timestamp 1698175906
transform 1 0 62608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__A2
timestamp 1698175906
transform -1 0 61040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A1
timestamp 1698175906
transform -1 0 59808 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A1
timestamp 1698175906
transform 1 0 60592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A2
timestamp 1698175906
transform 1 0 59360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__B2
timestamp 1698175906
transform -1 0 59136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__I
timestamp 1698175906
transform 1 0 73808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__S
timestamp 1698175906
transform 1 0 73136 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A1
timestamp 1698175906
transform 1 0 57344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__A1
timestamp 1698175906
transform 1 0 55440 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__A2
timestamp 1698175906
transform 1 0 49840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__B2
timestamp 1698175906
transform 1 0 50288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__I
timestamp 1698175906
transform 1 0 71344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__A2
timestamp 1698175906
transform -1 0 72352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__A1
timestamp 1698175906
transform 1 0 73920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__I
timestamp 1698175906
transform 1 0 40992 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__A1
timestamp 1698175906
transform 1 0 39200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__I
timestamp 1698175906
transform 1 0 43680 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__I1
timestamp 1698175906
transform 1 0 13552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__S
timestamp 1698175906
transform 1 0 14000 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__I1
timestamp 1698175906
transform 1 0 25984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__S
timestamp 1698175906
transform 1 0 28112 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__S
timestamp 1698175906
transform 1 0 9408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__S
timestamp 1698175906
transform 1 0 7280 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__I
timestamp 1698175906
transform -1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__I0
timestamp 1698175906
transform -1 0 7504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__S
timestamp 1698175906
transform 1 0 9632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__I1
timestamp 1698175906
transform 1 0 9632 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__S
timestamp 1698175906
transform 1 0 9184 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__I1
timestamp 1698175906
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__S
timestamp 1698175906
transform -1 0 32704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__I0
timestamp 1698175906
transform 1 0 40992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__I1
timestamp 1698175906
transform 1 0 41440 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__S
timestamp 1698175906
transform 1 0 40544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__I
timestamp 1698175906
transform 1 0 61040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__I1
timestamp 1698175906
transform 1 0 54320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__S
timestamp 1698175906
transform 1 0 56672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__I1
timestamp 1698175906
transform 1 0 61488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__S
timestamp 1698175906
transform 1 0 63392 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__S
timestamp 1698175906
transform 1 0 54432 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__S
timestamp 1698175906
transform 1 0 53424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__I
timestamp 1698175906
transform 1 0 76272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__I1
timestamp 1698175906
transform 1 0 77952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__I1
timestamp 1698175906
transform 1 0 74144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__I1
timestamp 1698175906
transform -1 0 76608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__I
timestamp 1698175906
transform 1 0 41776 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__A1
timestamp 1698175906
transform 1 0 16352 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__A2
timestamp 1698175906
transform 1 0 14448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__I
timestamp 1698175906
transform 1 0 45360 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__A2
timestamp 1698175906
transform -1 0 14224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__C
timestamp 1698175906
transform 1 0 16688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__I
timestamp 1698175906
transform 1 0 43904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__A1
timestamp 1698175906
transform -1 0 24864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__A2
timestamp 1698175906
transform 1 0 22848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__B
timestamp 1698175906
transform -1 0 24416 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__A1
timestamp 1698175906
transform 1 0 25312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__A2
timestamp 1698175906
transform -1 0 23744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A1
timestamp 1698175906
transform 1 0 20384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A2
timestamp 1698175906
transform 1 0 19936 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__I
timestamp 1698175906
transform 1 0 43904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__A1
timestamp 1698175906
transform 1 0 19488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__C
timestamp 1698175906
transform 1 0 19712 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__A1
timestamp 1698175906
transform 1 0 15904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__A1
timestamp 1698175906
transform -1 0 14000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__C
timestamp 1698175906
transform -1 0 15344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__A1
timestamp 1698175906
transform 1 0 26544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__A2
timestamp 1698175906
transform 1 0 26096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A1
timestamp 1698175906
transform 1 0 26656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__C
timestamp 1698175906
transform -1 0 26432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__A1
timestamp 1698175906
transform -1 0 20384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A1
timestamp 1698175906
transform 1 0 20944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A2
timestamp 1698175906
transform 1 0 22512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__C
timestamp 1698175906
transform 1 0 22960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A1
timestamp 1698175906
transform 1 0 42672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A2
timestamp 1698175906
transform -1 0 42112 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__A1
timestamp 1698175906
transform 1 0 42000 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__A2
timestamp 1698175906
transform 1 0 42784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__A3
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A1
timestamp 1698175906
transform 1 0 43904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A2
timestamp 1698175906
transform 1 0 45360 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__I0
timestamp 1698175906
transform 1 0 44688 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__I
timestamp 1698175906
transform 1 0 45584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__I
timestamp 1698175906
transform 1 0 56672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__A1
timestamp 1698175906
transform 1 0 44016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__A1
timestamp 1698175906
transform 1 0 43792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__A2
timestamp 1698175906
transform 1 0 44240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__A1
timestamp 1698175906
transform 1 0 44576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__A1
timestamp 1698175906
transform -1 0 45136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__A1
timestamp 1698175906
transform 1 0 42560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__A2
timestamp 1698175906
transform -1 0 43232 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__A1
timestamp 1698175906
transform 1 0 45808 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__A2
timestamp 1698175906
transform 1 0 48944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A1
timestamp 1698175906
transform 1 0 45360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__A1
timestamp 1698175906
transform -1 0 47600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__A1
timestamp 1698175906
transform -1 0 49616 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__A1
timestamp 1698175906
transform 1 0 44576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__A2
timestamp 1698175906
transform 1 0 43120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__A1
timestamp 1698175906
transform 1 0 43456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__A2
timestamp 1698175906
transform 1 0 49840 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__A2
timestamp 1698175906
transform -1 0 50512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__A1
timestamp 1698175906
transform 1 0 51408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__I
timestamp 1698175906
transform 1 0 46256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__A1
timestamp 1698175906
transform 1 0 54544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__A1
timestamp 1698175906
transform 1 0 53760 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__B
timestamp 1698175906
transform -1 0 60816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__A1
timestamp 1698175906
transform 1 0 60368 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__A2
timestamp 1698175906
transform 1 0 60368 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__A1
timestamp 1698175906
transform 1 0 56672 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__A2
timestamp 1698175906
transform 1 0 57120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__B
timestamp 1698175906
transform -1 0 58688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__A1
timestamp 1698175906
transform 1 0 58688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__A2
timestamp 1698175906
transform -1 0 58688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__A2
timestamp 1698175906
transform 1 0 50624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A2
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__I
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1934__I
timestamp 1698175906
transform -1 0 27440 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1935__A1
timestamp 1698175906
transform 1 0 18480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1935__A2
timestamp 1698175906
transform 1 0 17808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1937__I
timestamp 1698175906
transform -1 0 26992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1938__A1
timestamp 1698175906
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1938__A2
timestamp 1698175906
transform 1 0 25760 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__A2
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__A2
timestamp 1698175906
transform 1 0 17472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__A2
timestamp 1698175906
transform 1 0 21840 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__A2
timestamp 1698175906
transform 1 0 19264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A1
timestamp 1698175906
transform 1 0 22960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A2
timestamp 1698175906
transform -1 0 23632 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__A2
timestamp 1698175906
transform -1 0 24304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A1
timestamp 1698175906
transform 1 0 31920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A2
timestamp 1698175906
transform 1 0 32368 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__A2
timestamp 1698175906
transform 1 0 30128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__I1
timestamp 1698175906
transform 1 0 41664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__S
timestamp 1698175906
transform 1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__I
timestamp 1698175906
transform -1 0 65072 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__I1
timestamp 1698175906
transform 1 0 56784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__S
timestamp 1698175906
transform 1 0 61040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__I1
timestamp 1698175906
transform 1 0 63840 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__S
timestamp 1698175906
transform 1 0 67200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__S
timestamp 1698175906
transform -1 0 53536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__S
timestamp 1698175906
transform 1 0 54432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1961__I
timestamp 1698175906
transform 1 0 74144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__I1
timestamp 1698175906
transform 1 0 77952 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__I1
timestamp 1698175906
transform 1 0 73808 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__I1
timestamp 1698175906
transform 1 0 75600 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__I
timestamp 1698175906
transform 1 0 69776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__S
timestamp 1698175906
transform -1 0 19376 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__S
timestamp 1698175906
transform -1 0 24304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__I
timestamp 1698175906
transform 1 0 38192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1979__S
timestamp 1698175906
transform 1 0 6384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__I1
timestamp 1698175906
transform -1 0 5936 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__S
timestamp 1698175906
transform 1 0 7392 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__I1
timestamp 1698175906
transform 1 0 8288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__S
timestamp 1698175906
transform 1 0 8736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__I1
timestamp 1698175906
transform 1 0 11312 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__S
timestamp 1698175906
transform 1 0 11760 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__I
timestamp 1698175906
transform 1 0 65296 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__S
timestamp 1698175906
transform 1 0 35392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__S
timestamp 1698175906
transform -1 0 42896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__S
timestamp 1698175906
transform 1 0 59696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__S
timestamp 1698175906
transform 1 0 67200 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__S
timestamp 1698175906
transform 1 0 63504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1999__S
timestamp 1698175906
transform 1 0 50176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__S
timestamp 1698175906
transform 1 0 66192 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__S
timestamp 1698175906
transform 1 0 69216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__S
timestamp 1698175906
transform 1 0 73248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2007__A2
timestamp 1698175906
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__A2
timestamp 1698175906
transform 1 0 73248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__I
timestamp 1698175906
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__S
timestamp 1698175906
transform 1 0 15008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__S
timestamp 1698175906
transform -1 0 29456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__I
timestamp 1698175906
transform 1 0 10528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__S
timestamp 1698175906
transform 1 0 8064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__S
timestamp 1698175906
transform 1 0 6272 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__I1
timestamp 1698175906
transform 1 0 5712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__S
timestamp 1698175906
transform 1 0 6160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__S
timestamp 1698175906
transform 1 0 9632 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2025__I
timestamp 1698175906
transform 1 0 59920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__S
timestamp 1698175906
transform -1 0 35168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__S
timestamp 1698175906
transform -1 0 50512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__S
timestamp 1698175906
transform 1 0 59360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__S
timestamp 1698175906
transform -1 0 61824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__S
timestamp 1698175906
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__S
timestamp 1698175906
transform -1 0 49728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2039__S
timestamp 1698175906
transform 1 0 67872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__S
timestamp 1698175906
transform -1 0 72576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__S
timestamp 1698175906
transform 1 0 72240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A1
timestamp 1698175906
transform 1 0 73360 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A2
timestamp 1698175906
transform 1 0 72576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__A1
timestamp 1698175906
transform 1 0 71680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__A2
timestamp 1698175906
transform -1 0 72352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__I
timestamp 1698175906
transform -1 0 14336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__S
timestamp 1698175906
transform 1 0 14560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__S
timestamp 1698175906
transform 1 0 25760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2054__I
timestamp 1698175906
transform 1 0 9184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__S
timestamp 1698175906
transform 1 0 7616 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2057__S
timestamp 1698175906
transform 1 0 5712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__I1
timestamp 1698175906
transform 1 0 6608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__S
timestamp 1698175906
transform 1 0 7056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__S
timestamp 1698175906
transform 1 0 8624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__I
timestamp 1698175906
transform 1 0 60592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__S
timestamp 1698175906
transform -1 0 38752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2066__S
timestamp 1698175906
transform -1 0 50736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2068__S
timestamp 1698175906
transform -1 0 55104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2070__S
timestamp 1698175906
transform 1 0 63840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__S
timestamp 1698175906
transform 1 0 60032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2075__S
timestamp 1698175906
transform 1 0 46368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__S
timestamp 1698175906
transform 1 0 65856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__S
timestamp 1698175906
transform 1 0 69664 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2081__S
timestamp 1698175906
transform 1 0 71680 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2083__A1
timestamp 1698175906
transform -1 0 67200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2083__A2
timestamp 1698175906
transform -1 0 67424 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__A1
timestamp 1698175906
transform -1 0 68432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__A2
timestamp 1698175906
transform -1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__I
timestamp 1698175906
transform -1 0 68656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2088__I0
timestamp 1698175906
transform 1 0 17472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2088__S
timestamp 1698175906
transform -1 0 19600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__I0
timestamp 1698175906
transform 1 0 25312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__S
timestamp 1698175906
transform -1 0 25984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2092__I
timestamp 1698175906
transform -1 0 12208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2093__S
timestamp 1698175906
transform 1 0 11312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__S
timestamp 1698175906
transform -1 0 13776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2097__S
timestamp 1698175906
transform -1 0 11536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2099__I0
timestamp 1698175906
transform 1 0 15232 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2099__S
timestamp 1698175906
transform 1 0 13552 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2101__I
timestamp 1698175906
transform -1 0 38080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2102__I0
timestamp 1698175906
transform 1 0 34048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2102__S
timestamp 1698175906
transform 1 0 36176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2104__I0
timestamp 1698175906
transform 1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2104__S
timestamp 1698175906
transform -1 0 42672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2106__I0
timestamp 1698175906
transform 1 0 57120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2106__S
timestamp 1698175906
transform 1 0 56672 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2108__I0
timestamp 1698175906
transform 1 0 61264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2108__S
timestamp 1698175906
transform 1 0 60816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2111__S
timestamp 1698175906
transform 1 0 57792 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2113__S
timestamp 1698175906
transform 1 0 49280 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__I0
timestamp 1698175906
transform -1 0 64848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__S
timestamp 1698175906
transform 1 0 64176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__I0
timestamp 1698175906
transform 1 0 65632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__S
timestamp 1698175906
transform 1 0 65744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__I0
timestamp 1698175906
transform 1 0 70000 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__S
timestamp 1698175906
transform 1 0 68992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2121__A2
timestamp 1698175906
transform 1 0 70336 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__A1
timestamp 1698175906
transform 1 0 68096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__A2
timestamp 1698175906
transform 1 0 68544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__CLK
timestamp 1698175906
transform 1 0 53312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2155__CLK
timestamp 1698175906
transform 1 0 17696 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__CLK
timestamp 1698175906
transform 1 0 24976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2157__CLK
timestamp 1698175906
transform 1 0 13552 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2158__CLK
timestamp 1698175906
transform 1 0 14224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2159__CLK
timestamp 1698175906
transform -1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2160__CLK
timestamp 1698175906
transform -1 0 19152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2174__CLK
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2176__CLK
timestamp 1698175906
transform 1 0 23968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__CLK
timestamp 1698175906
transform -1 0 56112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__CLK
timestamp 1698175906
transform 1 0 56000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout84_I
timestamp 1698175906
transform -1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout85_I
timestamp 1698175906
transform -1 0 27776 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout95_I
timestamp 1698175906
transform -1 0 21392 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout98_I
timestamp 1698175906
transform 1 0 11760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout99_I
timestamp 1698175906
transform 1 0 9408 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout100_I
timestamp 1698175906
transform 1 0 12656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout101_I
timestamp 1698175906
transform -1 0 13328 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout108_I
timestamp 1698175906
transform 1 0 36848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout110_I
timestamp 1698175906
transform -1 0 38080 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout115_I
timestamp 1698175906
transform 1 0 57008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout117_I
timestamp 1698175906
transform 1 0 55328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout118_I
timestamp 1698175906
transform -1 0 50512 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout119_I
timestamp 1698175906
transform 1 0 55328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout123_I
timestamp 1698175906
transform -1 0 65520 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout124_I
timestamp 1698175906
transform -1 0 59808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout128_I
timestamp 1698175906
transform 1 0 69216 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout129_I
timestamp 1698175906
transform -1 0 68992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout132_I
timestamp 1698175906
transform 1 0 65072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout133_I
timestamp 1698175906
transform 1 0 66304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout136_I
timestamp 1698175906
transform -1 0 73584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout137_I
timestamp 1698175906
transform -1 0 69888 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout138_I
timestamp 1698175906
transform 1 0 72464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout140_I
timestamp 1698175906
transform -1 0 70448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698175906
transform -1 0 72240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698175906
transform -1 0 44016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698175906
transform -1 0 48048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698175906
transform -1 0 52080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698175906
transform -1 0 56112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698175906
transform -1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698175906
transform -1 0 64176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698175906
transform -1 0 7728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698175906
transform -1 0 11760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698175906
transform -1 0 15792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698175906
transform -1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698175906
transform -1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698175906
transform -1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698175906
transform -1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698175906
transform -1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698175906
transform -1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698175906
transform -1 0 38528 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698175906
transform -1 0 14000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698175906
transform -1 0 11536 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698175906
transform -1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698175906
transform -1 0 6608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698175906
transform -1 0 4480 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698175906
transform 1 0 3472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698175906
transform -1 0 35616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698175906
transform 1 0 34832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698175906
transform 1 0 31584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698175906
transform 1 0 31136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698175906
transform -1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698175906
transform -1 0 23744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698175906
transform -1 0 21392 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698175906
transform -1 0 18928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698175906
transform 1 0 16352 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698175906
transform -1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1698175906
transform 1 0 4704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1698175906
transform -1 0 4928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output37_I
timestamp 1698175906
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output38_I
timestamp 1698175906
transform -1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output39_I
timestamp 1698175906
transform -1 0 4928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output40_I
timestamp 1698175906
transform 1 0 5152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output41_I
timestamp 1698175906
transform -1 0 5824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output43_I
timestamp 1698175906
transform -1 0 4928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output45_I
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output46_I
timestamp 1698175906
transform -1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output47_I
timestamp 1698175906
transform -1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output49_I
timestamp 1698175906
transform -1 0 4928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output52_I
timestamp 1698175906
transform 1 0 76272 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output53_I
timestamp 1698175906
transform 1 0 72688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output54_I
timestamp 1698175906
transform -1 0 75488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output55_I
timestamp 1698175906
transform -1 0 75488 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output56_I
timestamp 1698175906
transform -1 0 72576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output57_I
timestamp 1698175906
transform 1 0 76272 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output64_I
timestamp 1698175906
transform -1 0 72576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output65_I
timestamp 1698175906
transform 1 0 75264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output66_I
timestamp 1698175906
transform 1 0 71680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output67_I
timestamp 1698175906
transform 1 0 68656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output68_I
timestamp 1698175906
transform 1 0 72352 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output73_I
timestamp 1698175906
transform 1 0 50400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output75_I
timestamp 1698175906
transform 1 0 76272 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output76_I
timestamp 1698175906
transform 1 0 73696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output77_I
timestamp 1698175906
transform 1 0 70448 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output78_I
timestamp 1698175906
transform -1 0 68656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output79_I
timestamp 1698175906
transform 1 0 65856 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output80_I
timestamp 1698175906
transform 1 0 63840 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout84
timestamp 1698175906
transform -1 0 27216 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout85
timestamp 1698175906
transform 1 0 28112 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout86
timestamp 1698175906
transform -1 0 10640 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout87
timestamp 1698175906
transform -1 0 2912 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout88
timestamp 1698175906
transform -1 0 11536 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout89
timestamp 1698175906
transform -1 0 2912 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout90
timestamp 1698175906
transform -1 0 8064 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout91
timestamp 1698175906
transform -1 0 11312 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout92
timestamp 1698175906
transform 1 0 15680 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout93
timestamp 1698175906
transform -1 0 20608 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout94
timestamp 1698175906
transform -1 0 20272 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout95
timestamp 1698175906
transform -1 0 20944 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout96
timestamp 1698175906
transform -1 0 2688 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout97
timestamp 1698175906
transform -1 0 11312 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout98
timestamp 1698175906
transform -1 0 11536 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout99
timestamp 1698175906
transform -1 0 9184 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout100
timestamp 1698175906
transform 1 0 14000 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout101
timestamp 1698175906
transform -1 0 14000 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout102
timestamp 1698175906
transform -1 0 21840 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout103
timestamp 1698175906
transform 1 0 26432 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout104
timestamp 1698175906
transform -1 0 26544 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout105
timestamp 1698175906
transform -1 0 32704 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout106
timestamp 1698175906
transform -1 0 38976 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout107
timestamp 1698175906
transform 1 0 35616 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout108
timestamp 1698175906
transform -1 0 36512 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout109
timestamp 1698175906
transform 1 0 36064 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout110
timestamp 1698175906
transform -1 0 37632 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout111
timestamp 1698175906
transform -1 0 43792 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout112
timestamp 1698175906
transform 1 0 46592 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout113
timestamp 1698175906
transform -1 0 44464 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout114
timestamp 1698175906
transform -1 0 53200 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout115
timestamp 1698175906
transform 1 0 55552 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout116
timestamp 1698175906
transform 1 0 55776 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout117
timestamp 1698175906
transform -1 0 56224 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout118
timestamp 1698175906
transform -1 0 51184 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout119
timestamp 1698175906
transform -1 0 55104 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout120
timestamp 1698175906
transform -1 0 57120 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout121
timestamp 1698175906
transform -1 0 61040 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout122
timestamp 1698175906
transform -1 0 65296 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout123
timestamp 1698175906
transform -1 0 66192 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout124
timestamp 1698175906
transform -1 0 60480 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout125
timestamp 1698175906
transform -1 0 71904 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout126
timestamp 1698175906
transform 1 0 76048 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout127
timestamp 1698175906
transform -1 0 70336 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout128
timestamp 1698175906
transform 1 0 68544 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout129
timestamp 1698175906
transform -1 0 69888 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout130
timestamp 1698175906
transform -1 0 60592 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout131
timestamp 1698175906
transform 1 0 64624 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout132
timestamp 1698175906
transform -1 0 65072 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout133
timestamp 1698175906
transform -1 0 65408 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout134
timestamp 1698175906
transform 1 0 69664 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout135
timestamp 1698175906
transform 1 0 74032 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout136
timestamp 1698175906
transform 1 0 73584 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout137
timestamp 1698175906
transform 1 0 68992 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout138
timestamp 1698175906
transform 1 0 72688 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout139
timestamp 1698175906
transform 1 0 70784 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout140
timestamp 1698175906
transform -1 0 70224 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout141
timestamp 1698175906
transform -1 0 70896 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_40 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_48 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6720 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_52
timestamp 1698175906
transform 1 0 7168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_54 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7392 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_63
timestamp 1698175906
transform 1 0 8400 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698175906
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_70 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_86
timestamp 1698175906
transform 1 0 10976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_90
timestamp 1698175906
transform 1 0 11424 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_99
timestamp 1698175906
transform 1 0 12432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698175906
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_120
timestamp 1698175906
transform 1 0 14784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_124
timestamp 1698175906
transform 1 0 15232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_126
timestamp 1698175906
transform 1 0 15456 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698175906
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_138
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_154
timestamp 1698175906
transform 1 0 18592 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_162
timestamp 1698175906
transform 1 0 19488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_166
timestamp 1698175906
transform 1 0 19936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_178
timestamp 1698175906
transform 1 0 21280 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_194
timestamp 1698175906
transform 1 0 23072 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_212
timestamp 1698175906
transform 1 0 25088 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_228
timestamp 1698175906
transform 1 0 26880 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_246
timestamp 1698175906
transform 1 0 28896 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_262
timestamp 1698175906
transform 1 0 30688 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_280
timestamp 1698175906
transform 1 0 32704 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_296
timestamp 1698175906
transform 1 0 34496 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_315
timestamp 1698175906
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_319
timestamp 1698175906
transform 1 0 37072 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_335
timestamp 1698175906
transform 1 0 38864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_337
timestamp 1698175906
transform 1 0 39088 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_344
timestamp 1698175906
transform 1 0 39872 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_351
timestamp 1698175906
transform 1 0 40656 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_367
timestamp 1698175906
transform 1 0 42448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_371
timestamp 1698175906
transform 1 0 42896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_373
timestamp 1698175906
transform 1 0 43120 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698175906
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_378
timestamp 1698175906
transform 1 0 43680 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_387
timestamp 1698175906
transform 1 0 44688 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_403
timestamp 1698175906
transform 1 0 46480 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_407
timestamp 1698175906
transform 1 0 46928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_410
timestamp 1698175906
transform 1 0 47264 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_414
timestamp 1698175906
transform 1 0 47712 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_423
timestamp 1698175906
transform 1 0 48720 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_439
timestamp 1698175906
transform 1 0 50512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_441
timestamp 1698175906
transform 1 0 50736 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_444
timestamp 1698175906
transform 1 0 51072 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_448
timestamp 1698175906
transform 1 0 51520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_450
timestamp 1698175906
transform 1 0 51744 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_459
timestamp 1698175906
transform 1 0 52752 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_475
timestamp 1698175906
transform 1 0 54544 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_478
timestamp 1698175906
transform 1 0 54880 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_486
timestamp 1698175906
transform 1 0 55776 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_495
timestamp 1698175906
transform 1 0 56784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_499
timestamp 1698175906
transform 1 0 57232 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_507
timestamp 1698175906
transform 1 0 58128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_509
timestamp 1698175906
transform 1 0 58352 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_512
timestamp 1698175906
transform 1 0 58688 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_520
timestamp 1698175906
transform 1 0 59584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_522
timestamp 1698175906
transform 1 0 59808 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_531
timestamp 1698175906
transform 1 0 60816 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_539
timestamp 1698175906
transform 1 0 61712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_543
timestamp 1698175906
transform 1 0 62160 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_546
timestamp 1698175906
transform 1 0 62496 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_554
timestamp 1698175906
transform 1 0 63392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_558
timestamp 1698175906
transform 1 0 63840 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_569
timestamp 1698175906
transform 1 0 65072 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_577
timestamp 1698175906
transform 1 0 65968 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_580
timestamp 1698175906
transform 1 0 66304 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_584
timestamp 1698175906
transform 1 0 66752 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_588
timestamp 1698175906
transform 1 0 67200 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_592
timestamp 1698175906
transform 1 0 67648 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_595
timestamp 1698175906
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_599
timestamp 1698175906
transform 1 0 68432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_603
timestamp 1698175906
transform 1 0 68880 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_611
timestamp 1698175906
transform 1 0 69776 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_614
timestamp 1698175906
transform 1 0 70112 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_630
timestamp 1698175906
transform 1 0 71904 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_639
timestamp 1698175906
transform 1 0 72912 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_643
timestamp 1698175906
transform 1 0 73360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_645
timestamp 1698175906
transform 1 0 73584 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_648
timestamp 1698175906
transform 1 0 73920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_652
timestamp 1698175906
transform 1 0 74368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_682
timestamp 1698175906
transform 1 0 77728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_686
timestamp 1698175906
transform 1 0 78176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_28
timestamp 1698175906
transform 1 0 4480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_32
timestamp 1698175906
transform 1 0 4928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5376 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_68
timestamp 1698175906
transform 1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_107
timestamp 1698175906
transform 1 0 13328 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_158
timestamp 1698175906
transform 1 0 19040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_162
timestamp 1698175906
transform 1 0 19488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_193
timestamp 1698175906
transform 1 0 22960 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_216
timestamp 1698175906
transform 1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_241
timestamp 1698175906
transform 1 0 28336 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_249
timestamp 1698175906
transform 1 0 29232 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_298
timestamp 1698175906
transform 1 0 34720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_302
timestamp 1698175906
transform 1 0 35168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_333
timestamp 1698175906
transform 1 0 38640 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_341
timestamp 1698175906
transform 1 0 39536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_343
timestamp 1698175906
transform 1 0 39760 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_367
timestamp 1698175906
transform 1 0 42448 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_371
timestamp 1698175906
transform 1 0 42896 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_375
timestamp 1698175906
transform 1 0 43344 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_407
timestamp 1698175906
transform 1 0 46928 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_411
timestamp 1698175906
transform 1 0 47376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_413
timestamp 1698175906
transform 1 0 47600 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_437
timestamp 1698175906
transform 1 0 50288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_441
timestamp 1698175906
transform 1 0 50736 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_449
timestamp 1698175906
transform 1 0 51632 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_482
timestamp 1698175906
transform 1 0 55328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_523
timestamp 1698175906
transform 1 0 59920 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_527
timestamp 1698175906
transform 1 0 60368 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_557
timestamp 1698175906
transform 1 0 63728 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_559
timestamp 1698175906
transform 1 0 63952 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_562
timestamp 1698175906
transform 1 0 64288 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_566
timestamp 1698175906
transform 1 0 64736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_568
timestamp 1698175906
transform 1 0 64960 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_624
timestamp 1698175906
transform 1 0 71232 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_628
timestamp 1698175906
transform 1 0 71680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_632
timestamp 1698175906
transform 1 0 72128 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_648
timestamp 1698175906
transform 1 0 73920 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_656
timestamp 1698175906
transform 1 0 74816 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_660
timestamp 1698175906
transform 1 0 75264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_59
timestamp 1698175906
transform 1 0 7952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_63
timestamp 1698175906
transform 1 0 8400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_65
timestamp 1698175906
transform 1 0 8624 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_72
timestamp 1698175906
transform 1 0 9408 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_122
timestamp 1698175906
transform 1 0 15008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_130
timestamp 1698175906
transform 1 0 15904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_161
timestamp 1698175906
transform 1 0 19376 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_207
timestamp 1698175906
transform 1 0 24528 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698175906
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_253
timestamp 1698175906
transform 1 0 29680 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_261
timestamp 1698175906
transform 1 0 30576 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_265
timestamp 1698175906
transform 1 0 31024 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_301
timestamp 1698175906
transform 1 0 35056 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698175906
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_332
timestamp 1698175906
transform 1 0 38528 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_363
timestamp 1698175906
transform 1 0 42000 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_402
timestamp 1698175906
transform 1 0 46368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_406
timestamp 1698175906
transform 1 0 46816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_410
timestamp 1698175906
transform 1 0 47264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_412
timestamp 1698175906
transform 1 0 47488 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_444
timestamp 1698175906
transform 1 0 51072 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_452
timestamp 1698175906
transform 1 0 51968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_454
timestamp 1698175906
transform 1 0 52192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_469
timestamp 1698175906
transform 1 0 53872 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_485
timestamp 1698175906
transform 1 0 55664 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_492
timestamp 1698175906
transform 1 0 56448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_494
timestamp 1698175906
transform 1 0 56672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_516
timestamp 1698175906
transform 1 0 59136 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_520
timestamp 1698175906
transform 1 0 59584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_522
timestamp 1698175906
transform 1 0 59808 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_556
timestamp 1698175906
transform 1 0 63616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_560
timestamp 1698175906
transform 1 0 64064 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_564
timestamp 1698175906
transform 1 0 64512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_586
timestamp 1698175906
transform 1 0 66976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_605
timestamp 1698175906
transform 1 0 69104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_638
timestamp 1698175906
transform 1 0 72800 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_654
timestamp 1698175906
transform 1 0 74592 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_662
timestamp 1698175906
transform 1 0 75488 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_667
timestamp 1698175906
transform 1 0 76048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_677
timestamp 1698175906
transform 1 0 77168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_685
timestamp 1698175906
transform 1 0 78064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_687
timestamp 1698175906
transform 1 0 78288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_34
timestamp 1698175906
transform 1 0 5152 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_38
timestamp 1698175906
transform 1 0 5600 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_40
timestamp 1698175906
transform 1 0 5824 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_76
timestamp 1698175906
transform 1 0 9856 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_112
timestamp 1698175906
transform 1 0 13888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_116
timestamp 1698175906
transform 1 0 14336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_120
timestamp 1698175906
transform 1 0 14784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_124
timestamp 1698175906
transform 1 0 15232 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_157
timestamp 1698175906
transform 1 0 18928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_161
timestamp 1698175906
transform 1 0 19376 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_175
timestamp 1698175906
transform 1 0 20944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_179
timestamp 1698175906
transform 1 0 21392 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_201
timestamp 1698175906
transform 1 0 23856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_205
timestamp 1698175906
transform 1 0 24304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698175906
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_216
timestamp 1698175906
transform 1 0 25536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_218
timestamp 1698175906
transform 1 0 25760 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_254
timestamp 1698175906
transform 1 0 29792 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_270
timestamp 1698175906
transform 1 0 31584 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_290
timestamp 1698175906
transform 1 0 33824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_307
timestamp 1698175906
transform 1 0 35728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_309
timestamp 1698175906
transform 1 0 35952 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_324
timestamp 1698175906
transform 1 0 37632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_328
timestamp 1698175906
transform 1 0 38080 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_334
timestamp 1698175906
transform 1 0 38752 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_352
timestamp 1698175906
transform 1 0 40768 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_360
timestamp 1698175906
transform 1 0 41664 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_364
timestamp 1698175906
transform 1 0 42112 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_400
timestamp 1698175906
transform 1 0 46144 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_408
timestamp 1698175906
transform 1 0 47040 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_412
timestamp 1698175906
transform 1 0 47488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_453
timestamp 1698175906
transform 1 0 52080 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_469
timestamp 1698175906
transform 1 0 53872 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_477
timestamp 1698175906
transform 1 0 54768 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_480
timestamp 1698175906
transform 1 0 55104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_498
timestamp 1698175906
transform 1 0 57120 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_528
timestamp 1698175906
transform 1 0 60480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_544
timestamp 1698175906
transform 1 0 62272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_562
timestamp 1698175906
transform 1 0 64288 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_570
timestamp 1698175906
transform 1 0 65184 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_637
timestamp 1698175906
transform 1 0 72688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_641
timestamp 1698175906
transform 1 0 73136 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_645
timestamp 1698175906
transform 1 0 73584 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_661
timestamp 1698175906
transform 1 0 75376 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_28
timestamp 1698175906
transform 1 0 4480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1698175906
transform 1 0 4928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_69
timestamp 1698175906
transform 1 0 9072 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_91
timestamp 1698175906
transform 1 0 11536 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_99
timestamp 1698175906
transform 1 0 12432 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698175906
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_113
timestamp 1698175906
transform 1 0 14000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_117
timestamp 1698175906
transform 1 0 14448 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_149
timestamp 1698175906
transform 1 0 18032 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_165
timestamp 1698175906
transform 1 0 19824 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698175906
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698175906
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_183
timestamp 1698175906
transform 1 0 21840 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_199
timestamp 1698175906
transform 1 0 23632 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_207
timestamp 1698175906
transform 1 0 24528 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_219
timestamp 1698175906
transform 1 0 25872 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_223
timestamp 1698175906
transform 1 0 26320 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_251
timestamp 1698175906
transform 1 0 29456 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_267
timestamp 1698175906
transform 1 0 31248 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_275
timestamp 1698175906
transform 1 0 32144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_277
timestamp 1698175906
transform 1 0 32368 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_280
timestamp 1698175906
transform 1 0 32704 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_296
timestamp 1698175906
transform 1 0 34496 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_312
timestamp 1698175906
transform 1 0 36288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_314
timestamp 1698175906
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_333
timestamp 1698175906
transform 1 0 38640 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_365
timestamp 1698175906
transform 1 0 42224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_369
timestamp 1698175906
transform 1 0 42672 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_379
timestamp 1698175906
transform 1 0 43792 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_383
timestamp 1698175906
transform 1 0 44240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_387
timestamp 1698175906
transform 1 0 44688 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_419
timestamp 1698175906
transform 1 0 48272 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_435
timestamp 1698175906
transform 1 0 50064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_439
timestamp 1698175906
transform 1 0 50512 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_457
timestamp 1698175906
transform 1 0 52528 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_461
timestamp 1698175906
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_469
timestamp 1698175906
transform 1 0 53872 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_486
timestamp 1698175906
transform 1 0 55776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_490
timestamp 1698175906
transform 1 0 56224 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_519
timestamp 1698175906
transform 1 0 59472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_523
timestamp 1698175906
transform 1 0 59920 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_527
timestamp 1698175906
transform 1 0 60368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_531
timestamp 1698175906
transform 1 0 60816 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_535
timestamp 1698175906
transform 1 0 61264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_537
timestamp 1698175906
transform 1 0 61488 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_569
timestamp 1698175906
transform 1 0 65072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_581
timestamp 1698175906
transform 1 0 66416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_585
timestamp 1698175906
transform 1 0 66864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_587
timestamp 1698175906
transform 1 0 67088 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_590
timestamp 1698175906
transform 1 0 67424 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_594
timestamp 1698175906
transform 1 0 67872 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_597
timestamp 1698175906
transform 1 0 68208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_599
timestamp 1698175906
transform 1 0 68432 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_626
timestamp 1698175906
transform 1 0 71456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_630
timestamp 1698175906
transform 1 0 71904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_634
timestamp 1698175906
transform 1 0 72352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_638
timestamp 1698175906
transform 1 0 72800 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_654
timestamp 1698175906
transform 1 0 74592 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_662
timestamp 1698175906
transform 1 0 75488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_664
timestamp 1698175906
transform 1 0 75712 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_667
timestamp 1698175906
transform 1 0 76048 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_683
timestamp 1698175906
transform 1 0 77840 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_687
timestamp 1698175906
transform 1 0 78288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_6
timestamp 1698175906
transform 1 0 2016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_43
timestamp 1698175906
transform 1 0 6160 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_51
timestamp 1698175906
transform 1 0 7056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_76
timestamp 1698175906
transform 1 0 9856 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_80
timestamp 1698175906
transform 1 0 10304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_82
timestamp 1698175906
transform 1 0 10528 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_89
timestamp 1698175906
transform 1 0 11312 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_121
timestamp 1698175906
transform 1 0 14896 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_125
timestamp 1698175906
transform 1 0 15344 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_132
timestamp 1698175906
transform 1 0 16128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_146
timestamp 1698175906
transform 1 0 17696 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_154
timestamp 1698175906
transform 1 0 18592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_158
timestamp 1698175906
transform 1 0 19040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_160
timestamp 1698175906
transform 1 0 19264 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_163
timestamp 1698175906
transform 1 0 19600 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_167
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_169
timestamp 1698175906
transform 1 0 20272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_172
timestamp 1698175906
transform 1 0 20608 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_188
timestamp 1698175906
transform 1 0 22400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_192
timestamp 1698175906
transform 1 0 22848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_194
timestamp 1698175906
transform 1 0 23072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_216
timestamp 1698175906
transform 1 0 25536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_220
timestamp 1698175906
transform 1 0 25984 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_252
timestamp 1698175906
transform 1 0 29568 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_260
timestamp 1698175906
transform 1 0 30464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_262
timestamp 1698175906
transform 1 0 30688 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_278
timestamp 1698175906
transform 1 0 32480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_286
timestamp 1698175906
transform 1 0 33376 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_323
timestamp 1698175906
transform 1 0 37520 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_331
timestamp 1698175906
transform 1 0 38416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_352
timestamp 1698175906
transform 1 0 40768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_356
timestamp 1698175906
transform 1 0 41216 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_360
timestamp 1698175906
transform 1 0 41664 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_364
timestamp 1698175906
transform 1 0 42112 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_366
timestamp 1698175906
transform 1 0 42336 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_384
timestamp 1698175906
transform 1 0 44352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_388
timestamp 1698175906
transform 1 0 44800 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_422
timestamp 1698175906
transform 1 0 48608 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_489
timestamp 1698175906
transform 1 0 56112 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_492
timestamp 1698175906
transform 1 0 56448 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_524
timestamp 1698175906
transform 1 0 60032 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_540
timestamp 1698175906
transform 1 0 61824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_544
timestamp 1698175906
transform 1 0 62272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_552
timestamp 1698175906
transform 1 0 63168 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_562
timestamp 1698175906
transform 1 0 64288 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_594
timestamp 1698175906
transform 1 0 67872 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_604
timestamp 1698175906
transform 1 0 68992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_608
timestamp 1698175906
transform 1 0 69440 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_629
timestamp 1698175906
transform 1 0 71792 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_640
timestamp 1698175906
transform 1 0 73024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_644
timestamp 1698175906
transform 1 0 73472 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_660
timestamp 1698175906
transform 1 0 75264 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_668
timestamp 1698175906
transform 1 0 76160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_678
timestamp 1698175906
transform 1 0 77280 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_686
timestamp 1698175906
transform 1 0 78176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_31
timestamp 1698175906
transform 1 0 4816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_43
timestamp 1698175906
transform 1 0 6160 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_59
timestamp 1698175906
transform 1 0 7952 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_67
timestamp 1698175906
transform 1 0 8848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_69
timestamp 1698175906
transform 1 0 9072 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_72
timestamp 1698175906
transform 1 0 9408 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698175906
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_111
timestamp 1698175906
transform 1 0 13776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_115
timestamp 1698175906
transform 1 0 14224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_181
timestamp 1698175906
transform 1 0 21616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_212
timestamp 1698175906
transform 1 0 25088 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_237
timestamp 1698175906
transform 1 0 27888 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_280
timestamp 1698175906
transform 1 0 32704 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_288
timestamp 1698175906
transform 1 0 33600 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_292
timestamp 1698175906
transform 1 0 34048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_294
timestamp 1698175906
transform 1 0 34272 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_303
timestamp 1698175906
transform 1 0 35280 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_310
timestamp 1698175906
transform 1 0 36064 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698175906
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_332
timestamp 1698175906
transform 1 0 38528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_336
timestamp 1698175906
transform 1 0 38976 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_346
timestamp 1698175906
transform 1 0 40096 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_352
timestamp 1698175906
transform 1 0 40768 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_384
timestamp 1698175906
transform 1 0 44352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_393
timestamp 1698175906
transform 1 0 45360 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_401
timestamp 1698175906
transform 1 0 46256 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_433
timestamp 1698175906
transform 1 0 49840 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_449
timestamp 1698175906
transform 1 0 51632 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_453
timestamp 1698175906
transform 1 0 52080 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_457
timestamp 1698175906
transform 1 0 52528 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_473
timestamp 1698175906
transform 1 0 54320 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_483
timestamp 1698175906
transform 1 0 55440 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_491
timestamp 1698175906
transform 1 0 56336 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_493
timestamp 1698175906
transform 1 0 56560 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_496
timestamp 1698175906
transform 1 0 56896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_500
timestamp 1698175906
transform 1 0 57344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_517
timestamp 1698175906
transform 1 0 59248 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_527
timestamp 1698175906
transform 1 0 60368 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_543
timestamp 1698175906
transform 1 0 62160 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_551
timestamp 1698175906
transform 1 0 63056 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_554
timestamp 1698175906
transform 1 0 63392 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_585
timestamp 1698175906
transform 1 0 66864 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_589
timestamp 1698175906
transform 1 0 67312 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_593
timestamp 1698175906
transform 1 0 67760 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_597
timestamp 1698175906
transform 1 0 68208 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_605
timestamp 1698175906
transform 1 0 69104 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_609
timestamp 1698175906
transform 1 0 69552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_613
timestamp 1698175906
transform 1 0 70000 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_617
timestamp 1698175906
transform 1 0 70448 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_647
timestamp 1698175906
transform 1 0 73808 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_663
timestamp 1698175906
transform 1 0 75600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_667
timestamp 1698175906
transform 1 0 76048 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_683
timestamp 1698175906
transform 1 0 77840 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_687
timestamp 1698175906
transform 1 0 78288 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_28
timestamp 1698175906
transform 1 0 4480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_45
timestamp 1698175906
transform 1 0 6384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_49
timestamp 1698175906
transform 1 0 6832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_53
timestamp 1698175906
transform 1 0 7280 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_60
timestamp 1698175906
transform 1 0 8064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_87
timestamp 1698175906
transform 1 0 11088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_111
timestamp 1698175906
transform 1 0 13776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_115
timestamp 1698175906
transform 1 0 14224 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_119
timestamp 1698175906
transform 1 0 14672 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_122
timestamp 1698175906
transform 1 0 15008 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_138
timestamp 1698175906
transform 1 0 16800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_150
timestamp 1698175906
transform 1 0 18144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_183
timestamp 1698175906
transform 1 0 21840 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_191
timestamp 1698175906
transform 1 0 22736 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_198
timestamp 1698175906
transform 1 0 23520 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_249
timestamp 1698175906
transform 1 0 29232 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_257
timestamp 1698175906
transform 1 0 30128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_265
timestamp 1698175906
transform 1 0 31024 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_273
timestamp 1698175906
transform 1 0 31920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_277
timestamp 1698175906
transform 1 0 32368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698175906
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_290
timestamp 1698175906
transform 1 0 33824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_309
timestamp 1698175906
transform 1 0 35952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_313
timestamp 1698175906
transform 1 0 36400 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_321
timestamp 1698175906
transform 1 0 37296 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_325
timestamp 1698175906
transform 1 0 37744 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_328
timestamp 1698175906
transform 1 0 38080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_342
timestamp 1698175906
transform 1 0 39648 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_352
timestamp 1698175906
transform 1 0 40768 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_368
timestamp 1698175906
transform 1 0 42560 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_372
timestamp 1698175906
transform 1 0 43008 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_402
timestamp 1698175906
transform 1 0 46368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_404
timestamp 1698175906
transform 1 0 46592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_428
timestamp 1698175906
transform 1 0 49280 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_432
timestamp 1698175906
transform 1 0 49728 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_436
timestamp 1698175906
transform 1 0 50176 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_466
timestamp 1698175906
transform 1 0 53536 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_482
timestamp 1698175906
transform 1 0 55328 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_486
timestamp 1698175906
transform 1 0 55776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_492
timestamp 1698175906
transform 1 0 56448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_523
timestamp 1698175906
transform 1 0 59920 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_533
timestamp 1698175906
transform 1 0 61040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_537
timestamp 1698175906
transform 1 0 61488 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_562
timestamp 1698175906
transform 1 0 64288 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_566
timestamp 1698175906
transform 1 0 64736 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_596
timestamp 1698175906
transform 1 0 68096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_598
timestamp 1698175906
transform 1 0 68320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_614
timestamp 1698175906
transform 1 0 70112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_618
timestamp 1698175906
transform 1 0 70560 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_622
timestamp 1698175906
transform 1 0 71008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_624
timestamp 1698175906
transform 1 0 71232 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_627
timestamp 1698175906
transform 1 0 71568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_629
timestamp 1698175906
transform 1 0 71792 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_637
timestamp 1698175906
transform 1 0 72688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_641
timestamp 1698175906
transform 1 0 73136 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_643
timestamp 1698175906
transform 1 0 73360 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_646
timestamp 1698175906
transform 1 0 73696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_650
timestamp 1698175906
transform 1 0 74144 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_658
timestamp 1698175906
transform 1 0 75040 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_10
timestamp 1698175906
transform 1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_18
timestamp 1698175906
transform 1 0 3360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_41
timestamp 1698175906
transform 1 0 5936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_45
timestamp 1698175906
transform 1 0 6384 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_82
timestamp 1698175906
transform 1 0 10528 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_90
timestamp 1698175906
transform 1 0 11424 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_94
timestamp 1698175906
transform 1 0 11872 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_140
timestamp 1698175906
transform 1 0 17024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_144
timestamp 1698175906
transform 1 0 17472 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_146
timestamp 1698175906
transform 1 0 17696 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_149
timestamp 1698175906
transform 1 0 18032 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_157
timestamp 1698175906
transform 1 0 18928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_159
timestamp 1698175906
transform 1 0 19152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_181
timestamp 1698175906
transform 1 0 21616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_185
timestamp 1698175906
transform 1 0 22064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_189
timestamp 1698175906
transform 1 0 22512 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_193
timestamp 1698175906
transform 1 0 22960 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_211
timestamp 1698175906
transform 1 0 24976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_215
timestamp 1698175906
transform 1 0 25424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_219
timestamp 1698175906
transform 1 0 25872 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_223
timestamp 1698175906
transform 1 0 26320 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_230
timestamp 1698175906
transform 1 0 27104 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_238
timestamp 1698175906
transform 1 0 28000 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_242
timestamp 1698175906
transform 1 0 28448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698175906
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_263
timestamp 1698175906
transform 1 0 30800 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_265
timestamp 1698175906
transform 1 0 31024 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_271
timestamp 1698175906
transform 1 0 31696 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_275
timestamp 1698175906
transform 1 0 32144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_279
timestamp 1698175906
transform 1 0 32592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_310
timestamp 1698175906
transform 1 0 36064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698175906
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_326
timestamp 1698175906
transform 1 0 37856 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_328
timestamp 1698175906
transform 1 0 38080 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_358
timestamp 1698175906
transform 1 0 41440 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_362
timestamp 1698175906
transform 1 0 41888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_366
timestamp 1698175906
transform 1 0 42336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_370
timestamp 1698175906
transform 1 0 42784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_374
timestamp 1698175906
transform 1 0 43232 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_378
timestamp 1698175906
transform 1 0 43680 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_382
timestamp 1698175906
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698175906
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_402
timestamp 1698175906
transform 1 0 46368 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_410
timestamp 1698175906
transform 1 0 47264 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_463
timestamp 1698175906
transform 1 0 53200 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_467
timestamp 1698175906
transform 1 0 53648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_498
timestamp 1698175906
transform 1 0 57120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_506
timestamp 1698175906
transform 1 0 58016 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_522
timestamp 1698175906
transform 1 0 59808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_524
timestamp 1698175906
transform 1 0 60032 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_527
timestamp 1698175906
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_531
timestamp 1698175906
transform 1 0 60816 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_561
timestamp 1698175906
transform 1 0 64176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_565
timestamp 1698175906
transform 1 0 64624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_567
timestamp 1698175906
transform 1 0 64848 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_584
timestamp 1698175906
transform 1 0 66752 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_592
timestamp 1698175906
transform 1 0 67648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_594
timestamp 1698175906
transform 1 0 67872 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_597
timestamp 1698175906
transform 1 0 68208 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_633
timestamp 1698175906
transform 1 0 72240 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_637
timestamp 1698175906
transform 1 0 72688 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_654
timestamp 1698175906
transform 1 0 74592 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_662
timestamp 1698175906
transform 1 0 75488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_664
timestamp 1698175906
transform 1 0 75712 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_667
timestamp 1698175906
transform 1 0 76048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_669
timestamp 1698175906
transform 1 0 76272 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_678
timestamp 1698175906
transform 1 0 77280 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_686
timestamp 1698175906
transform 1 0 78176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_43
timestamp 1698175906
transform 1 0 6160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_47
timestamp 1698175906
transform 1 0 6608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_51
timestamp 1698175906
transform 1 0 7056 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_59
timestamp 1698175906
transform 1 0 7952 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698175906
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_80
timestamp 1698175906
transform 1 0 10304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_84
timestamp 1698175906
transform 1 0 10752 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_92
timestamp 1698175906
transform 1 0 11648 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698175906
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_147
timestamp 1698175906
transform 1 0 17808 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_151
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_155
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_163
timestamp 1698175906
transform 1 0 19600 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_172
timestamp 1698175906
transform 1 0 20608 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_178
timestamp 1698175906
transform 1 0 21280 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_184
timestamp 1698175906
transform 1 0 21952 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_188
timestamp 1698175906
transform 1 0 22400 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_192
timestamp 1698175906
transform 1 0 22848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_196
timestamp 1698175906
transform 1 0 23296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_214
timestamp 1698175906
transform 1 0 25312 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_217
timestamp 1698175906
transform 1 0 25648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_219
timestamp 1698175906
transform 1 0 25872 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_222
timestamp 1698175906
transform 1 0 26208 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_230
timestamp 1698175906
transform 1 0 27104 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_238
timestamp 1698175906
transform 1 0 28000 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_242
timestamp 1698175906
transform 1 0 28448 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_245
timestamp 1698175906
transform 1 0 28784 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_249
timestamp 1698175906
transform 1 0 29232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_296
timestamp 1698175906
transform 1 0 34496 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_312
timestamp 1698175906
transform 1 0 36288 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_320
timestamp 1698175906
transform 1 0 37184 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_324
timestamp 1698175906
transform 1 0 37632 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_327
timestamp 1698175906
transform 1 0 37968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_331
timestamp 1698175906
transform 1 0 38416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_352
timestamp 1698175906
transform 1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_356
timestamp 1698175906
transform 1 0 41216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_358
timestamp 1698175906
transform 1 0 41440 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_366
timestamp 1698175906
transform 1 0 42336 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_370
timestamp 1698175906
transform 1 0 42784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_381
timestamp 1698175906
transform 1 0 44016 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_385
timestamp 1698175906
transform 1 0 44464 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_401
timestamp 1698175906
transform 1 0 46256 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_404
timestamp 1698175906
transform 1 0 46592 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_412
timestamp 1698175906
transform 1 0 47488 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_422
timestamp 1698175906
transform 1 0 48608 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_438
timestamp 1698175906
transform 1 0 50400 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_440
timestamp 1698175906
transform 1 0 50624 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_470
timestamp 1698175906
transform 1 0 53984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_472
timestamp 1698175906
transform 1 0 54208 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_492
timestamp 1698175906
transform 1 0 56448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_496
timestamp 1698175906
transform 1 0 56896 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_500
timestamp 1698175906
transform 1 0 57344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_502
timestamp 1698175906
transform 1 0 57568 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_532
timestamp 1698175906
transform 1 0 60928 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_536
timestamp 1698175906
transform 1 0 61376 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_544
timestamp 1698175906
transform 1 0 62272 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_552
timestamp 1698175906
transform 1 0 63168 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_556
timestamp 1698175906
transform 1 0 63616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_562
timestamp 1698175906
transform 1 0 64288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_564
timestamp 1698175906
transform 1 0 64512 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_586
timestamp 1698175906
transform 1 0 66976 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_590
timestamp 1698175906
transform 1 0 67424 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_594
timestamp 1698175906
transform 1 0 67872 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_598
timestamp 1698175906
transform 1 0 68320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_602
timestamp 1698175906
transform 1 0 68768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_612
timestamp 1698175906
transform 1 0 69888 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_628
timestamp 1698175906
transform 1 0 71680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_632
timestamp 1698175906
transform 1 0 72128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_634
timestamp 1698175906
transform 1 0 72352 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_664
timestamp 1698175906
transform 1 0 75712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_668
timestamp 1698175906
transform 1 0 76160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_684
timestamp 1698175906
transform 1 0 77952 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_31
timestamp 1698175906
transform 1 0 4816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_60
timestamp 1698175906
transform 1 0 8064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_64
timestamp 1698175906
transform 1 0 8512 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_68
timestamp 1698175906
transform 1 0 8960 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_84
timestamp 1698175906
transform 1 0 10752 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_90
timestamp 1698175906
transform 1 0 11424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_98
timestamp 1698175906
transform 1 0 12320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_100
timestamp 1698175906
transform 1 0 12544 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_120
timestamp 1698175906
transform 1 0 14784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_122
timestamp 1698175906
transform 1 0 15008 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_169
timestamp 1698175906
transform 1 0 20272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_173
timestamp 1698175906
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_187
timestamp 1698175906
transform 1 0 22288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_220
timestamp 1698175906
transform 1 0 25984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_222
timestamp 1698175906
transform 1 0 26208 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_225
timestamp 1698175906
transform 1 0 26544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698175906
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_251
timestamp 1698175906
transform 1 0 29456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_255
timestamp 1698175906
transform 1 0 29904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_267
timestamp 1698175906
transform 1 0 31248 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_275
timestamp 1698175906
transform 1 0 32144 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_285
timestamp 1698175906
transform 1 0 33264 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_295
timestamp 1698175906
transform 1 0 34384 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_303
timestamp 1698175906
transform 1 0 35280 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_307
timestamp 1698175906
transform 1 0 35728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_323
timestamp 1698175906
transform 1 0 37520 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_325
timestamp 1698175906
transform 1 0 37744 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_332
timestamp 1698175906
transform 1 0 38528 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_338
timestamp 1698175906
transform 1 0 39200 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_342
timestamp 1698175906
transform 1 0 39648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_346
timestamp 1698175906
transform 1 0 40096 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_350
timestamp 1698175906
transform 1 0 40544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_368
timestamp 1698175906
transform 1 0 42560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_372
timestamp 1698175906
transform 1 0 43008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_383
timestamp 1698175906
transform 1 0 44240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_387
timestamp 1698175906
transform 1 0 44688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_391
timestamp 1698175906
transform 1 0 45136 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_399
timestamp 1698175906
transform 1 0 46032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_403
timestamp 1698175906
transform 1 0 46480 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_406
timestamp 1698175906
transform 1 0 46816 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_410
timestamp 1698175906
transform 1 0 47264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_412
timestamp 1698175906
transform 1 0 47488 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_434
timestamp 1698175906
transform 1 0 49952 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_438
timestamp 1698175906
transform 1 0 50400 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_446
timestamp 1698175906
transform 1 0 51296 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_448
timestamp 1698175906
transform 1 0 51520 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_472
timestamp 1698175906
transform 1 0 54208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_482
timestamp 1698175906
transform 1 0 55328 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_486
timestamp 1698175906
transform 1 0 55776 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_489
timestamp 1698175906
transform 1 0 56112 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_493
timestamp 1698175906
transform 1 0 56560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_497
timestamp 1698175906
transform 1 0 57008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_522
timestamp 1698175906
transform 1 0 59808 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_524
timestamp 1698175906
transform 1 0 60032 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_527
timestamp 1698175906
transform 1 0 60368 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_531
timestamp 1698175906
transform 1 0 60816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_535
timestamp 1698175906
transform 1 0 61264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_539
timestamp 1698175906
transform 1 0 61712 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_555
timestamp 1698175906
transform 1 0 63504 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_563
timestamp 1698175906
transform 1 0 64400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_565
timestamp 1698175906
transform 1 0 64624 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_597
timestamp 1698175906
transform 1 0 68208 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_629
timestamp 1698175906
transform 1 0 71792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_631
timestamp 1698175906
transform 1 0 72016 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_667
timestamp 1698175906
transform 1 0 76048 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_669
timestamp 1698175906
transform 1 0 76272 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_678
timestamp 1698175906
transform 1 0 77280 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_686
timestamp 1698175906
transform 1 0 78176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_10
timestamp 1698175906
transform 1 0 2464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_18
timestamp 1698175906
transform 1 0 3360 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_34
timestamp 1698175906
transform 1 0 5152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_65
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698175906
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_88
timestamp 1698175906
transform 1 0 11200 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_92
timestamp 1698175906
transform 1 0 11648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_94
timestamp 1698175906
transform 1 0 11872 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_162
timestamp 1698175906
transform 1 0 19488 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_193
timestamp 1698175906
transform 1 0 22960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_197
timestamp 1698175906
transform 1 0 23408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_222
timestamp 1698175906
transform 1 0 26208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_224
timestamp 1698175906
transform 1 0 26432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_251
timestamp 1698175906
transform 1 0 29456 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_267
timestamp 1698175906
transform 1 0 31248 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_271
timestamp 1698175906
transform 1 0 31696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_273
timestamp 1698175906
transform 1 0 31920 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_293
timestamp 1698175906
transform 1 0 34160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_297
timestamp 1698175906
transform 1 0 34608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_313
timestamp 1698175906
transform 1 0 36400 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_315
timestamp 1698175906
transform 1 0 36624 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_330
timestamp 1698175906
transform 1 0 38304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_352
timestamp 1698175906
transform 1 0 40768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_354
timestamp 1698175906
transform 1 0 40992 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_378
timestamp 1698175906
transform 1 0 43680 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_382
timestamp 1698175906
transform 1 0 44128 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_412
timestamp 1698175906
transform 1 0 47488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698175906
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_422
timestamp 1698175906
transform 1 0 48608 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_430
timestamp 1698175906
transform 1 0 49504 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_483
timestamp 1698175906
transform 1 0 55440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_487
timestamp 1698175906
transform 1 0 55888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_489
timestamp 1698175906
transform 1 0 56112 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_492
timestamp 1698175906
transform 1 0 56448 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_496
timestamp 1698175906
transform 1 0 56896 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_498
timestamp 1698175906
transform 1 0 57120 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_501
timestamp 1698175906
transform 1 0 57456 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_512
timestamp 1698175906
transform 1 0 58688 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_530
timestamp 1698175906
transform 1 0 60704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_534
timestamp 1698175906
transform 1 0 61152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_536
timestamp 1698175906
transform 1 0 61376 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_552
timestamp 1698175906
transform 1 0 63168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_556
timestamp 1698175906
transform 1 0 63616 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_562
timestamp 1698175906
transform 1 0 64288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_566
timestamp 1698175906
transform 1 0 64736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_570
timestamp 1698175906
transform 1 0 65184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_588
timestamp 1698175906
transform 1 0 67200 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_604
timestamp 1698175906
transform 1 0 68992 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_608
timestamp 1698175906
transform 1 0 69440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_622
timestamp 1698175906
transform 1 0 71008 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_632
timestamp 1698175906
transform 1 0 72128 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_648
timestamp 1698175906
transform 1 0 73920 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_685
timestamp 1698175906
transform 1 0 78064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_687
timestamp 1698175906
transform 1 0 78288 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_6
timestamp 1698175906
transform 1 0 2016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_14
timestamp 1698175906
transform 1 0 2912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_22
timestamp 1698175906
transform 1 0 3808 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_30
timestamp 1698175906
transform 1 0 4704 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_41
timestamp 1698175906
transform 1 0 5936 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_48
timestamp 1698175906
transform 1 0 6720 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_81
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_89
timestamp 1698175906
transform 1 0 11312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_91
timestamp 1698175906
transform 1 0 11536 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_96
timestamp 1698175906
transform 1 0 12096 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_100
timestamp 1698175906
transform 1 0 12544 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_120
timestamp 1698175906
transform 1 0 14784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_124
timestamp 1698175906
transform 1 0 15232 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_137
timestamp 1698175906
transform 1 0 16688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_160
timestamp 1698175906
transform 1 0 19264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_164
timestamp 1698175906
transform 1 0 19712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_184
timestamp 1698175906
transform 1 0 21952 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_192
timestamp 1698175906
transform 1 0 22848 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_195
timestamp 1698175906
transform 1 0 23184 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_217
timestamp 1698175906
transform 1 0 25648 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_251
timestamp 1698175906
transform 1 0 29456 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_259
timestamp 1698175906
transform 1 0 30352 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_263
timestamp 1698175906
transform 1 0 30800 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_265
timestamp 1698175906
transform 1 0 31024 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_308
timestamp 1698175906
transform 1 0 35840 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_327
timestamp 1698175906
transform 1 0 37968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_329
timestamp 1698175906
transform 1 0 38192 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_381
timestamp 1698175906
transform 1 0 44016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_387
timestamp 1698175906
transform 1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_453
timestamp 1698175906
transform 1 0 52080 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_457
timestamp 1698175906
transform 1 0 52528 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_473
timestamp 1698175906
transform 1 0 54320 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_481
timestamp 1698175906
transform 1 0 55216 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_484
timestamp 1698175906
transform 1 0 55552 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_488
timestamp 1698175906
transform 1 0 56000 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_501
timestamp 1698175906
transform 1 0 57456 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_519
timestamp 1698175906
transform 1 0 59472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_523
timestamp 1698175906
transform 1 0 59920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_527
timestamp 1698175906
transform 1 0 60368 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_529
timestamp 1698175906
transform 1 0 60592 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_559
timestamp 1698175906
transform 1 0 63952 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_588
timestamp 1698175906
transform 1 0 67200 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_592
timestamp 1698175906
transform 1 0 67648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_594
timestamp 1698175906
transform 1 0 67872 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_597
timestamp 1698175906
transform 1 0 68208 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_605
timestamp 1698175906
transform 1 0 69104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_607
timestamp 1698175906
transform 1 0 69328 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_639
timestamp 1698175906
transform 1 0 72912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_641
timestamp 1698175906
transform 1 0 73136 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_667
timestamp 1698175906
transform 1 0 76048 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_683
timestamp 1698175906
transform 1 0 77840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_687
timestamp 1698175906
transform 1 0 78288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_35
timestamp 1698175906
transform 1 0 5264 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_51
timestamp 1698175906
transform 1 0 7056 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_54
timestamp 1698175906
transform 1 0 7392 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698175906
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_87
timestamp 1698175906
transform 1 0 11088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_105
timestamp 1698175906
transform 1 0 13104 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_109
timestamp 1698175906
transform 1 0 13552 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_115
timestamp 1698175906
transform 1 0 14224 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_123
timestamp 1698175906
transform 1 0 15120 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_137
timestamp 1698175906
transform 1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698175906
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_151
timestamp 1698175906
transform 1 0 18256 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_167
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_177
timestamp 1698175906
transform 1 0 21168 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_185
timestamp 1698175906
transform 1 0 22064 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_189
timestamp 1698175906
transform 1 0 22512 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_200
timestamp 1698175906
transform 1 0 23744 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698175906
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_217
timestamp 1698175906
transform 1 0 25648 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_221
timestamp 1698175906
transform 1 0 26096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_245
timestamp 1698175906
transform 1 0 28784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_249
timestamp 1698175906
transform 1 0 29232 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_253
timestamp 1698175906
transform 1 0 29680 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_257
timestamp 1698175906
transform 1 0 30128 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698175906
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698175906
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_297
timestamp 1698175906
transform 1 0 34608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_301
timestamp 1698175906
transform 1 0 35056 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_305
timestamp 1698175906
transform 1 0 35504 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_308
timestamp 1698175906
transform 1 0 35840 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_312
timestamp 1698175906
transform 1 0 36288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_314
timestamp 1698175906
transform 1 0 36512 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_317
timestamp 1698175906
transform 1 0 36848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_321
timestamp 1698175906
transform 1 0 37296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_334
timestamp 1698175906
transform 1 0 38752 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_340
timestamp 1698175906
transform 1 0 39424 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_358
timestamp 1698175906
transform 1 0 41440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_362
timestamp 1698175906
transform 1 0 41888 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_366
timestamp 1698175906
transform 1 0 42336 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_383
timestamp 1698175906
transform 1 0 44240 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_387
timestamp 1698175906
transform 1 0 44688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_389
timestamp 1698175906
transform 1 0 44912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_396
timestamp 1698175906
transform 1 0 45696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_400
timestamp 1698175906
transform 1 0 46144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_458
timestamp 1698175906
transform 1 0 52640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_462
timestamp 1698175906
transform 1 0 53088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_466
timestamp 1698175906
transform 1 0 53536 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_476
timestamp 1698175906
transform 1 0 54656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_486
timestamp 1698175906
transform 1 0 55776 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_492
timestamp 1698175906
transform 1 0 56448 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_546
timestamp 1698175906
transform 1 0 62496 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_548
timestamp 1698175906
transform 1 0 62720 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_609
timestamp 1698175906
transform 1 0 69552 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_626
timestamp 1698175906
transform 1 0 71456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_647
timestamp 1698175906
transform 1 0 73808 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_683
timestamp 1698175906
transform 1 0 77840 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_687
timestamp 1698175906
transform 1 0 78288 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_28
timestamp 1698175906
transform 1 0 4480 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_32
timestamp 1698175906
transform 1 0 4928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_52
timestamp 1698175906
transform 1 0 7168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_60
timestamp 1698175906
transform 1 0 8064 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_92
timestamp 1698175906
transform 1 0 11648 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_96
timestamp 1698175906
transform 1 0 12096 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_100
timestamp 1698175906
transform 1 0 12544 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698175906
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_121
timestamp 1698175906
transform 1 0 14896 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_125
timestamp 1698175906
transform 1 0 15344 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_133
timestamp 1698175906
transform 1 0 16240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_135
timestamp 1698175906
transform 1 0 16464 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_145
timestamp 1698175906
transform 1 0 17584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_159
timestamp 1698175906
transform 1 0 19152 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_183
timestamp 1698175906
transform 1 0 21840 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_187
timestamp 1698175906
transform 1 0 22288 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_219
timestamp 1698175906
transform 1 0 25872 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_227
timestamp 1698175906
transform 1 0 26768 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_230
timestamp 1698175906
transform 1 0 27104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_232
timestamp 1698175906
transform 1 0 27328 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698175906
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_255
timestamp 1698175906
transform 1 0 29904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_300
timestamp 1698175906
transform 1 0 34944 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_304
timestamp 1698175906
transform 1 0 35392 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_313
timestamp 1698175906
transform 1 0 36400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_338
timestamp 1698175906
transform 1 0 39200 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_340
timestamp 1698175906
transform 1 0 39424 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_361
timestamp 1698175906
transform 1 0 41776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_365
timestamp 1698175906
transform 1 0 42224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_369
timestamp 1698175906
transform 1 0 42672 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_387
timestamp 1698175906
transform 1 0 44688 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_451
timestamp 1698175906
transform 1 0 51856 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_471
timestamp 1698175906
transform 1 0 54096 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_524
timestamp 1698175906
transform 1 0 60032 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_527
timestamp 1698175906
transform 1 0 60368 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_543
timestamp 1698175906
transform 1 0 62160 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_551
timestamp 1698175906
transform 1 0 63056 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_566
timestamp 1698175906
transform 1 0 64736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_568
timestamp 1698175906
transform 1 0 64960 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_597
timestamp 1698175906
transform 1 0 68208 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_601
timestamp 1698175906
transform 1 0 68656 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_631
timestamp 1698175906
transform 1 0 72016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_635
timestamp 1698175906
transform 1 0 72464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_679
timestamp 1698175906
transform 1 0 77392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_683
timestamp 1698175906
transform 1 0 77840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_687
timestamp 1698175906
transform 1 0 78288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_54
timestamp 1698175906
transform 1 0 7392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_58
timestamp 1698175906
transform 1 0 7840 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698175906
transform 1 0 10304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_84
timestamp 1698175906
transform 1 0 10752 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_86
timestamp 1698175906
transform 1 0 10976 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_130
timestamp 1698175906
transform 1 0 15904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_134
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_161
timestamp 1698175906
transform 1 0 19376 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_177
timestamp 1698175906
transform 1 0 21168 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_184
timestamp 1698175906
transform 1 0 21952 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_188
timestamp 1698175906
transform 1 0 22400 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_204
timestamp 1698175906
transform 1 0 24192 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_228
timestamp 1698175906
transform 1 0 26880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_232
timestamp 1698175906
transform 1 0 27328 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_257
timestamp 1698175906
transform 1 0 30128 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_261
timestamp 1698175906
transform 1 0 30576 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_264
timestamp 1698175906
transform 1 0 30912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_268
timestamp 1698175906
transform 1 0 31360 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_270
timestamp 1698175906
transform 1 0 31584 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_294
timestamp 1698175906
transform 1 0 34272 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_335
timestamp 1698175906
transform 1 0 38864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_337
timestamp 1698175906
transform 1 0 39088 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_370
timestamp 1698175906
transform 1 0 42784 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_401
timestamp 1698175906
transform 1 0 46256 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_409
timestamp 1698175906
transform 1 0 47152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_411
timestamp 1698175906
transform 1 0 47376 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_438
timestamp 1698175906
transform 1 0 50400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_442
timestamp 1698175906
transform 1 0 50848 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_455
timestamp 1698175906
transform 1 0 52304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_459
timestamp 1698175906
transform 1 0 52752 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_463
timestamp 1698175906
transform 1 0 53200 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_471
timestamp 1698175906
transform 1 0 54096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_475
timestamp 1698175906
transform 1 0 54544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_485
timestamp 1698175906
transform 1 0 55664 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_487
timestamp 1698175906
transform 1 0 55888 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_504
timestamp 1698175906
transform 1 0 57792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1698175906
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_535
timestamp 1698175906
transform 1 0 61264 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_551
timestamp 1698175906
transform 1 0 63056 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_555
timestamp 1698175906
transform 1 0 63504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_557
timestamp 1698175906
transform 1 0 63728 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_562
timestamp 1698175906
transform 1 0 64288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_564
timestamp 1698175906
transform 1 0 64512 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_578
timestamp 1698175906
transform 1 0 66080 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_595
timestamp 1698175906
transform 1 0 67984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_599
timestamp 1698175906
transform 1 0 68432 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_603
timestamp 1698175906
transform 1 0 68880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_607
timestamp 1698175906
transform 1 0 69328 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_615
timestamp 1698175906
transform 1 0 70224 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_623
timestamp 1698175906
transform 1 0 71120 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_627
timestamp 1698175906
transform 1 0 71568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_629
timestamp 1698175906
transform 1 0 71792 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_632
timestamp 1698175906
transform 1 0 72128 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_640
timestamp 1698175906
transform 1 0 73024 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_658
timestamp 1698175906
transform 1 0 75040 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_10
timestamp 1698175906
transform 1 0 2464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_14
timestamp 1698175906
transform 1 0 2912 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_16
timestamp 1698175906
transform 1 0 3136 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_29
timestamp 1698175906
transform 1 0 4592 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_33
timestamp 1698175906
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_53
timestamp 1698175906
transform 1 0 7280 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_70
timestamp 1698175906
transform 1 0 9184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_74
timestamp 1698175906
transform 1 0 9632 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_78
timestamp 1698175906
transform 1 0 10080 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_83
timestamp 1698175906
transform 1 0 10640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_98
timestamp 1698175906
transform 1 0 12320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_100
timestamp 1698175906
transform 1 0 12544 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698175906
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698175906
transform 1 0 13776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_126
timestamp 1698175906
transform 1 0 15456 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_136
timestamp 1698175906
transform 1 0 16576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_159
timestamp 1698175906
transform 1 0 19152 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_163
timestamp 1698175906
transform 1 0 19600 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_170
timestamp 1698175906
transform 1 0 20384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_181
timestamp 1698175906
transform 1 0 21616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_183
timestamp 1698175906
transform 1 0 21840 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_213
timestamp 1698175906
transform 1 0 25200 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_221
timestamp 1698175906
transform 1 0 26096 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_231
timestamp 1698175906
transform 1 0 27216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_235
timestamp 1698175906
transform 1 0 27664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_263
timestamp 1698175906
transform 1 0 30800 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_287
timestamp 1698175906
transform 1 0 33488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_291
timestamp 1698175906
transform 1 0 33936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_293
timestamp 1698175906
transform 1 0 34160 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_296
timestamp 1698175906
transform 1 0 34496 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_304
timestamp 1698175906
transform 1 0 35392 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_350
timestamp 1698175906
transform 1 0 40544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_352
timestamp 1698175906
transform 1 0 40768 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_375
timestamp 1698175906
transform 1 0 43344 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_383
timestamp 1698175906
transform 1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_409
timestamp 1698175906
transform 1 0 47152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_411
timestamp 1698175906
transform 1 0 47376 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_420
timestamp 1698175906
transform 1 0 48384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_430
timestamp 1698175906
transform 1 0 49504 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_438
timestamp 1698175906
transform 1 0 50400 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_450
timestamp 1698175906
transform 1 0 51744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_452
timestamp 1698175906
transform 1 0 51968 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_512
timestamp 1698175906
transform 1 0 58688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_516
timestamp 1698175906
transform 1 0 59136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_520
timestamp 1698175906
transform 1 0 59584 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_524
timestamp 1698175906
transform 1 0 60032 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_527
timestamp 1698175906
transform 1 0 60368 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_559
timestamp 1698175906
transform 1 0 63952 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_569
timestamp 1698175906
transform 1 0 65072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_607
timestamp 1698175906
transform 1 0 69328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_611
timestamp 1698175906
transform 1 0 69776 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_643
timestamp 1698175906
transform 1 0 73360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_655
timestamp 1698175906
transform 1 0 74704 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_663
timestamp 1698175906
transform 1 0 75600 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_667
timestamp 1698175906
transform 1 0 76048 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_669
timestamp 1698175906
transform 1 0 76272 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_678
timestamp 1698175906
transform 1 0 77280 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_686
timestamp 1698175906
transform 1 0 78176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_32
timestamp 1698175906
transform 1 0 4928 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_40
timestamp 1698175906
transform 1 0 5824 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_76
timestamp 1698175906
transform 1 0 9856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_78
timestamp 1698175906
transform 1 0 10080 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_163
timestamp 1698175906
transform 1 0 19600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_167
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_169
timestamp 1698175906
transform 1 0 20272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_172
timestamp 1698175906
transform 1 0 20608 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_188
timestamp 1698175906
transform 1 0 22400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_192
timestamp 1698175906
transform 1 0 22848 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_201
timestamp 1698175906
transform 1 0 23856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_216
timestamp 1698175906
transform 1 0 25536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_220
timestamp 1698175906
transform 1 0 25984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_224
timestamp 1698175906
transform 1 0 26432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_247
timestamp 1698175906
transform 1 0 29008 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_251
timestamp 1698175906
transform 1 0 29456 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_290
timestamp 1698175906
transform 1 0 33824 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_300
timestamp 1698175906
transform 1 0 34944 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_336
timestamp 1698175906
transform 1 0 38976 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_340
timestamp 1698175906
transform 1 0 39424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_344
timestamp 1698175906
transform 1 0 39872 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698175906
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698175906
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_385
timestamp 1698175906
transform 1 0 44464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_387
timestamp 1698175906
transform 1 0 44688 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_418
timestamp 1698175906
transform 1 0 48160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_422
timestamp 1698175906
transform 1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_426
timestamp 1698175906
transform 1 0 49056 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_430
timestamp 1698175906
transform 1 0 49504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_432
timestamp 1698175906
transform 1 0 49728 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_462
timestamp 1698175906
transform 1 0 53088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_466
timestamp 1698175906
transform 1 0 53536 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_470
timestamp 1698175906
transform 1 0 53984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_508
timestamp 1698175906
transform 1 0 58240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_512
timestamp 1698175906
transform 1 0 58688 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_528
timestamp 1698175906
transform 1 0 60480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_530
timestamp 1698175906
transform 1 0 60704 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_562
timestamp 1698175906
transform 1 0 64288 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_570
timestamp 1698175906
transform 1 0 65184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_572
timestamp 1698175906
transform 1 0 65408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_613
timestamp 1698175906
transform 1 0 70000 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_638
timestamp 1698175906
transform 1 0 72800 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_654
timestamp 1698175906
transform 1 0 74592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_685
timestamp 1698175906
transform 1 0 78064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_687
timestamp 1698175906
transform 1 0 78288 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_58
timestamp 1698175906
transform 1 0 7840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_62
timestamp 1698175906
transform 1 0 8288 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_78
timestamp 1698175906
transform 1 0 10080 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_86
timestamp 1698175906
transform 1 0 10976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_117
timestamp 1698175906
transform 1 0 14448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_121
timestamp 1698175906
transform 1 0 14896 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_160
timestamp 1698175906
transform 1 0 19264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_162
timestamp 1698175906
transform 1 0 19488 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_170
timestamp 1698175906
transform 1 0 20384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_172
timestamp 1698175906
transform 1 0 20608 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_181
timestamp 1698175906
transform 1 0 21616 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_187
timestamp 1698175906
transform 1 0 22288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_205
timestamp 1698175906
transform 1 0 24304 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_214
timestamp 1698175906
transform 1 0 25312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_218
timestamp 1698175906
transform 1 0 25760 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_232
timestamp 1698175906
transform 1 0 27328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_256
timestamp 1698175906
transform 1 0 30016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_260
timestamp 1698175906
transform 1 0 30464 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_277
timestamp 1698175906
transform 1 0 32368 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698175906
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_376
timestamp 1698175906
transform 1 0 43456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1698175906
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_389
timestamp 1698175906
transform 1 0 44912 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_404
timestamp 1698175906
transform 1 0 46592 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_426
timestamp 1698175906
transform 1 0 49056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_430
timestamp 1698175906
transform 1 0 49504 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_438
timestamp 1698175906
transform 1 0 50400 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_448
timestamp 1698175906
transform 1 0 51520 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_452
timestamp 1698175906
transform 1 0 51968 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_454
timestamp 1698175906
transform 1 0 52192 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_472
timestamp 1698175906
transform 1 0 54208 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_520
timestamp 1698175906
transform 1 0 59584 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_524
timestamp 1698175906
transform 1 0 60032 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_579
timestamp 1698175906
transform 1 0 66192 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_589
timestamp 1698175906
transform 1 0 67312 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_605
timestamp 1698175906
transform 1 0 69104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_607
timestamp 1698175906
transform 1 0 69328 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_657
timestamp 1698175906
transform 1 0 74928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_680
timestamp 1698175906
transform 1 0 77504 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_43
timestamp 1698175906
transform 1 0 6160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_47
timestamp 1698175906
transform 1 0 6608 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_63
timestamp 1698175906
transform 1 0 8400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_67
timestamp 1698175906
transform 1 0 8848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698175906
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 10304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_84
timestamp 1698175906
transform 1 0 10752 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_86
timestamp 1698175906
transform 1 0 10976 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_130
timestamp 1698175906
transform 1 0 15904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_134
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_161
timestamp 1698175906
transform 1 0 19376 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_177
timestamp 1698175906
transform 1 0 21168 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_185
timestamp 1698175906
transform 1 0 22064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_206
timestamp 1698175906
transform 1 0 24416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_216
timestamp 1698175906
transform 1 0 25536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_218
timestamp 1698175906
transform 1 0 25760 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_225
timestamp 1698175906
transform 1 0 26544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_229
timestamp 1698175906
transform 1 0 26992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_241
timestamp 1698175906
transform 1 0 28336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_245
timestamp 1698175906
transform 1 0 28784 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_262
timestamp 1698175906
transform 1 0 30688 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_290
timestamp 1698175906
transform 1 0 33824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_334
timestamp 1698175906
transform 1 0 38752 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_336
timestamp 1698175906
transform 1 0 38976 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_339
timestamp 1698175906
transform 1 0 39312 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_343
timestamp 1698175906
transform 1 0 39760 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_374
timestamp 1698175906
transform 1 0 43232 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_431
timestamp 1698175906
transform 1 0 49616 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_463
timestamp 1698175906
transform 1 0 53200 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_508
timestamp 1698175906
transform 1 0 58240 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_553
timestamp 1698175906
transform 1 0 63280 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_557
timestamp 1698175906
transform 1 0 63728 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_559
timestamp 1698175906
transform 1 0 63952 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_562
timestamp 1698175906
transform 1 0 64288 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_566
timestamp 1698175906
transform 1 0 64736 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_577
timestamp 1698175906
transform 1 0 65968 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_581
timestamp 1698175906
transform 1 0 66416 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_598
timestamp 1698175906
transform 1 0 68320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_602
timestamp 1698175906
transform 1 0 68768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_604
timestamp 1698175906
transform 1 0 68992 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_658
timestamp 1698175906
transform 1 0 75040 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_33
timestamp 1698175906
transform 1 0 5040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_72
timestamp 1698175906
transform 1 0 9408 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_80
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_99
timestamp 1698175906
transform 1 0 12432 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698175906
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_113
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_125
timestamp 1698175906
transform 1 0 15344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_127
timestamp 1698175906
transform 1 0 15568 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_159
timestamp 1698175906
transform 1 0 19152 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_167
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_171
timestamp 1698175906
transform 1 0 20496 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_179
timestamp 1698175906
transform 1 0 21392 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_188
timestamp 1698175906
transform 1 0 22400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_190
timestamp 1698175906
transform 1 0 22624 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_201
timestamp 1698175906
transform 1 0 23856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_205
timestamp 1698175906
transform 1 0 24304 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_215
timestamp 1698175906
transform 1 0 25424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_219
timestamp 1698175906
transform 1 0 25872 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_223
timestamp 1698175906
transform 1 0 26320 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_227
timestamp 1698175906
transform 1 0 26768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_240
timestamp 1698175906
transform 1 0 28224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_242
timestamp 1698175906
transform 1 0 28448 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_260
timestamp 1698175906
transform 1 0 30464 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_276
timestamp 1698175906
transform 1 0 32256 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_280
timestamp 1698175906
transform 1 0 32704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_282
timestamp 1698175906
transform 1 0 32928 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_319
timestamp 1698175906
transform 1 0 37072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_383
timestamp 1698175906
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_387
timestamp 1698175906
transform 1 0 44688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_391
timestamp 1698175906
transform 1 0 45136 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_399
timestamp 1698175906
transform 1 0 46032 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_403
timestamp 1698175906
transform 1 0 46480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_405
timestamp 1698175906
transform 1 0 46704 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_414
timestamp 1698175906
transform 1 0 47712 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_446
timestamp 1698175906
transform 1 0 51296 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_449
timestamp 1698175906
transform 1 0 51632 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_453
timestamp 1698175906
transform 1 0 52080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_486
timestamp 1698175906
transform 1 0 55776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_490
timestamp 1698175906
transform 1 0 56224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_500
timestamp 1698175906
transform 1 0 57344 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_521
timestamp 1698175906
transform 1 0 59696 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_527
timestamp 1698175906
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_531
timestamp 1698175906
transform 1 0 60816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_543
timestamp 1698175906
transform 1 0 62160 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_575
timestamp 1698175906
transform 1 0 65744 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_591
timestamp 1698175906
transform 1 0 67536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_605
timestamp 1698175906
transform 1 0 69104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_607
timestamp 1698175906
transform 1 0 69328 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_659
timestamp 1698175906
transform 1 0 75152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_687
timestamp 1698175906
transform 1 0 78288 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_10
timestamp 1698175906
transform 1 0 2464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_14
timestamp 1698175906
transform 1 0 2912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_25
timestamp 1698175906
transform 1 0 4144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_29
timestamp 1698175906
transform 1 0 4592 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_45
timestamp 1698175906
transform 1 0 6384 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_146
timestamp 1698175906
transform 1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_150
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_166
timestamp 1698175906
transform 1 0 19936 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_200
timestamp 1698175906
transform 1 0 23744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_204
timestamp 1698175906
transform 1 0 24192 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698175906
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_216
timestamp 1698175906
transform 1 0 25536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_220
timestamp 1698175906
transform 1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_232
timestamp 1698175906
transform 1 0 27328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_234
timestamp 1698175906
transform 1 0 27552 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_261
timestamp 1698175906
transform 1 0 30576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_263
timestamp 1698175906
transform 1 0 30800 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_272
timestamp 1698175906
transform 1 0 31808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_276
timestamp 1698175906
transform 1 0 32256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_319
timestamp 1698175906
transform 1 0 37072 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_321
timestamp 1698175906
transform 1 0 37296 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698175906
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_372
timestamp 1698175906
transform 1 0 43008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_376
timestamp 1698175906
transform 1 0 43456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_380
timestamp 1698175906
transform 1 0 43904 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_386
timestamp 1698175906
transform 1 0 44576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_390
timestamp 1698175906
transform 1 0 45024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_394
timestamp 1698175906
transform 1 0 45472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_398
timestamp 1698175906
transform 1 0 45920 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_414
timestamp 1698175906
transform 1 0 47712 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_418
timestamp 1698175906
transform 1 0 48160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_427
timestamp 1698175906
transform 1 0 49168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_431
timestamp 1698175906
transform 1 0 49616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_435
timestamp 1698175906
transform 1 0 50064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_439
timestamp 1698175906
transform 1 0 50512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_481
timestamp 1698175906
transform 1 0 55216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_485
timestamp 1698175906
transform 1 0 55664 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_489
timestamp 1698175906
transform 1 0 56112 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_492
timestamp 1698175906
transform 1 0 56448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_525
timestamp 1698175906
transform 1 0 60144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_529
timestamp 1698175906
transform 1 0 60592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_536
timestamp 1698175906
transform 1 0 61376 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_552
timestamp 1698175906
transform 1 0 63168 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_556
timestamp 1698175906
transform 1 0 63616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_585
timestamp 1698175906
transform 1 0 66864 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_601
timestamp 1698175906
transform 1 0 68656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_603
timestamp 1698175906
transform 1 0 68880 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_632
timestamp 1698175906
transform 1 0 72128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_53
timestamp 1698175906
transform 1 0 7280 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_55
timestamp 1698175906
transform 1 0 7504 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_62
timestamp 1698175906
transform 1 0 8288 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_70
timestamp 1698175906
transform 1 0 9184 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_74
timestamp 1698175906
transform 1 0 9632 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_94
timestamp 1698175906
transform 1 0 11872 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_102
timestamp 1698175906
transform 1 0 12768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698175906
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_145
timestamp 1698175906
transform 1 0 17584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_149
timestamp 1698175906
transform 1 0 18032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_153
timestamp 1698175906
transform 1 0 18480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_155
timestamp 1698175906
transform 1 0 18704 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_162
timestamp 1698175906
transform 1 0 19488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_166
timestamp 1698175906
transform 1 0 19936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_170
timestamp 1698175906
transform 1 0 20384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_172
timestamp 1698175906
transform 1 0 20608 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_191
timestamp 1698175906
transform 1 0 22736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_195
timestamp 1698175906
transform 1 0 23184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_199
timestamp 1698175906
transform 1 0 23632 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_203
timestamp 1698175906
transform 1 0 24080 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_206
timestamp 1698175906
transform 1 0 24416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_210
timestamp 1698175906
transform 1 0 24864 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_214
timestamp 1698175906
transform 1 0 25312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_249
timestamp 1698175906
transform 1 0 29232 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_256
timestamp 1698175906
transform 1 0 30016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_260
timestamp 1698175906
transform 1 0 30464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_264
timestamp 1698175906
transform 1 0 30912 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_268
timestamp 1698175906
transform 1 0 31360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_272
timestamp 1698175906
transform 1 0 31808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_350
timestamp 1698175906
transform 1 0 40544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_374
timestamp 1698175906
transform 1 0 43232 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_378
timestamp 1698175906
transform 1 0 43680 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_382
timestamp 1698175906
transform 1 0 44128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698175906
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_396
timestamp 1698175906
transform 1 0 45696 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_400
timestamp 1698175906
transform 1 0 46144 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_404
timestamp 1698175906
transform 1 0 46592 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_407
timestamp 1698175906
transform 1 0 46928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_411
timestamp 1698175906
transform 1 0 47376 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_415
timestamp 1698175906
transform 1 0 47824 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_419
timestamp 1698175906
transform 1 0 48272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_421
timestamp 1698175906
transform 1 0 48496 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_431
timestamp 1698175906
transform 1 0 49616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_454
timestamp 1698175906
transform 1 0 52192 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_462
timestamp 1698175906
transform 1 0 53088 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_470
timestamp 1698175906
transform 1 0 53984 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_510
timestamp 1698175906
transform 1 0 58464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_516
timestamp 1698175906
transform 1 0 59136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_520
timestamp 1698175906
transform 1 0 59584 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_524
timestamp 1698175906
transform 1 0 60032 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_527
timestamp 1698175906
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_531
timestamp 1698175906
transform 1 0 60816 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_590
timestamp 1698175906
transform 1 0 67424 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_594
timestamp 1698175906
transform 1 0 67872 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_597
timestamp 1698175906
transform 1 0 68208 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_615
timestamp 1698175906
transform 1 0 70224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_619
timestamp 1698175906
transform 1 0 70672 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_621
timestamp 1698175906
transform 1 0 70896 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_648
timestamp 1698175906
transform 1 0 73920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_652
timestamp 1698175906
transform 1 0 74368 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_662
timestamp 1698175906
transform 1 0 75488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_664
timestamp 1698175906
transform 1 0 75712 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_667
timestamp 1698175906
transform 1 0 76048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_671
timestamp 1698175906
transform 1 0 76496 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_687
timestamp 1698175906
transform 1 0 78288 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_76
timestamp 1698175906
transform 1 0 9856 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_78
timestamp 1698175906
transform 1 0 10080 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_93
timestamp 1698175906
transform 1 0 11760 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_99
timestamp 1698175906
transform 1 0 12432 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_103
timestamp 1698175906
transform 1 0 12880 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_119
timestamp 1698175906
transform 1 0 14672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_121
timestamp 1698175906
transform 1 0 14896 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_132
timestamp 1698175906
transform 1 0 16128 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698175906
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_146
timestamp 1698175906
transform 1 0 17696 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_174
timestamp 1698175906
transform 1 0 20832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_178
timestamp 1698175906
transform 1 0 21280 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_182
timestamp 1698175906
transform 1 0 21728 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_186
timestamp 1698175906
transform 1 0 22176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_190
timestamp 1698175906
transform 1 0 22624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_194
timestamp 1698175906
transform 1 0 23072 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698175906
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_228
timestamp 1698175906
transform 1 0 26880 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_239
timestamp 1698175906
transform 1 0 28112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_270
timestamp 1698175906
transform 1 0 31584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_274
timestamp 1698175906
transform 1 0 32032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_286
timestamp 1698175906
transform 1 0 33376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_328
timestamp 1698175906
transform 1 0 38080 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1698175906
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_356
timestamp 1698175906
transform 1 0 41216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_360
timestamp 1698175906
transform 1 0 41664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_364
timestamp 1698175906
transform 1 0 42112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_368
timestamp 1698175906
transform 1 0 42560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_372
timestamp 1698175906
transform 1 0 43008 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_422
timestamp 1698175906
transform 1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_426
timestamp 1698175906
transform 1 0 49056 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_435
timestamp 1698175906
transform 1 0 50064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_439
timestamp 1698175906
transform 1 0 50512 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_458
timestamp 1698175906
transform 1 0 52640 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_527
timestamp 1698175906
transform 1 0 60368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_562
timestamp 1698175906
transform 1 0 64288 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_582
timestamp 1698175906
transform 1 0 66528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_584
timestamp 1698175906
transform 1 0 66752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_590
timestamp 1698175906
transform 1 0 67424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_594
timestamp 1698175906
transform 1 0 67872 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_610
timestamp 1698175906
transform 1 0 69664 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_641
timestamp 1698175906
transform 1 0 73136 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_8
timestamp 1698175906
transform 1 0 2240 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_18
timestamp 1698175906
transform 1 0 3360 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_41
timestamp 1698175906
transform 1 0 5936 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_73
timestamp 1698175906
transform 1 0 9520 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_89
timestamp 1698175906
transform 1 0 11312 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_99
timestamp 1698175906
transform 1 0 12432 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_103
timestamp 1698175906
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_113
timestamp 1698175906
transform 1 0 14000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_117
timestamp 1698175906
transform 1 0 14448 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_144
timestamp 1698175906
transform 1 0 17472 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_157
timestamp 1698175906
transform 1 0 18928 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_163
timestamp 1698175906
transform 1 0 19600 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_167
timestamp 1698175906
transform 1 0 20048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698175906
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_181
timestamp 1698175906
transform 1 0 21616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_183
timestamp 1698175906
transform 1 0 21840 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_189
timestamp 1698175906
transform 1 0 22512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_193
timestamp 1698175906
transform 1 0 22960 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698175906
transform 1 0 25312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_257
timestamp 1698175906
transform 1 0 30128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_283
timestamp 1698175906
transform 1 0 33040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_285
timestamp 1698175906
transform 1 0 33264 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_300
timestamp 1698175906
transform 1 0 34944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_351
timestamp 1698175906
transform 1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_372
timestamp 1698175906
transform 1 0 43008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_376
timestamp 1698175906
transform 1 0 43456 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_396
timestamp 1698175906
transform 1 0 45696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_398
timestamp 1698175906
transform 1 0 45920 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_439
timestamp 1698175906
transform 1 0 50512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_451
timestamp 1698175906
transform 1 0 51856 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_457
timestamp 1698175906
transform 1 0 52528 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_465
timestamp 1698175906
transform 1 0 53424 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_469
timestamp 1698175906
transform 1 0 53872 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_471
timestamp 1698175906
transform 1 0 54096 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_524
timestamp 1698175906
transform 1 0 60032 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_536
timestamp 1698175906
transform 1 0 61376 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_573
timestamp 1698175906
transform 1 0 65520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_577
timestamp 1698175906
transform 1 0 65968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_594
timestamp 1698175906
transform 1 0 67872 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_597
timestamp 1698175906
transform 1 0 68208 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_661
timestamp 1698175906
transform 1 0 75376 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_31
timestamp 1698175906
transform 1 0 4816 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_47
timestamp 1698175906
transform 1 0 6608 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_54
timestamp 1698175906
transform 1 0 7392 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_62
timestamp 1698175906
transform 1 0 8288 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_64
timestamp 1698175906
transform 1 0 8512 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_67
timestamp 1698175906
transform 1 0 8848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698175906
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_104
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_120
timestamp 1698175906
transform 1 0 14784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_134
timestamp 1698175906
transform 1 0 16352 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698175906
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_146
timestamp 1698175906
transform 1 0 17696 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_160
timestamp 1698175906
transform 1 0 19264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_164
timestamp 1698175906
transform 1 0 19712 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_180
timestamp 1698175906
transform 1 0 21504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_182
timestamp 1698175906
transform 1 0 21728 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_194
timestamp 1698175906
transform 1 0 23072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_198
timestamp 1698175906
transform 1 0 23520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_200
timestamp 1698175906
transform 1 0 23744 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_228
timestamp 1698175906
transform 1 0 26880 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_286
timestamp 1698175906
transform 1 0 33376 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_299
timestamp 1698175906
transform 1 0 34832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_301
timestamp 1698175906
transform 1 0 35056 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_312
timestamp 1698175906
transform 1 0 36288 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_317
timestamp 1698175906
transform 1 0 36848 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_332
timestamp 1698175906
transform 1 0 38528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_334
timestamp 1698175906
transform 1 0 38752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_360
timestamp 1698175906
transform 1 0 41664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_364
timestamp 1698175906
transform 1 0 42112 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_373
timestamp 1698175906
transform 1 0 43120 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_377
timestamp 1698175906
transform 1 0 43568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_381
timestamp 1698175906
transform 1 0 44016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_387
timestamp 1698175906
transform 1 0 44688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_389
timestamp 1698175906
transform 1 0 44912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_392
timestamp 1698175906
transform 1 0 45248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_402
timestamp 1698175906
transform 1 0 46368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_406
timestamp 1698175906
transform 1 0 46816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_414
timestamp 1698175906
transform 1 0 47712 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_418
timestamp 1698175906
transform 1 0 48160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_422
timestamp 1698175906
transform 1 0 48608 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_426
timestamp 1698175906
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_428
timestamp 1698175906
transform 1 0 49280 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_431
timestamp 1698175906
transform 1 0 49616 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_433
timestamp 1698175906
transform 1 0 49840 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_454
timestamp 1698175906
transform 1 0 52192 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_537
timestamp 1698175906
transform 1 0 61488 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_541
timestamp 1698175906
transform 1 0 61936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_545
timestamp 1698175906
transform 1 0 62384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_549
timestamp 1698175906
transform 1 0 62832 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_555
timestamp 1698175906
transform 1 0 63504 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_559
timestamp 1698175906
transform 1 0 63952 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_562
timestamp 1698175906
transform 1 0 64288 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_566
timestamp 1698175906
transform 1 0 64736 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_568
timestamp 1698175906
transform 1 0 64960 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_571
timestamp 1698175906
transform 1 0 65296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_573
timestamp 1698175906
transform 1 0 65520 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_605
timestamp 1698175906
transform 1 0 69104 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_613
timestamp 1698175906
transform 1 0 70000 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_632
timestamp 1698175906
transform 1 0 72128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_634
timestamp 1698175906
transform 1 0 72352 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_687
timestamp 1698175906
transform 1 0 78288 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_82
timestamp 1698175906
transform 1 0 10528 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_86
timestamp 1698175906
transform 1 0 10976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_94
timestamp 1698175906
transform 1 0 11872 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_102
timestamp 1698175906
transform 1 0 12768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698175906
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_111
timestamp 1698175906
transform 1 0 13776 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_119
timestamp 1698175906
transform 1 0 14672 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_123
timestamp 1698175906
transform 1 0 15120 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_169
timestamp 1698175906
transform 1 0 20272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_198
timestamp 1698175906
transform 1 0 23520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_202
timestamp 1698175906
transform 1 0 23968 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_210
timestamp 1698175906
transform 1 0 24864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_212
timestamp 1698175906
transform 1 0 25088 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_215
timestamp 1698175906
transform 1 0 25424 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_231
timestamp 1698175906
transform 1 0 27216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_235
timestamp 1698175906
transform 1 0 27664 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_256
timestamp 1698175906
transform 1 0 30016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_260
timestamp 1698175906
transform 1 0 30464 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_263
timestamp 1698175906
transform 1 0 30800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_297
timestamp 1698175906
transform 1 0 34608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_299
timestamp 1698175906
transform 1 0 34832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_380
timestamp 1698175906
transform 1 0 43904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698175906
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_387
timestamp 1698175906
transform 1 0 44688 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_391
timestamp 1698175906
transform 1 0 45136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_395
timestamp 1698175906
transform 1 0 45584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_397
timestamp 1698175906
transform 1 0 45808 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_400
timestamp 1698175906
transform 1 0 46144 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_431
timestamp 1698175906
transform 1 0 49616 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_439
timestamp 1698175906
transform 1 0 50512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_442
timestamp 1698175906
transform 1 0 50848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_450
timestamp 1698175906
transform 1 0 51744 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_452
timestamp 1698175906
transform 1 0 51968 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_457
timestamp 1698175906
transform 1 0 52528 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_522
timestamp 1698175906
transform 1 0 59808 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_524
timestamp 1698175906
transform 1 0 60032 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_527
timestamp 1698175906
transform 1 0 60368 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_531
timestamp 1698175906
transform 1 0 60816 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_547
timestamp 1698175906
transform 1 0 62608 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_555
timestamp 1698175906
transform 1 0 63504 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_559
timestamp 1698175906
transform 1 0 63952 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_563
timestamp 1698175906
transform 1 0 64400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_567
timestamp 1698175906
transform 1 0 64848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_575
timestamp 1698175906
transform 1 0 65744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_579
timestamp 1698175906
transform 1 0 66192 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_586
timestamp 1698175906
transform 1 0 66976 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_594
timestamp 1698175906
transform 1 0 67872 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_597
timestamp 1698175906
transform 1 0 68208 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_601
timestamp 1698175906
transform 1 0 68656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_603
timestamp 1698175906
transform 1 0 68880 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_629
timestamp 1698175906
transform 1 0 71792 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_667
timestamp 1698175906
transform 1 0 76048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_669
timestamp 1698175906
transform 1 0 76272 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_672
timestamp 1698175906
transform 1 0 76608 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_18
timestamp 1698175906
transform 1 0 3360 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_34
timestamp 1698175906
transform 1 0 5152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_42
timestamp 1698175906
transform 1 0 6048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_46
timestamp 1698175906
transform 1 0 6496 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_62
timestamp 1698175906
transform 1 0 8288 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_78
timestamp 1698175906
transform 1 0 10080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_166
timestamp 1698175906
transform 1 0 19936 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_216
timestamp 1698175906
transform 1 0 25536 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_218
timestamp 1698175906
transform 1 0 25760 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_221
timestamp 1698175906
transform 1 0 26096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_225
timestamp 1698175906
transform 1 0 26544 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_228
timestamp 1698175906
transform 1 0 26880 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_232
timestamp 1698175906
transform 1 0 27328 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_249
timestamp 1698175906
transform 1 0 29232 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_251
timestamp 1698175906
transform 1 0 29456 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_260
timestamp 1698175906
transform 1 0 30464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_264
timestamp 1698175906
transform 1 0 30912 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_268
timestamp 1698175906
transform 1 0 31360 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_270
timestamp 1698175906
transform 1 0 31584 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_328
timestamp 1698175906
transform 1 0 38080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_332
timestamp 1698175906
transform 1 0 38528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698175906
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_352
timestamp 1698175906
transform 1 0 40768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_354
timestamp 1698175906
transform 1 0 40992 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_372
timestamp 1698175906
transform 1 0 43008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_376
timestamp 1698175906
transform 1 0 43456 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_380
timestamp 1698175906
transform 1 0 43904 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_408
timestamp 1698175906
transform 1 0 47040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_410
timestamp 1698175906
transform 1 0 47264 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_413
timestamp 1698175906
transform 1 0 47600 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_417
timestamp 1698175906
transform 1 0 48048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_419
timestamp 1698175906
transform 1 0 48272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_422
timestamp 1698175906
transform 1 0 48608 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_426
timestamp 1698175906
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_428
timestamp 1698175906
transform 1 0 49280 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_431
timestamp 1698175906
transform 1 0 49616 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_439
timestamp 1698175906
transform 1 0 50512 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_451
timestamp 1698175906
transform 1 0 51856 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_455
timestamp 1698175906
transform 1 0 52304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_457
timestamp 1698175906
transform 1 0 52528 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_478
timestamp 1698175906
transform 1 0 54880 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_500
timestamp 1698175906
transform 1 0 57344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_502
timestamp 1698175906
transform 1 0 57568 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_511
timestamp 1698175906
transform 1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_515
timestamp 1698175906
transform 1 0 59024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_519
timestamp 1698175906
transform 1 0 59472 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_529
timestamp 1698175906
transform 1 0 60592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_533
timestamp 1698175906
transform 1 0 61040 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_541
timestamp 1698175906
transform 1 0 61936 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_550
timestamp 1698175906
transform 1 0 62944 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_562
timestamp 1698175906
transform 1 0 64288 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_564
timestamp 1698175906
transform 1 0 64512 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_580
timestamp 1698175906
transform 1 0 66304 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_596
timestamp 1698175906
transform 1 0 68096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_598
timestamp 1698175906
transform 1 0 68320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_615
timestamp 1698175906
transform 1 0 70224 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_623
timestamp 1698175906
transform 1 0 71120 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_627
timestamp 1698175906
transform 1 0 71568 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_657
timestamp 1698175906
transform 1 0 74928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_69
timestamp 1698175906
transform 1 0 9072 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_77
timestamp 1698175906
transform 1 0 9968 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_80
timestamp 1698175906
transform 1 0 10304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_82
timestamp 1698175906
transform 1 0 10528 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_89
timestamp 1698175906
transform 1 0 11312 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_111
timestamp 1698175906
transform 1 0 13776 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_162
timestamp 1698175906
transform 1 0 19488 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_225
timestamp 1698175906
transform 1 0 26544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_241
timestamp 1698175906
transform 1 0 28336 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_252
timestamp 1698175906
transform 1 0 29568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_256
timestamp 1698175906
transform 1 0 30016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_260
timestamp 1698175906
transform 1 0 30464 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_276
timestamp 1698175906
transform 1 0 32256 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_280
timestamp 1698175906
transform 1 0 32704 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_284
timestamp 1698175906
transform 1 0 33152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_293
timestamp 1698175906
transform 1 0 34160 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_305
timestamp 1698175906
transform 1 0 35504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698175906
transform 1 0 35952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698175906
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_325
timestamp 1698175906
transform 1 0 37744 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_339
timestamp 1698175906
transform 1 0 39312 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_350
timestamp 1698175906
transform 1 0 40544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_354
timestamp 1698175906
transform 1 0 40992 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_358
timestamp 1698175906
transform 1 0 41440 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_362
timestamp 1698175906
transform 1 0 41888 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_378
timestamp 1698175906
transform 1 0 43680 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_381
timestamp 1698175906
transform 1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_387
timestamp 1698175906
transform 1 0 44688 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_396
timestamp 1698175906
transform 1 0 45696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_400
timestamp 1698175906
transform 1 0 46144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_412
timestamp 1698175906
transform 1 0 47488 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_443
timestamp 1698175906
transform 1 0 50960 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_451
timestamp 1698175906
transform 1 0 51856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_457
timestamp 1698175906
transform 1 0 52528 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_461
timestamp 1698175906
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_479
timestamp 1698175906
transform 1 0 54992 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_506
timestamp 1698175906
transform 1 0 58016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_510
timestamp 1698175906
transform 1 0 58464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_512
timestamp 1698175906
transform 1 0 58688 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_527
timestamp 1698175906
transform 1 0 60368 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_543
timestamp 1698175906
transform 1 0 62160 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_551
timestamp 1698175906
transform 1 0 63056 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_581
timestamp 1698175906
transform 1 0 66416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_585
timestamp 1698175906
transform 1 0 66864 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_613
timestamp 1698175906
transform 1 0 70000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_615
timestamp 1698175906
transform 1 0 70224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_663
timestamp 1698175906
transform 1 0 75600 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_682
timestamp 1698175906
transform 1 0 77728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_686
timestamp 1698175906
transform 1 0 78176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_31
timestamp 1698175906
transform 1 0 4816 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_47
timestamp 1698175906
transform 1 0 6608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_76
timestamp 1698175906
transform 1 0 9856 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_84
timestamp 1698175906
transform 1 0 10752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_91
timestamp 1698175906
transform 1 0 11536 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_95
timestamp 1698175906
transform 1 0 11984 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_111
timestamp 1698175906
transform 1 0 13776 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_119
timestamp 1698175906
transform 1 0 14672 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_144
timestamp 1698175906
transform 1 0 17472 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_163
timestamp 1698175906
transform 1 0 19600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_167
timestamp 1698175906
transform 1 0 20048 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_192
timestamp 1698175906
transform 1 0 22848 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_196
timestamp 1698175906
transform 1 0 23296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_216
timestamp 1698175906
transform 1 0 25536 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_240
timestamp 1698175906
transform 1 0 28224 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_257
timestamp 1698175906
transform 1 0 30128 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_261
timestamp 1698175906
transform 1 0 30576 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_273
timestamp 1698175906
transform 1 0 31920 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_319
timestamp 1698175906
transform 1 0 37072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_352
timestamp 1698175906
transform 1 0 40768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_360
timestamp 1698175906
transform 1 0 41664 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_364
timestamp 1698175906
transform 1 0 42112 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_373
timestamp 1698175906
transform 1 0 43120 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_377
timestamp 1698175906
transform 1 0 43568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_385
timestamp 1698175906
transform 1 0 44464 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_404
timestamp 1698175906
transform 1 0 46592 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_412
timestamp 1698175906
transform 1 0 47488 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_416
timestamp 1698175906
transform 1 0 47936 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_446
timestamp 1698175906
transform 1 0 51296 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_454
timestamp 1698175906
transform 1 0 52192 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_464
timestamp 1698175906
transform 1 0 53312 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_468
timestamp 1698175906
transform 1 0 53760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_470
timestamp 1698175906
transform 1 0 53984 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_473
timestamp 1698175906
transform 1 0 54320 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_489
timestamp 1698175906
transform 1 0 56112 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_492
timestamp 1698175906
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_496
timestamp 1698175906
transform 1 0 56896 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_502
timestamp 1698175906
transform 1 0 57568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_526
timestamp 1698175906
transform 1 0 60256 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_534
timestamp 1698175906
transform 1 0 61152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_536
timestamp 1698175906
transform 1 0 61376 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_543
timestamp 1698175906
transform 1 0 62160 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_556
timestamp 1698175906
transform 1 0 63616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_562
timestamp 1698175906
transform 1 0 64288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_648
timestamp 1698175906
transform 1 0 73920 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_678
timestamp 1698175906
transform 1 0 77280 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_686
timestamp 1698175906
transform 1 0 78176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_10
timestamp 1698175906
transform 1 0 2464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_18
timestamp 1698175906
transform 1 0 3360 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_26
timestamp 1698175906
transform 1 0 4256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_30
timestamp 1698175906
transform 1 0 4704 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_45
timestamp 1698175906
transform 1 0 6384 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_75
timestamp 1698175906
transform 1 0 9744 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_123
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_131
timestamp 1698175906
transform 1 0 16016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_133
timestamp 1698175906
transform 1 0 16240 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_136
timestamp 1698175906
transform 1 0 16576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_148
timestamp 1698175906
transform 1 0 17920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_156
timestamp 1698175906
transform 1 0 18816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_160
timestamp 1698175906
transform 1 0 19264 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_168
timestamp 1698175906
transform 1 0 20160 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698175906
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_184
timestamp 1698175906
transform 1 0 21952 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_188
timestamp 1698175906
transform 1 0 22400 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_194
timestamp 1698175906
transform 1 0 23072 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_202
timestamp 1698175906
transform 1 0 23968 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_255
timestamp 1698175906
transform 1 0 29904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_349
timestamp 1698175906
transform 1 0 40432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_353
timestamp 1698175906
transform 1 0 40880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_355
timestamp 1698175906
transform 1 0 41104 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_358
timestamp 1698175906
transform 1 0 41440 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_362
timestamp 1698175906
transform 1 0 41888 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_399
timestamp 1698175906
transform 1 0 46032 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_415
timestamp 1698175906
transform 1 0 47824 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_419
timestamp 1698175906
transform 1 0 48272 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_422
timestamp 1698175906
transform 1 0 48608 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_430
timestamp 1698175906
transform 1 0 49504 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_434
timestamp 1698175906
transform 1 0 49952 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_436
timestamp 1698175906
transform 1 0 50176 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_439
timestamp 1698175906
transform 1 0 50512 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_457
timestamp 1698175906
transform 1 0 52528 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_476
timestamp 1698175906
transform 1 0 54656 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_508
timestamp 1698175906
transform 1 0 58240 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_524
timestamp 1698175906
transform 1 0 60032 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_527
timestamp 1698175906
transform 1 0 60368 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_531
timestamp 1698175906
transform 1 0 60816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_533
timestamp 1698175906
transform 1 0 61040 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_549
timestamp 1698175906
transform 1 0 62832 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_565
timestamp 1698175906
transform 1 0 64624 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_573
timestamp 1698175906
transform 1 0 65520 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_577
timestamp 1698175906
transform 1 0 65968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_649
timestamp 1698175906
transform 1 0 74032 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_673
timestamp 1698175906
transform 1 0 76720 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_681
timestamp 1698175906
transform 1 0 77616 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_685
timestamp 1698175906
transform 1 0 78064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_687
timestamp 1698175906
transform 1 0 78288 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_43
timestamp 1698175906
transform 1 0 6160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_47
timestamp 1698175906
transform 1 0 6608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_51
timestamp 1698175906
transform 1 0 7056 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_67
timestamp 1698175906
transform 1 0 8848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698175906
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_87
timestamp 1698175906
transform 1 0 11088 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_94
timestamp 1698175906
transform 1 0 11872 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_98
timestamp 1698175906
transform 1 0 12320 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_114
timestamp 1698175906
transform 1 0 14112 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_118
timestamp 1698175906
transform 1 0 14560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_120
timestamp 1698175906
transform 1 0 14784 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_129
timestamp 1698175906
transform 1 0 15792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_131
timestamp 1698175906
transform 1 0 16016 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_157
timestamp 1698175906
transform 1 0 18928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_178
timestamp 1698175906
transform 1 0 21280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_180
timestamp 1698175906
transform 1 0 21504 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_185
timestamp 1698175906
transform 1 0 22064 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_189
timestamp 1698175906
transform 1 0 22512 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_199
timestamp 1698175906
transform 1 0 23632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_201
timestamp 1698175906
transform 1 0 23856 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_225
timestamp 1698175906
transform 1 0 26544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_229
timestamp 1698175906
transform 1 0 26992 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_233
timestamp 1698175906
transform 1 0 27440 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_235
timestamp 1698175906
transform 1 0 27664 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_241
timestamp 1698175906
transform 1 0 28336 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_245
timestamp 1698175906
transform 1 0 28784 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_249
timestamp 1698175906
transform 1 0 29232 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_302
timestamp 1698175906
transform 1 0 35168 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_306
timestamp 1698175906
transform 1 0 35616 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_314
timestamp 1698175906
transform 1 0 36512 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_318
timestamp 1698175906
transform 1 0 36960 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698175906
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_352
timestamp 1698175906
transform 1 0 40768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_354
timestamp 1698175906
transform 1 0 40992 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_360
timestamp 1698175906
transform 1 0 41664 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_364
timestamp 1698175906
transform 1 0 42112 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_366
timestamp 1698175906
transform 1 0 42336 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_372
timestamp 1698175906
transform 1 0 43008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_376
timestamp 1698175906
transform 1 0 43456 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_387
timestamp 1698175906
transform 1 0 44688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_391
timestamp 1698175906
transform 1 0 45136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_395
timestamp 1698175906
transform 1 0 45584 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_403
timestamp 1698175906
transform 1 0 46480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_422
timestamp 1698175906
transform 1 0 48608 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_429
timestamp 1698175906
transform 1 0 49392 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_445
timestamp 1698175906
transform 1 0 51184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_473
timestamp 1698175906
transform 1 0 54320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_483
timestamp 1698175906
transform 1 0 55440 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_487
timestamp 1698175906
transform 1 0 55888 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_489
timestamp 1698175906
transform 1 0 56112 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_492
timestamp 1698175906
transform 1 0 56448 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_496
timestamp 1698175906
transform 1 0 56896 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_504
timestamp 1698175906
transform 1 0 57792 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698175906
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_522
timestamp 1698175906
transform 1 0 59808 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_538
timestamp 1698175906
transform 1 0 61600 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_555
timestamp 1698175906
transform 1 0 63504 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_559
timestamp 1698175906
transform 1 0 63952 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_562
timestamp 1698175906
transform 1 0 64288 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_594
timestamp 1698175906
transform 1 0 67872 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_607
timestamp 1698175906
transform 1 0 69328 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_611
timestamp 1698175906
transform 1 0 69776 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_629
timestamp 1698175906
transform 1 0 71792 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_648
timestamp 1698175906
transform 1 0 73920 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_652
timestamp 1698175906
transform 1 0 74368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_660
timestamp 1698175906
transform 1 0 75264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_43
timestamp 1698175906
transform 1 0 6160 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_47
timestamp 1698175906
transform 1 0 6608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_49
timestamp 1698175906
transform 1 0 6832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_79
timestamp 1698175906
transform 1 0 10192 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_89
timestamp 1698175906
transform 1 0 11312 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_211
timestamp 1698175906
transform 1 0 24976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_213
timestamp 1698175906
transform 1 0 25200 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_220
timestamp 1698175906
transform 1 0 25984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_232
timestamp 1698175906
transform 1 0 27328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_234
timestamp 1698175906
transform 1 0 27552 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_305
timestamp 1698175906
transform 1 0 35504 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_307
timestamp 1698175906
transform 1 0 35728 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_364
timestamp 1698175906
transform 1 0 42112 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_368
timestamp 1698175906
transform 1 0 42560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_372
timestamp 1698175906
transform 1 0 43008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_380
timestamp 1698175906
transform 1 0 43904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698175906
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_387
timestamp 1698175906
transform 1 0 44688 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_395
timestamp 1698175906
transform 1 0 45584 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_406
timestamp 1698175906
transform 1 0 46816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_408
timestamp 1698175906
transform 1 0 47040 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_422
timestamp 1698175906
transform 1 0 48608 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_430
timestamp 1698175906
transform 1 0 49504 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_466
timestamp 1698175906
transform 1 0 53536 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_481
timestamp 1698175906
transform 1 0 55216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_483
timestamp 1698175906
transform 1 0 55440 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_492
timestamp 1698175906
transform 1 0 56448 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_527
timestamp 1698175906
transform 1 0 60368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_549
timestamp 1698175906
transform 1 0 62832 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_565
timestamp 1698175906
transform 1 0 64624 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_573
timestamp 1698175906
transform 1 0 65520 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_575
timestamp 1698175906
transform 1 0 65744 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_593
timestamp 1698175906
transform 1 0 67760 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_597
timestamp 1698175906
transform 1 0 68208 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_629
timestamp 1698175906
transform 1 0 71792 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_632
timestamp 1698175906
transform 1 0 72128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_636
timestamp 1698175906
transform 1 0 72576 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_667
timestamp 1698175906
transform 1 0 76048 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_671
timestamp 1698175906
transform 1 0 76496 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_687
timestamp 1698175906
transform 1 0 78288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_6
timestamp 1698175906
transform 1 0 2016 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_52
timestamp 1698175906
transform 1 0 7168 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_56
timestamp 1698175906
transform 1 0 7616 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_64
timestamp 1698175906
transform 1 0 8512 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698175906
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_87
timestamp 1698175906
transform 1 0 11088 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_91
timestamp 1698175906
transform 1 0 11536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_95
timestamp 1698175906
transform 1 0 11984 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_103
timestamp 1698175906
transform 1 0 12880 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698175906
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_150
timestamp 1698175906
transform 1 0 18144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_162
timestamp 1698175906
transform 1 0 19488 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_166
timestamp 1698175906
transform 1 0 19936 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_214
timestamp 1698175906
transform 1 0 25312 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_240
timestamp 1698175906
transform 1 0 28224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_244
timestamp 1698175906
transform 1 0 28672 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698175906
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_295
timestamp 1698175906
transform 1 0 34384 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_299
timestamp 1698175906
transform 1 0 34832 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_326
timestamp 1698175906
transform 1 0 37856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_328
timestamp 1698175906
transform 1 0 38080 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_352
timestamp 1698175906
transform 1 0 40768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_354
timestamp 1698175906
transform 1 0 40992 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_357
timestamp 1698175906
transform 1 0 41328 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_361
timestamp 1698175906
transform 1 0 41776 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_385
timestamp 1698175906
transform 1 0 44464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_389
timestamp 1698175906
transform 1 0 44912 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_393
timestamp 1698175906
transform 1 0 45360 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_395
timestamp 1698175906
transform 1 0 45584 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698175906
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_435
timestamp 1698175906
transform 1 0 50064 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_443
timestamp 1698175906
transform 1 0 50960 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_456
timestamp 1698175906
transform 1 0 52416 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_458
timestamp 1698175906
transform 1 0 52640 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_487
timestamp 1698175906
transform 1 0 55888 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_489
timestamp 1698175906
transform 1 0 56112 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_492
timestamp 1698175906
transform 1 0 56448 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_500
timestamp 1698175906
transform 1 0 57344 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_525
timestamp 1698175906
transform 1 0 60144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_529
timestamp 1698175906
transform 1 0 60592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_553
timestamp 1698175906
transform 1 0 63280 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_557
timestamp 1698175906
transform 1 0 63728 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_559
timestamp 1698175906
transform 1 0 63952 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_562
timestamp 1698175906
transform 1 0 64288 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_564
timestamp 1698175906
transform 1 0 64512 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_592
timestamp 1698175906
transform 1 0 67648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_596
timestamp 1698175906
transform 1 0 68096 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_604
timestamp 1698175906
transform 1 0 68992 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_608
timestamp 1698175906
transform 1 0 69440 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_627
timestamp 1698175906
transform 1 0 71568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_629
timestamp 1698175906
transform 1 0 71792 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_638
timestamp 1698175906
transform 1 0 72800 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_646
timestamp 1698175906
transform 1 0 73696 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_684
timestamp 1698175906
transform 1 0 77952 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_10
timestamp 1698175906
transform 1 0 2464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_14
timestamp 1698175906
transform 1 0 2912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_16
timestamp 1698175906
transform 1 0 3136 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_23
timestamp 1698175906
transform 1 0 3920 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_31
timestamp 1698175906
transform 1 0 4816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_41
timestamp 1698175906
transform 1 0 5936 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_57
timestamp 1698175906
transform 1 0 7728 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_61
timestamp 1698175906
transform 1 0 8176 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_91
timestamp 1698175906
transform 1 0 11536 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_99
timestamp 1698175906
transform 1 0 12432 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698175906
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_151
timestamp 1698175906
transform 1 0 18256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_153
timestamp 1698175906
transform 1 0 18480 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_173
timestamp 1698175906
transform 1 0 20720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_179
timestamp 1698175906
transform 1 0 21392 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_223
timestamp 1698175906
transform 1 0 26320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_227
timestamp 1698175906
transform 1 0 26768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_304
timestamp 1698175906
transform 1 0 35392 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_306
timestamp 1698175906
transform 1 0 35616 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_366
timestamp 1698175906
transform 1 0 42336 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_370
timestamp 1698175906
transform 1 0 42784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_374
timestamp 1698175906
transform 1 0 43232 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698175906
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_387
timestamp 1698175906
transform 1 0 44688 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_394
timestamp 1698175906
transform 1 0 45472 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_398
timestamp 1698175906
transform 1 0 45920 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_402
timestamp 1698175906
transform 1 0 46368 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_419
timestamp 1698175906
transform 1 0 48272 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698175906
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_457
timestamp 1698175906
transform 1 0 52528 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_473
timestamp 1698175906
transform 1 0 54320 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_489
timestamp 1698175906
transform 1 0 56112 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_493
timestamp 1698175906
transform 1 0 56560 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_496
timestamp 1698175906
transform 1 0 56896 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_500
timestamp 1698175906
transform 1 0 57344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_544
timestamp 1698175906
transform 1 0 62272 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_560
timestamp 1698175906
transform 1 0 64064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_562
timestamp 1698175906
transform 1 0 64288 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_594
timestamp 1698175906
transform 1 0 67872 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_649
timestamp 1698175906
transform 1 0 74032 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_682
timestamp 1698175906
transform 1 0 77728 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_686
timestamp 1698175906
transform 1 0 78176 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_78
timestamp 1698175906
transform 1 0 10080 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_110
timestamp 1698175906
transform 1 0 13664 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_144
timestamp 1698175906
transform 1 0 17472 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_171
timestamp 1698175906
transform 1 0 20496 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_175
timestamp 1698175906
transform 1 0 20944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_177
timestamp 1698175906
transform 1 0 21168 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_247
timestamp 1698175906
transform 1 0 29008 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_251
timestamp 1698175906
transform 1 0 29456 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_272
timestamp 1698175906
transform 1 0 31808 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_288
timestamp 1698175906
transform 1 0 33600 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_298
timestamp 1698175906
transform 1 0 34720 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_352
timestamp 1698175906
transform 1 0 40768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_356
timestamp 1698175906
transform 1 0 41216 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_360
timestamp 1698175906
transform 1 0 41664 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_371
timestamp 1698175906
transform 1 0 42896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_375
timestamp 1698175906
transform 1 0 43344 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_384
timestamp 1698175906
transform 1 0 44352 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_388
timestamp 1698175906
transform 1 0 44800 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_404
timestamp 1698175906
transform 1 0 46592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_408
timestamp 1698175906
transform 1 0 47040 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_410
timestamp 1698175906
transform 1 0 47264 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_419
timestamp 1698175906
transform 1 0 48272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_422
timestamp 1698175906
transform 1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_424
timestamp 1698175906
transform 1 0 48832 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_432
timestamp 1698175906
transform 1 0 49728 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_455
timestamp 1698175906
transform 1 0 52304 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_487
timestamp 1698175906
transform 1 0 55888 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_489
timestamp 1698175906
transform 1 0 56112 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_492
timestamp 1698175906
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_496
timestamp 1698175906
transform 1 0 56896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_508
timestamp 1698175906
transform 1 0 58240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_512
timestamp 1698175906
transform 1 0 58688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_525
timestamp 1698175906
transform 1 0 60144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_529
timestamp 1698175906
transform 1 0 60592 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_545
timestamp 1698175906
transform 1 0 62384 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_553
timestamp 1698175906
transform 1 0 63280 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_557
timestamp 1698175906
transform 1 0 63728 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_559
timestamp 1698175906
transform 1 0 63952 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_562
timestamp 1698175906
transform 1 0 64288 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_593
timestamp 1698175906
transform 1 0 67760 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_597
timestamp 1698175906
transform 1 0 68208 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_605
timestamp 1698175906
transform 1 0 69104 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_609
timestamp 1698175906
transform 1 0 69552 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_616
timestamp 1698175906
transform 1 0 70336 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_620
timestamp 1698175906
transform 1 0 70784 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_627
timestamp 1698175906
transform 1 0 71568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_629
timestamp 1698175906
transform 1 0 71792 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_632
timestamp 1698175906
transform 1 0 72128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_636
timestamp 1698175906
transform 1 0 72576 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_644
timestamp 1698175906
transform 1 0 73472 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_648
timestamp 1698175906
transform 1 0 73920 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_684
timestamp 1698175906
transform 1 0 77952 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_28
timestamp 1698175906
transform 1 0 4480 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_32
timestamp 1698175906
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_53
timestamp 1698175906
transform 1 0 7280 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_61
timestamp 1698175906
transform 1 0 8176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_63
timestamp 1698175906
transform 1 0 8400 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_70
timestamp 1698175906
transform 1 0 9184 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_74
timestamp 1698175906
transform 1 0 9632 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_90
timestamp 1698175906
transform 1 0 11424 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_98
timestamp 1698175906
transform 1 0 12320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_102
timestamp 1698175906
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698175906
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_125
timestamp 1698175906
transform 1 0 15344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_127
timestamp 1698175906
transform 1 0 15568 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_134
timestamp 1698175906
transform 1 0 16352 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_142
timestamp 1698175906
transform 1 0 17248 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_181
timestamp 1698175906
transform 1 0 21616 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_194
timestamp 1698175906
transform 1 0 23072 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_213
timestamp 1698175906
transform 1 0 25200 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_217
timestamp 1698175906
transform 1 0 25648 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_237
timestamp 1698175906
transform 1 0 27888 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_261
timestamp 1698175906
transform 1 0 30576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_290
timestamp 1698175906
transform 1 0 33824 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_306
timestamp 1698175906
transform 1 0 35616 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698175906
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_325
timestamp 1698175906
transform 1 0 37744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_369
timestamp 1698175906
transform 1 0 42672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_378
timestamp 1698175906
transform 1 0 43680 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_382
timestamp 1698175906
transform 1 0 44128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698175906
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_391
timestamp 1698175906
transform 1 0 45136 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_395
timestamp 1698175906
transform 1 0 45584 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_407
timestamp 1698175906
transform 1 0 46928 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_415
timestamp 1698175906
transform 1 0 47824 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_419
timestamp 1698175906
transform 1 0 48272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_427
timestamp 1698175906
transform 1 0 49168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_429
timestamp 1698175906
transform 1 0 49392 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_438
timestamp 1698175906
transform 1 0 50400 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_444
timestamp 1698175906
transform 1 0 51072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_454
timestamp 1698175906
transform 1 0 52192 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_457
timestamp 1698175906
transform 1 0 52528 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_461
timestamp 1698175906
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_471
timestamp 1698175906
transform 1 0 54096 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_503
timestamp 1698175906
transform 1 0 57680 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_511
timestamp 1698175906
transform 1 0 58576 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_514
timestamp 1698175906
transform 1 0 58912 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_518
timestamp 1698175906
transform 1 0 59360 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_522
timestamp 1698175906
transform 1 0 59808 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_524
timestamp 1698175906
transform 1 0 60032 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_527
timestamp 1698175906
transform 1 0 60368 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_540
timestamp 1698175906
transform 1 0 61824 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_556
timestamp 1698175906
transform 1 0 63616 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_564
timestamp 1698175906
transform 1 0 64512 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_578
timestamp 1698175906
transform 1 0 66080 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_582
timestamp 1698175906
transform 1 0 66528 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_590
timestamp 1698175906
transform 1 0 67424 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_594
timestamp 1698175906
transform 1 0 67872 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_597
timestamp 1698175906
transform 1 0 68208 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_601
timestamp 1698175906
transform 1 0 68656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_603
timestamp 1698175906
transform 1 0 68880 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_645
timestamp 1698175906
transform 1 0 73584 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_653
timestamp 1698175906
transform 1 0 74480 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_657
timestamp 1698175906
transform 1 0 74928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_667
timestamp 1698175906
transform 1 0 76048 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_683
timestamp 1698175906
transform 1 0 77840 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_687
timestamp 1698175906
transform 1 0 78288 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_104
timestamp 1698175906
transform 1 0 12992 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_108
timestamp 1698175906
transform 1 0 13440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_110
timestamp 1698175906
transform 1 0 13664 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_128
timestamp 1698175906
transform 1 0 15680 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_132
timestamp 1698175906
transform 1 0 16128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_150
timestamp 1698175906
transform 1 0 18144 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_154
timestamp 1698175906
transform 1 0 18592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_156
timestamp 1698175906
transform 1 0 18816 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_164
timestamp 1698175906
transform 1 0 19712 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_168
timestamp 1698175906
transform 1 0 20160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_172
timestamp 1698175906
transform 1 0 20608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_174
timestamp 1698175906
transform 1 0 20832 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_177
timestamp 1698175906
transform 1 0 21168 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_185
timestamp 1698175906
transform 1 0 22064 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_191
timestamp 1698175906
transform 1 0 22736 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_195
timestamp 1698175906
transform 1 0 23184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_203
timestamp 1698175906
transform 1 0 24080 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_207
timestamp 1698175906
transform 1 0 24528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698175906
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_219
timestamp 1698175906
transform 1 0 25872 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_223
timestamp 1698175906
transform 1 0 26320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_227
timestamp 1698175906
transform 1 0 26768 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_231
timestamp 1698175906
transform 1 0 27216 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_234
timestamp 1698175906
transform 1 0 27552 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_278
timestamp 1698175906
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_292
timestamp 1698175906
transform 1 0 34048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_296
timestamp 1698175906
transform 1 0 34496 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_304
timestamp 1698175906
transform 1 0 35392 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_306
timestamp 1698175906
transform 1 0 35616 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_309
timestamp 1698175906
transform 1 0 35952 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_333
timestamp 1698175906
transform 1 0 38640 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_352
timestamp 1698175906
transform 1 0 40768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_360
timestamp 1698175906
transform 1 0 41664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_364
timestamp 1698175906
transform 1 0 42112 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_368
timestamp 1698175906
transform 1 0 42560 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_385
timestamp 1698175906
transform 1 0 44464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_393
timestamp 1698175906
transform 1 0 45360 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_397
timestamp 1698175906
transform 1 0 45808 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_399
timestamp 1698175906
transform 1 0 46032 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_406
timestamp 1698175906
transform 1 0 46816 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_414
timestamp 1698175906
transform 1 0 47712 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_418
timestamp 1698175906
transform 1 0 48160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_422
timestamp 1698175906
transform 1 0 48608 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_430
timestamp 1698175906
transform 1 0 49504 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_432
timestamp 1698175906
transform 1 0 49728 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_435
timestamp 1698175906
transform 1 0 50064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_444
timestamp 1698175906
transform 1 0 51072 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_446
timestamp 1698175906
transform 1 0 51296 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_476
timestamp 1698175906
transform 1 0 54656 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_484
timestamp 1698175906
transform 1 0 55552 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_488
timestamp 1698175906
transform 1 0 56000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_492
timestamp 1698175906
transform 1 0 56448 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_526
timestamp 1698175906
transform 1 0 60256 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_528
timestamp 1698175906
transform 1 0 60480 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_562
timestamp 1698175906
transform 1 0 64288 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_578
timestamp 1698175906
transform 1 0 66080 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_596
timestamp 1698175906
transform 1 0 68096 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_604
timestamp 1698175906
transform 1 0 68992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_608
timestamp 1698175906
transform 1 0 69440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_612
timestamp 1698175906
transform 1 0 69888 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_614
timestamp 1698175906
transform 1 0 70112 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_632
timestamp 1698175906
transform 1 0 72128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_10
timestamp 1698175906
transform 1 0 2464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_14
timestamp 1698175906
transform 1 0 2912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_16
timestamp 1698175906
transform 1 0 3136 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_19
timestamp 1698175906
transform 1 0 3472 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_69
timestamp 1698175906
transform 1 0 9072 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_85
timestamp 1698175906
transform 1 0 10864 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_93
timestamp 1698175906
transform 1 0 11760 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_97
timestamp 1698175906
transform 1 0 12208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_103
timestamp 1698175906
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_111
timestamp 1698175906
transform 1 0 13776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_115
timestamp 1698175906
transform 1 0 14224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_135
timestamp 1698175906
transform 1 0 16464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_139
timestamp 1698175906
transform 1 0 16912 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_147
timestamp 1698175906
transform 1 0 17808 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_151
timestamp 1698175906
transform 1 0 18256 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_162
timestamp 1698175906
transform 1 0 19488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_166
timestamp 1698175906
transform 1 0 19936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_187
timestamp 1698175906
transform 1 0 22288 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_191
timestamp 1698175906
transform 1 0 22736 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_202
timestamp 1698175906
transform 1 0 23968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_206
timestamp 1698175906
transform 1 0 24416 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_220
timestamp 1698175906
transform 1 0 25984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_224
timestamp 1698175906
transform 1 0 26432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_228
timestamp 1698175906
transform 1 0 26880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_232
timestamp 1698175906
transform 1 0 27328 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_236
timestamp 1698175906
transform 1 0 27776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_238
timestamp 1698175906
transform 1 0 28000 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_261
timestamp 1698175906
transform 1 0 30576 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_296
timestamp 1698175906
transform 1 0 34496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_300
timestamp 1698175906
transform 1 0 34944 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_304
timestamp 1698175906
transform 1 0 35392 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_306
timestamp 1698175906
transform 1 0 35616 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_358
timestamp 1698175906
transform 1 0 41440 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_366
timestamp 1698175906
transform 1 0 42336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_374
timestamp 1698175906
transform 1 0 43232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_378
timestamp 1698175906
transform 1 0 43680 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_382
timestamp 1698175906
transform 1 0 44128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_384
timestamp 1698175906
transform 1 0 44352 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_395
timestamp 1698175906
transform 1 0 45584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_399
timestamp 1698175906
transform 1 0 46032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_403
timestamp 1698175906
transform 1 0 46480 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_419
timestamp 1698175906
transform 1 0 48272 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_429
timestamp 1698175906
transform 1 0 49392 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_445
timestamp 1698175906
transform 1 0 51184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_447
timestamp 1698175906
transform 1 0 51408 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_453
timestamp 1698175906
transform 1 0 52080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_457
timestamp 1698175906
transform 1 0 52528 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_493
timestamp 1698175906
transform 1 0 56560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_495
timestamp 1698175906
transform 1 0 56784 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_511
timestamp 1698175906
transform 1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_527
timestamp 1698175906
transform 1 0 60368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_557
timestamp 1698175906
transform 1 0 63728 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_573
timestamp 1698175906
transform 1 0 65520 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_594
timestamp 1698175906
transform 1 0 67872 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_597
timestamp 1698175906
transform 1 0 68208 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_605
timestamp 1698175906
transform 1 0 69104 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_609
timestamp 1698175906
transform 1 0 69552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_611
timestamp 1698175906
transform 1 0 69776 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_641
timestamp 1698175906
transform 1 0 73136 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_657
timestamp 1698175906
transform 1 0 74928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_659
timestamp 1698175906
transform 1 0 75152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_662
timestamp 1698175906
transform 1 0 75488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_664
timestamp 1698175906
transform 1 0 75712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_667
timestamp 1698175906
transform 1 0 76048 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_671
timestamp 1698175906
transform 1 0 76496 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_687
timestamp 1698175906
transform 1 0 78288 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_28
timestamp 1698175906
transform 1 0 4480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_32
timestamp 1698175906
transform 1 0 4928 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_64
timestamp 1698175906
transform 1 0 8512 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_68
timestamp 1698175906
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_80
timestamp 1698175906
transform 1 0 10304 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_133
timestamp 1698175906
transform 1 0 16240 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_137
timestamp 1698175906
transform 1 0 16688 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_155
timestamp 1698175906
transform 1 0 18704 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_159
timestamp 1698175906
transform 1 0 19152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_161
timestamp 1698175906
transform 1 0 19376 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_164
timestamp 1698175906
transform 1 0 19712 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_168
timestamp 1698175906
transform 1 0 20160 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_173
timestamp 1698175906
transform 1 0 20720 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_181
timestamp 1698175906
transform 1 0 21616 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698175906
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_216
timestamp 1698175906
transform 1 0 25536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_220
timestamp 1698175906
transform 1 0 25984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_224
timestamp 1698175906
transform 1 0 26432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_228
timestamp 1698175906
transform 1 0 26880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_232
timestamp 1698175906
transform 1 0 27328 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_365
timestamp 1698175906
transform 1 0 42224 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_373
timestamp 1698175906
transform 1 0 43120 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_375
timestamp 1698175906
transform 1 0 43344 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_378
timestamp 1698175906
transform 1 0 43680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_380
timestamp 1698175906
transform 1 0 43904 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_434
timestamp 1698175906
transform 1 0 49952 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_442
timestamp 1698175906
transform 1 0 50848 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_487
timestamp 1698175906
transform 1 0 55888 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_489
timestamp 1698175906
transform 1 0 56112 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_518
timestamp 1698175906
transform 1 0 59360 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_522
timestamp 1698175906
transform 1 0 59808 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_562
timestamp 1698175906
transform 1 0 64288 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_566
timestamp 1698175906
transform 1 0 64736 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_602
timestamp 1698175906
transform 1 0 68768 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_606
timestamp 1698175906
transform 1 0 69216 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_632
timestamp 1698175906
transform 1 0 72128 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_11
timestamp 1698175906
transform 1 0 2576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_17
timestamp 1698175906
transform 1 0 3248 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_21
timestamp 1698175906
transform 1 0 3696 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_25
timestamp 1698175906
transform 1 0 4144 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_28
timestamp 1698175906
transform 1 0 4480 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698175906
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_111
timestamp 1698175906
transform 1 0 13776 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_117
timestamp 1698175906
transform 1 0 14448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_121
timestamp 1698175906
transform 1 0 14896 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_155
timestamp 1698175906
transform 1 0 18704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_159
timestamp 1698175906
transform 1 0 19152 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_209
timestamp 1698175906
transform 1 0 24752 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_217
timestamp 1698175906
transform 1 0 25648 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_235
timestamp 1698175906
transform 1 0 27664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_249
timestamp 1698175906
transform 1 0 29232 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_303
timestamp 1698175906
transform 1 0 35280 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_305
timestamp 1698175906
transform 1 0 35504 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_319
timestamp 1698175906
transform 1 0 37072 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_328
timestamp 1698175906
transform 1 0 38080 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_353
timestamp 1698175906
transform 1 0 40880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_357
timestamp 1698175906
transform 1 0 41328 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_365
timestamp 1698175906
transform 1 0 42224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_367
timestamp 1698175906
transform 1 0 42448 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_370
timestamp 1698175906
transform 1 0 42784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_374
timestamp 1698175906
transform 1 0 43232 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_387
timestamp 1698175906
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_391
timestamp 1698175906
transform 1 0 45136 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_403
timestamp 1698175906
transform 1 0 46480 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_405
timestamp 1698175906
transform 1 0 46704 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_424
timestamp 1698175906
transform 1 0 48832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_457
timestamp 1698175906
transform 1 0 52528 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_465
timestamp 1698175906
transform 1 0 53424 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_467
timestamp 1698175906
transform 1 0 53648 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_507
timestamp 1698175906
transform 1 0 58128 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_523
timestamp 1698175906
transform 1 0 59920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_558
timestamp 1698175906
transform 1 0 63840 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_562
timestamp 1698175906
transform 1 0 64288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_564
timestamp 1698175906
transform 1 0 64512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_594
timestamp 1698175906
transform 1 0 67872 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_597
timestamp 1698175906
transform 1 0 68208 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_601
timestamp 1698175906
transform 1 0 68656 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_609
timestamp 1698175906
transform 1 0 69552 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_642
timestamp 1698175906
transform 1 0 73248 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_648
timestamp 1698175906
transform 1 0 73920 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_656
timestamp 1698175906
transform 1 0 74816 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_662
timestamp 1698175906
transform 1 0 75488 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_664
timestamp 1698175906
transform 1 0 75712 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_667
timestamp 1698175906
transform 1 0 76048 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_671
timestamp 1698175906
transform 1 0 76496 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_687
timestamp 1698175906
transform 1 0 78288 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_36
timestamp 1698175906
transform 1 0 5376 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_68
timestamp 1698175906
transform 1 0 8960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_76
timestamp 1698175906
transform 1 0 9856 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_149
timestamp 1698175906
transform 1 0 18032 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_153
timestamp 1698175906
transform 1 0 18480 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_190
timestamp 1698175906
transform 1 0 22624 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_200
timestamp 1698175906
transform 1 0 23744 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_254
timestamp 1698175906
transform 1 0 29792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_270
timestamp 1698175906
transform 1 0 31584 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698175906
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_292
timestamp 1698175906
transform 1 0 34048 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_300
timestamp 1698175906
transform 1 0 34944 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_302
timestamp 1698175906
transform 1 0 35168 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_305
timestamp 1698175906
transform 1 0 35504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_322
timestamp 1698175906
transform 1 0 37408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_340
timestamp 1698175906
transform 1 0 39424 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_342
timestamp 1698175906
transform 1 0 39648 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_347
timestamp 1698175906
transform 1 0 40208 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698175906
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_352
timestamp 1698175906
transform 1 0 40768 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_360
timestamp 1698175906
transform 1 0 41664 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_405
timestamp 1698175906
transform 1 0 46704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_409
timestamp 1698175906
transform 1 0 47152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_411
timestamp 1698175906
transform 1 0 47376 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_432
timestamp 1698175906
transform 1 0 49728 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_436
timestamp 1698175906
transform 1 0 50176 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_480
timestamp 1698175906
transform 1 0 55104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_484
timestamp 1698175906
transform 1 0 55552 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_488
timestamp 1698175906
transform 1 0 56000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_492
timestamp 1698175906
transform 1 0 56448 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_500
timestamp 1698175906
transform 1 0 57344 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_535
timestamp 1698175906
transform 1 0 61264 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_551
timestamp 1698175906
transform 1 0 63056 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_555
timestamp 1698175906
transform 1 0 63504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_557
timestamp 1698175906
transform 1 0 63728 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_594
timestamp 1698175906
transform 1 0 67872 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_596
timestamp 1698175906
transform 1 0 68096 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_629
timestamp 1698175906
transform 1 0 71792 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_632
timestamp 1698175906
transform 1 0 72128 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_28
timestamp 1698175906
transform 1 0 4480 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_32
timestamp 1698175906
transform 1 0 4928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_36
timestamp 1698175906
transform 1 0 5376 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_44
timestamp 1698175906
transform 1 0 6272 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_55
timestamp 1698175906
transform 1 0 7504 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_63
timestamp 1698175906
transform 1 0 8400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_65
timestamp 1698175906
transform 1 0 8624 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_78
timestamp 1698175906
transform 1 0 10080 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_86
timestamp 1698175906
transform 1 0 10976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_88
timestamp 1698175906
transform 1 0 11200 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_99
timestamp 1698175906
transform 1 0 12432 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_104
timestamp 1698175906
transform 1 0 12992 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_108
timestamp 1698175906
transform 1 0 13440 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_110
timestamp 1698175906
transform 1 0 13664 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_119
timestamp 1698175906
transform 1 0 14672 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_127
timestamp 1698175906
transform 1 0 15568 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_131
timestamp 1698175906
transform 1 0 16016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_133
timestamp 1698175906
transform 1 0 16240 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_144
timestamp 1698175906
transform 1 0 17472 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_148
timestamp 1698175906
transform 1 0 17920 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_152
timestamp 1698175906
transform 1 0 18368 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_154
timestamp 1698175906
transform 1 0 18592 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_165
timestamp 1698175906
transform 1 0 19824 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_169
timestamp 1698175906
transform 1 0 20272 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_172
timestamp 1698175906
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_176
timestamp 1698175906
transform 1 0 21056 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_187
timestamp 1698175906
transform 1 0 22288 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_195
timestamp 1698175906
transform 1 0 23184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_197
timestamp 1698175906
transform 1 0 23408 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_200
timestamp 1698175906
transform 1 0 23744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_214
timestamp 1698175906
transform 1 0 25312 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_218
timestamp 1698175906
transform 1 0 25760 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_221
timestamp 1698175906
transform 1 0 26096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_237
timestamp 1698175906
transform 1 0 27888 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_240
timestamp 1698175906
transform 1 0 28224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_242
timestamp 1698175906
transform 1 0 28448 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_251
timestamp 1698175906
transform 1 0 29456 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_255
timestamp 1698175906
transform 1 0 29904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_257
timestamp 1698175906
transform 1 0 30128 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_264
timestamp 1698175906
transform 1 0 30912 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_268
timestamp 1698175906
transform 1 0 31360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_286
timestamp 1698175906
transform 1 0 33376 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_288
timestamp 1698175906
transform 1 0 33600 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_297
timestamp 1698175906
transform 1 0 34608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_301
timestamp 1698175906
transform 1 0 35056 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_303
timestamp 1698175906
transform 1 0 35280 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_308
timestamp 1698175906
transform 1 0 35840 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_310
timestamp 1698175906
transform 1 0 36064 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_325
timestamp 1698175906
transform 1 0 37744 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_329
timestamp 1698175906
transform 1 0 38192 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_342
timestamp 1698175906
transform 1 0 39648 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_346
timestamp 1698175906
transform 1 0 40096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_376
timestamp 1698175906
transform 1 0 43456 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_403
timestamp 1698175906
transform 1 0 46480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_407
timestamp 1698175906
transform 1 0 46928 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_436
timestamp 1698175906
transform 1 0 50176 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_440
timestamp 1698175906
transform 1 0 50624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_470
timestamp 1698175906
transform 1 0 53984 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_474
timestamp 1698175906
transform 1 0 54432 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_504
timestamp 1698175906
transform 1 0 57792 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_508
timestamp 1698175906
transform 1 0 58240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_538
timestamp 1698175906
transform 1 0 61600 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_542
timestamp 1698175906
transform 1 0 62048 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_572
timestamp 1698175906
transform 1 0 65408 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_606
timestamp 1698175906
transform 1 0 69216 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_610
timestamp 1698175906
transform 1 0 69664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_614
timestamp 1698175906
transform 1 0 70112 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_616
timestamp 1698175906
transform 1 0 70336 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_645
timestamp 1698175906
transform 1 0 73584 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_674
timestamp 1698175906
transform 1 0 76832 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_678
timestamp 1698175906
transform 1 0 77280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_682
timestamp 1698175906
transform 1 0 77728 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_686
timestamp 1698175906
transform 1 0 78176 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698175906
transform -1 0 72912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698175906
transform 1 0 4480 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698175906
transform 1 0 44016 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698175906
transform 1 0 48048 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698175906
transform 1 0 52080 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698175906
transform 1 0 56112 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698175906
transform 1 0 60144 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input8
timestamp 1698175906
transform 1 0 64176 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698175906
transform 1 0 7728 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698175906
transform 1 0 11760 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698175906
transform 1 0 15792 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698175906
transform -1 0 21280 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698175906
transform -1 0 25088 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698175906
transform 1 0 35952 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698175906
transform 1 0 39984 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input18
timestamp 1698175906
transform 1 0 38528 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input19
timestamp 1698175906
transform 1 0 14000 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input20
timestamp 1698175906
transform 1 0 11536 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input21
timestamp 1698175906
transform 1 0 9184 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input22
timestamp 1698175906
transform 1 0 6608 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input23
timestamp 1698175906
transform 1 0 4480 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input24
timestamp 1698175906
transform 1 0 1680 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input25
timestamp 1698175906
transform -1 0 36848 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input26
timestamp 1698175906
transform 1 0 33712 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input27
timestamp 1698175906
transform 1 0 32704 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input28
timestamp 1698175906
transform -1 0 29456 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698175906
transform 1 0 27216 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input30
timestamp 1698175906
transform 1 0 24416 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input31
timestamp 1698175906
transform 1 0 21392 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input32
timestamp 1698175906
transform 1 0 18928 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input33
timestamp 1698175906
transform 1 0 16800 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input34
timestamp 1698175906
transform 1 0 76272 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output35 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4480 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output36
timestamp 1698175906
transform -1 0 4480 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output37
timestamp 1698175906
transform -1 0 4480 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output38
timestamp 1698175906
transform -1 0 4480 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output39
timestamp 1698175906
transform -1 0 4480 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output40
timestamp 1698175906
transform -1 0 4480 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output41
timestamp 1698175906
transform -1 0 4480 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output42
timestamp 1698175906
transform -1 0 4480 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output43
timestamp 1698175906
transform -1 0 4480 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output44
timestamp 1698175906
transform -1 0 4480 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output45
timestamp 1698175906
transform -1 0 4480 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output46
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output47
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output48
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output49
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output50
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output51
timestamp 1698175906
transform -1 0 77504 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output52
timestamp 1698175906
transform 1 0 75488 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output53
timestamp 1698175906
transform 1 0 72912 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output54
timestamp 1698175906
transform 1 0 75488 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output55
timestamp 1698175906
transform 1 0 75488 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output56
timestamp 1698175906
transform 1 0 72576 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output57
timestamp 1698175906
transform 1 0 72576 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output58
timestamp 1698175906
transform 1 0 75488 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output59
timestamp 1698175906
transform 1 0 75488 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output60
timestamp 1698175906
transform 1 0 75488 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output61
timestamp 1698175906
transform -1 0 75824 0 1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output62
timestamp 1698175906
transform -1 0 75824 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output63
timestamp 1698175906
transform 1 0 75488 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output64
timestamp 1698175906
transform 1 0 72576 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output65
timestamp 1698175906
transform 1 0 75488 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output66
timestamp 1698175906
transform 1 0 72912 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output67
timestamp 1698175906
transform 1 0 68320 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output68
timestamp 1698175906
transform 1 0 72576 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output69
timestamp 1698175906
transform 1 0 54880 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output70
timestamp 1698175906
transform -1 0 53872 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output71
timestamp 1698175906
transform -1 0 53984 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output72
timestamp 1698175906
transform -1 0 50176 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output73
timestamp 1698175906
transform -1 0 46480 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output74
timestamp 1698175906
transform -1 0 43232 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output75
timestamp 1698175906
transform 1 0 75488 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output76
timestamp 1698175906
transform 1 0 73920 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output77
timestamp 1698175906
transform 1 0 70672 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output78
timestamp 1698175906
transform 1 0 68208 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output79
timestamp 1698175906
transform 1 0 66304 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output80
timestamp 1698175906
transform 1 0 64288 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output81
timestamp 1698175906
transform 1 0 60816 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output82
timestamp 1698175906
transform 1 0 62496 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output83
timestamp 1698175906
transform 1 0 58688 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_43 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_44
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_45
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_86 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_87
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_88
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_89
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_100
timestamp 1698175906
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_101
timestamp 1698175906
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_102
timestamp 1698175906
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_103
timestamp 1698175906
transform 1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_104
timestamp 1698175906
transform 1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698175906
transform 1 0 77504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_106
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_107
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_108
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_109
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_110
timestamp 1698175906
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_111
timestamp 1698175906
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_112
timestamp 1698175906
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_113
timestamp 1698175906
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_114
timestamp 1698175906
transform 1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_115
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_116
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_117
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_118
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_119
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_120
timestamp 1698175906
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_121
timestamp 1698175906
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_122
timestamp 1698175906
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_123
timestamp 1698175906
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_124
timestamp 1698175906
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_125
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_126
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_127
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_128
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_129
timestamp 1698175906
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_130
timestamp 1698175906
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_131
timestamp 1698175906
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_132
timestamp 1698175906
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_133
timestamp 1698175906
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_134
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_135
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_136
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_137
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_138
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_139
timestamp 1698175906
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_140
timestamp 1698175906
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_141
timestamp 1698175906
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_142
timestamp 1698175906
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_143
timestamp 1698175906
transform 1 0 75824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_144
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_145
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_146
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_147
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_148
timestamp 1698175906
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_149
timestamp 1698175906
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_150
timestamp 1698175906
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_151
timestamp 1698175906
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_152
timestamp 1698175906
transform 1 0 71904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_153
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_154
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_155
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_156
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_157
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_158
timestamp 1698175906
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_159
timestamp 1698175906
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_160
timestamp 1698175906
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_161
timestamp 1698175906
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_162
timestamp 1698175906
transform 1 0 75824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_163
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_164
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_165
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_166
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_167
timestamp 1698175906
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_168
timestamp 1698175906
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_169
timestamp 1698175906
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_170
timestamp 1698175906
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_171
timestamp 1698175906
transform 1 0 71904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_172
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_173
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_174
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_175
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_176
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_177
timestamp 1698175906
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_178
timestamp 1698175906
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_179
timestamp 1698175906
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_180
timestamp 1698175906
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_181
timestamp 1698175906
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_182
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_183
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_184
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_185
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_186
timestamp 1698175906
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_187
timestamp 1698175906
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_188
timestamp 1698175906
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_189
timestamp 1698175906
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_190
timestamp 1698175906
transform 1 0 71904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_191
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_192
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_193
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_194
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_195
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_196
timestamp 1698175906
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_197
timestamp 1698175906
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_198
timestamp 1698175906
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_199
timestamp 1698175906
transform 1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_200
timestamp 1698175906
transform 1 0 75824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_201
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_202
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_203
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_204
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_205
timestamp 1698175906
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_206
timestamp 1698175906
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_207
timestamp 1698175906
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_208
timestamp 1698175906
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_209
timestamp 1698175906
transform 1 0 71904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_210
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_211
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_212
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_213
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_214
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_215
timestamp 1698175906
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_216
timestamp 1698175906
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_217
timestamp 1698175906
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_218
timestamp 1698175906
transform 1 0 67984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_219
timestamp 1698175906
transform 1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_220
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_221
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_222
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_223
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_224
timestamp 1698175906
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_225
timestamp 1698175906
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_226
timestamp 1698175906
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_227
timestamp 1698175906
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_228
timestamp 1698175906
transform 1 0 71904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_229
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_230
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_231
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_232
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_233
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_234
timestamp 1698175906
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_235
timestamp 1698175906
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_236
timestamp 1698175906
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_237
timestamp 1698175906
transform 1 0 67984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_238
timestamp 1698175906
transform 1 0 75824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_239
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_240
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_241
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_242
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_243
timestamp 1698175906
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_244
timestamp 1698175906
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_245
timestamp 1698175906
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_246
timestamp 1698175906
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_247
timestamp 1698175906
transform 1 0 71904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_248
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_249
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_250
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_251
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_252
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_253
timestamp 1698175906
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_254
timestamp 1698175906
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698175906
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698175906
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698175906
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_258
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_259
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_260
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_261
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698175906
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698175906
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698175906
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698175906
transform 1 0 64064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698175906
transform 1 0 71904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_267
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_268
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698175906
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698175906
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698175906
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698175906
transform 1 0 67984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_276
timestamp 1698175906
transform 1 0 75824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698175906
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698175906
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_283
timestamp 1698175906
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_284
timestamp 1698175906
transform 1 0 64064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_285
timestamp 1698175906
transform 1 0 71904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_290
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_291
timestamp 1698175906
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_292
timestamp 1698175906
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_293
timestamp 1698175906
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_294
timestamp 1698175906
transform 1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_295
timestamp 1698175906
transform 1 0 75824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_297
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_298
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_299
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_300
timestamp 1698175906
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_301
timestamp 1698175906
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_302
timestamp 1698175906
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_303
timestamp 1698175906
transform 1 0 64064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_304
timestamp 1698175906
transform 1 0 71904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_305
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_306
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_307
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_308
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_309
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_310
timestamp 1698175906
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_311
timestamp 1698175906
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_312
timestamp 1698175906
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_313
timestamp 1698175906
transform 1 0 67984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_314
timestamp 1698175906
transform 1 0 75824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_315
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_316
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_317
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_318
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_319
timestamp 1698175906
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_320
timestamp 1698175906
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_321
timestamp 1698175906
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_322
timestamp 1698175906
transform 1 0 64064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_323
timestamp 1698175906
transform 1 0 71904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_324
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_325
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_326
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_327
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_328
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_329
timestamp 1698175906
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_330
timestamp 1698175906
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_331
timestamp 1698175906
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_332
timestamp 1698175906
transform 1 0 67984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_333
timestamp 1698175906
transform 1 0 75824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_334
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_335
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_336
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_337
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_338
timestamp 1698175906
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_339
timestamp 1698175906
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_340
timestamp 1698175906
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_341
timestamp 1698175906
transform 1 0 64064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_342
timestamp 1698175906
transform 1 0 71904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_343
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_344
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_345
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_346
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_347
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_348
timestamp 1698175906
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_349
timestamp 1698175906
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_350
timestamp 1698175906
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_351
timestamp 1698175906
transform 1 0 67984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_352
timestamp 1698175906
transform 1 0 75824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_353
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_354
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_355
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_356
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_357
timestamp 1698175906
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_358
timestamp 1698175906
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_359
timestamp 1698175906
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_360
timestamp 1698175906
transform 1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_361
timestamp 1698175906
transform 1 0 71904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_362
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_363
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_364
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_365
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_366
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_367
timestamp 1698175906
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_368
timestamp 1698175906
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_369
timestamp 1698175906
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_370
timestamp 1698175906
transform 1 0 67984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_371
timestamp 1698175906
transform 1 0 75824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_372
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_373
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_374
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_375
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_376
timestamp 1698175906
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_377
timestamp 1698175906
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_378
timestamp 1698175906
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_379
timestamp 1698175906
transform 1 0 64064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_380
timestamp 1698175906
transform 1 0 71904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_381
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_382
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_383
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_384
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_385
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_386
timestamp 1698175906
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_387
timestamp 1698175906
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_388
timestamp 1698175906
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_389
timestamp 1698175906
transform 1 0 67984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_390
timestamp 1698175906
transform 1 0 75824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_391
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_392
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_393
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_394
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_395
timestamp 1698175906
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_396
timestamp 1698175906
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_397
timestamp 1698175906
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_398
timestamp 1698175906
transform 1 0 64064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_399
timestamp 1698175906
transform 1 0 71904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_400
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_401
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_402
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_403
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_404
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_405
timestamp 1698175906
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_406
timestamp 1698175906
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_407
timestamp 1698175906
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_408
timestamp 1698175906
transform 1 0 67984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_409
timestamp 1698175906
transform 1 0 75824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_410
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_411
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_412
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_413
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_414
timestamp 1698175906
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_415
timestamp 1698175906
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_416
timestamp 1698175906
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_417
timestamp 1698175906
transform 1 0 64064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_418
timestamp 1698175906
transform 1 0 71904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_419
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_420
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_421
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_422
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_423
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_424
timestamp 1698175906
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_425
timestamp 1698175906
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_426
timestamp 1698175906
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_427
timestamp 1698175906
transform 1 0 67984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_428
timestamp 1698175906
transform 1 0 75824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_429
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_430
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_431
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_432
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_433
timestamp 1698175906
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_434
timestamp 1698175906
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_435
timestamp 1698175906
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_436
timestamp 1698175906
transform 1 0 64064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_437
timestamp 1698175906
transform 1 0 71904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_438
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_439
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_440
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_441
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_442
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_443
timestamp 1698175906
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_444
timestamp 1698175906
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_445
timestamp 1698175906
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_446
timestamp 1698175906
transform 1 0 67984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_447
timestamp 1698175906
transform 1 0 75824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_448
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_449
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_450
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_451
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_452
timestamp 1698175906
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_453
timestamp 1698175906
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_454
timestamp 1698175906
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_455
timestamp 1698175906
transform 1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_456
timestamp 1698175906
transform 1 0 71904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_457
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_458
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_459
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_460
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_461
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_462
timestamp 1698175906
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_463
timestamp 1698175906
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_464
timestamp 1698175906
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_465
timestamp 1698175906
transform 1 0 67984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_466
timestamp 1698175906
transform 1 0 75824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_467
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_468
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_469
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_470
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_471
timestamp 1698175906
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_472
timestamp 1698175906
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_473
timestamp 1698175906
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_474
timestamp 1698175906
transform 1 0 64064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_475
timestamp 1698175906
transform 1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_476
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_477
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_478
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_479
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_480
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_481
timestamp 1698175906
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_482
timestamp 1698175906
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_483
timestamp 1698175906
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_484
timestamp 1698175906
transform 1 0 67984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_485
timestamp 1698175906
transform 1 0 75824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_486
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_487
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_488
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_489
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_490
timestamp 1698175906
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_491
timestamp 1698175906
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_492
timestamp 1698175906
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_493
timestamp 1698175906
transform 1 0 64064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_494
timestamp 1698175906
transform 1 0 71904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_495
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_496
timestamp 1698175906
transform 1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_497
timestamp 1698175906
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_498
timestamp 1698175906
transform 1 0 16576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_499
timestamp 1698175906
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_500
timestamp 1698175906
transform 1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_501
timestamp 1698175906
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_502
timestamp 1698175906
transform 1 0 31808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_503
timestamp 1698175906
transform 1 0 35616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_504
timestamp 1698175906
transform 1 0 39424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_505
timestamp 1698175906
transform 1 0 43232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_506
timestamp 1698175906
transform 1 0 47040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_507
timestamp 1698175906
transform 1 0 50848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_508
timestamp 1698175906
transform 1 0 54656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_509
timestamp 1698175906
transform 1 0 58464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_510
timestamp 1698175906
transform 1 0 62272 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_511
timestamp 1698175906
transform 1 0 66080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_512
timestamp 1698175906
transform 1 0 69888 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_513
timestamp 1698175906
transform 1 0 73696 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_514
timestamp 1698175906
transform 1 0 77504 0 1 36064
box -86 -86 310 870
<< labels >>
flabel metal2 s 72128 0 72240 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 38304 800 38416 0 FreeSans 448 0 0 0 dmem_addr[0]
port 1 nsew signal tristate
flabel metal3 s 0 13664 800 13776 0 FreeSans 448 0 0 0 dmem_addr[10]
port 2 nsew signal tristate
flabel metal3 s 0 11200 800 11312 0 FreeSans 448 0 0 0 dmem_addr[11]
port 3 nsew signal tristate
flabel metal3 s 0 8736 800 8848 0 FreeSans 448 0 0 0 dmem_addr[12]
port 4 nsew signal tristate
flabel metal3 s 0 6272 800 6384 0 FreeSans 448 0 0 0 dmem_addr[13]
port 5 nsew signal tristate
flabel metal3 s 0 3808 800 3920 0 FreeSans 448 0 0 0 dmem_addr[14]
port 6 nsew signal tristate
flabel metal3 s 0 1344 800 1456 0 FreeSans 448 0 0 0 dmem_addr[15]
port 7 nsew signal tristate
flabel metal3 s 0 35840 800 35952 0 FreeSans 448 0 0 0 dmem_addr[1]
port 8 nsew signal tristate
flabel metal3 s 0 33376 800 33488 0 FreeSans 448 0 0 0 dmem_addr[2]
port 9 nsew signal tristate
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 dmem_addr[3]
port 10 nsew signal tristate
flabel metal3 s 0 28448 800 28560 0 FreeSans 448 0 0 0 dmem_addr[4]
port 11 nsew signal tristate
flabel metal3 s 0 25984 800 26096 0 FreeSans 448 0 0 0 dmem_addr[5]
port 12 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 dmem_addr[6]
port 13 nsew signal tristate
flabel metal3 s 0 21056 800 21168 0 FreeSans 448 0 0 0 dmem_addr[7]
port 14 nsew signal tristate
flabel metal3 s 0 18592 800 18704 0 FreeSans 448 0 0 0 dmem_addr[8]
port 15 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 dmem_addr[9]
port 16 nsew signal tristate
flabel metal3 s 79200 1344 80000 1456 0 FreeSans 448 0 0 0 dmem_data_in[0]
port 17 nsew signal tristate
flabel metal3 s 79200 25984 80000 26096 0 FreeSans 448 0 0 0 dmem_data_in[10]
port 18 nsew signal tristate
flabel metal3 s 79200 28448 80000 28560 0 FreeSans 448 0 0 0 dmem_data_in[11]
port 19 nsew signal tristate
flabel metal3 s 79200 30912 80000 31024 0 FreeSans 448 0 0 0 dmem_data_in[12]
port 20 nsew signal tristate
flabel metal3 s 79200 33376 80000 33488 0 FreeSans 448 0 0 0 dmem_data_in[13]
port 21 nsew signal tristate
flabel metal3 s 79200 35840 80000 35952 0 FreeSans 448 0 0 0 dmem_data_in[14]
port 22 nsew signal tristate
flabel metal3 s 79200 38304 80000 38416 0 FreeSans 448 0 0 0 dmem_data_in[15]
port 23 nsew signal tristate
flabel metal3 s 79200 3808 80000 3920 0 FreeSans 448 0 0 0 dmem_data_in[1]
port 24 nsew signal tristate
flabel metal3 s 79200 6272 80000 6384 0 FreeSans 448 0 0 0 dmem_data_in[2]
port 25 nsew signal tristate
flabel metal3 s 79200 8736 80000 8848 0 FreeSans 448 0 0 0 dmem_data_in[3]
port 26 nsew signal tristate
flabel metal3 s 79200 11200 80000 11312 0 FreeSans 448 0 0 0 dmem_data_in[4]
port 27 nsew signal tristate
flabel metal3 s 79200 13664 80000 13776 0 FreeSans 448 0 0 0 dmem_data_in[5]
port 28 nsew signal tristate
flabel metal3 s 79200 16128 80000 16240 0 FreeSans 448 0 0 0 dmem_data_in[6]
port 29 nsew signal tristate
flabel metal3 s 79200 18592 80000 18704 0 FreeSans 448 0 0 0 dmem_data_in[7]
port 30 nsew signal tristate
flabel metal3 s 79200 21056 80000 21168 0 FreeSans 448 0 0 0 dmem_data_in[8]
port 31 nsew signal tristate
flabel metal3 s 79200 23520 80000 23632 0 FreeSans 448 0 0 0 dmem_data_in[9]
port 32 nsew signal tristate
flabel metal2 s 3584 0 3696 800 0 FreeSans 448 90 0 0 dmem_data_out[0]
port 33 nsew signal input
flabel metal2 s 43904 0 44016 800 0 FreeSans 448 90 0 0 dmem_data_out[10]
port 34 nsew signal input
flabel metal2 s 47936 0 48048 800 0 FreeSans 448 90 0 0 dmem_data_out[11]
port 35 nsew signal input
flabel metal2 s 51968 0 52080 800 0 FreeSans 448 90 0 0 dmem_data_out[12]
port 36 nsew signal input
flabel metal2 s 56000 0 56112 800 0 FreeSans 448 90 0 0 dmem_data_out[13]
port 37 nsew signal input
flabel metal2 s 60032 0 60144 800 0 FreeSans 448 90 0 0 dmem_data_out[14]
port 38 nsew signal input
flabel metal2 s 64064 0 64176 800 0 FreeSans 448 90 0 0 dmem_data_out[15]
port 39 nsew signal input
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 dmem_data_out[1]
port 40 nsew signal input
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 dmem_data_out[2]
port 41 nsew signal input
flabel metal2 s 15680 0 15792 800 0 FreeSans 448 90 0 0 dmem_data_out[3]
port 42 nsew signal input
flabel metal2 s 19712 0 19824 800 0 FreeSans 448 90 0 0 dmem_data_out[4]
port 43 nsew signal input
flabel metal2 s 23744 0 23856 800 0 FreeSans 448 90 0 0 dmem_data_out[5]
port 44 nsew signal input
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 dmem_data_out[6]
port 45 nsew signal input
flabel metal2 s 31808 0 31920 800 0 FreeSans 448 90 0 0 dmem_data_out[7]
port 46 nsew signal input
flabel metal2 s 35840 0 35952 800 0 FreeSans 448 90 0 0 dmem_data_out[8]
port 47 nsew signal input
flabel metal2 s 39872 0 39984 800 0 FreeSans 448 90 0 0 dmem_data_out[9]
port 48 nsew signal input
flabel metal2 s 68096 0 68208 800 0 FreeSans 448 90 0 0 dmem_we
port 49 nsew signal tristate
flabel metal2 s 38528 39200 38640 40000 0 FreeSans 448 90 0 0 instr[0]
port 50 nsew signal input
flabel metal2 s 13888 39200 14000 40000 0 FreeSans 448 90 0 0 instr[10]
port 51 nsew signal input
flabel metal2 s 11424 39200 11536 40000 0 FreeSans 448 90 0 0 instr[11]
port 52 nsew signal input
flabel metal2 s 8960 39200 9072 40000 0 FreeSans 448 90 0 0 instr[12]
port 53 nsew signal input
flabel metal2 s 6496 39200 6608 40000 0 FreeSans 448 90 0 0 instr[13]
port 54 nsew signal input
flabel metal2 s 4032 39200 4144 40000 0 FreeSans 448 90 0 0 instr[14]
port 55 nsew signal input
flabel metal2 s 1568 39200 1680 40000 0 FreeSans 448 90 0 0 instr[15]
port 56 nsew signal input
flabel metal2 s 36064 39200 36176 40000 0 FreeSans 448 90 0 0 instr[1]
port 57 nsew signal input
flabel metal2 s 33600 39200 33712 40000 0 FreeSans 448 90 0 0 instr[2]
port 58 nsew signal input
flabel metal2 s 31136 39200 31248 40000 0 FreeSans 448 90 0 0 instr[3]
port 59 nsew signal input
flabel metal2 s 28672 39200 28784 40000 0 FreeSans 448 90 0 0 instr[4]
port 60 nsew signal input
flabel metal2 s 26208 39200 26320 40000 0 FreeSans 448 90 0 0 instr[5]
port 61 nsew signal input
flabel metal2 s 23744 39200 23856 40000 0 FreeSans 448 90 0 0 instr[6]
port 62 nsew signal input
flabel metal2 s 21280 39200 21392 40000 0 FreeSans 448 90 0 0 instr[7]
port 63 nsew signal input
flabel metal2 s 18816 39200 18928 40000 0 FreeSans 448 90 0 0 instr[8]
port 64 nsew signal input
flabel metal2 s 16352 39200 16464 40000 0 FreeSans 448 90 0 0 instr[9]
port 65 nsew signal input
flabel metal2 s 77952 39200 78064 40000 0 FreeSans 448 90 0 0 pc[0]
port 66 nsew signal tristate
flabel metal2 s 53312 39200 53424 40000 0 FreeSans 448 90 0 0 pc[10]
port 67 nsew signal tristate
flabel metal2 s 50848 39200 50960 40000 0 FreeSans 448 90 0 0 pc[11]
port 68 nsew signal tristate
flabel metal2 s 48384 39200 48496 40000 0 FreeSans 448 90 0 0 pc[12]
port 69 nsew signal tristate
flabel metal2 s 45920 39200 46032 40000 0 FreeSans 448 90 0 0 pc[13]
port 70 nsew signal tristate
flabel metal2 s 43456 39200 43568 40000 0 FreeSans 448 90 0 0 pc[14]
port 71 nsew signal tristate
flabel metal2 s 40992 39200 41104 40000 0 FreeSans 448 90 0 0 pc[15]
port 72 nsew signal tristate
flabel metal2 s 75488 39200 75600 40000 0 FreeSans 448 90 0 0 pc[1]
port 73 nsew signal tristate
flabel metal2 s 73024 39200 73136 40000 0 FreeSans 448 90 0 0 pc[2]
port 74 nsew signal tristate
flabel metal2 s 70560 39200 70672 40000 0 FreeSans 448 90 0 0 pc[3]
port 75 nsew signal tristate
flabel metal2 s 68096 39200 68208 40000 0 FreeSans 448 90 0 0 pc[4]
port 76 nsew signal tristate
flabel metal2 s 65632 39200 65744 40000 0 FreeSans 448 90 0 0 pc[5]
port 77 nsew signal tristate
flabel metal2 s 63168 39200 63280 40000 0 FreeSans 448 90 0 0 pc[6]
port 78 nsew signal tristate
flabel metal2 s 60704 39200 60816 40000 0 FreeSans 448 90 0 0 pc[7]
port 79 nsew signal tristate
flabel metal2 s 58240 39200 58352 40000 0 FreeSans 448 90 0 0 pc[8]
port 80 nsew signal tristate
flabel metal2 s 55776 39200 55888 40000 0 FreeSans 448 90 0 0 pc[9]
port 81 nsew signal tristate
flabel metal2 s 76160 0 76272 800 0 FreeSans 448 90 0 0 rst_n
port 82 nsew signal input
flabel metal4 s 10844 3076 11164 36908 0 FreeSans 1280 90 0 0 vdd
port 83 nsew power bidirectional
flabel metal4 s 30164 3076 30484 36908 0 FreeSans 1280 90 0 0 vdd
port 83 nsew power bidirectional
flabel metal4 s 49484 3076 49804 36908 0 FreeSans 1280 90 0 0 vdd
port 83 nsew power bidirectional
flabel metal4 s 68804 3076 69124 36908 0 FreeSans 1280 90 0 0 vdd
port 83 nsew power bidirectional
flabel metal4 s 20504 3076 20824 36908 0 FreeSans 1280 90 0 0 vss
port 84 nsew ground bidirectional
flabel metal4 s 39824 3076 40144 36908 0 FreeSans 1280 90 0 0 vss
port 84 nsew ground bidirectional
flabel metal4 s 59144 3076 59464 36908 0 FreeSans 1280 90 0 0 vss
port 84 nsew ground bidirectional
flabel metal4 s 78464 3076 78784 36908 0 FreeSans 1280 90 0 0 vss
port 84 nsew ground bidirectional
rlabel metal1 39984 36848 39984 36848 0 vdd
rlabel via1 40064 36064 40064 36064 0 vss
rlabel metal2 17080 5600 17080 5600 0 _0000_
rlabel metal2 22232 5600 22232 5600 0 _0001_
rlabel metal2 3304 13216 3304 13216 0 _0002_
rlabel metal2 5656 28560 5656 28560 0 _0003_
rlabel metal2 2520 11872 2520 11872 0 _0004_
rlabel metal2 7952 28728 7952 28728 0 _0005_
rlabel metal2 36568 7784 36568 7784 0 _0006_
rlabel metal2 44408 4648 44408 4648 0 _0007_
rlabel metal2 53368 6944 53368 6944 0 _0008_
rlabel metal2 65800 9184 65800 9184 0 _0009_
rlabel metal2 64176 20664 64176 20664 0 _0010_
rlabel metal2 45192 13048 45192 13048 0 _0011_
rlabel metal2 65352 34552 65352 34552 0 _0012_
rlabel metal3 70560 34328 70560 34328 0 _0013_
rlabel metal3 75656 13832 75656 13832 0 _0014_
rlabel metal2 73472 9576 73472 9576 0 _0015_
rlabel metal2 10808 7896 10808 7896 0 _0016_
rlabel metal2 26936 9352 26936 9352 0 _0017_
rlabel metal2 6888 17192 6888 17192 0 _0018_
rlabel metal2 4648 21056 4648 21056 0 _0019_
rlabel metal2 7784 5376 7784 5376 0 _0020_
rlabel metal2 7784 21056 7784 21056 0 _0021_
rlabel metal2 30520 8344 30520 8344 0 _0022_
rlabel metal2 39704 7392 39704 7392 0 _0023_
rlabel metal2 54768 9912 54768 9912 0 _0024_
rlabel metal2 61656 13440 61656 13440 0 _0025_
rlabel metal2 50792 17192 50792 17192 0 _0026_
rlabel metal2 52584 9352 52584 9352 0 _0027_
rlabel metal2 76160 24808 76160 24808 0 _0028_
rlabel metal2 75040 26376 75040 26376 0 _0029_
rlabel metal3 76888 21672 76888 21672 0 _0030_
rlabel metal2 77112 17024 77112 17024 0 _0031_
rlabel metal2 14504 35000 14504 35000 0 _0032_
rlabel metal2 24248 34552 24248 34552 0 _0033_
rlabel metal3 12376 33432 12376 33432 0 _0034_
rlabel metal3 12152 33544 12152 33544 0 _0035_
rlabel metal2 25480 35336 25480 35336 0 _0036_
rlabel metal2 20440 34496 20440 34496 0 _0037_
rlabel metal2 43232 31528 43232 31528 0 _0038_
rlabel metal3 59136 34776 59136 34776 0 _0039_
rlabel metal2 50008 33152 50008 33152 0 _0040_
rlabel metal3 45304 34216 45304 34216 0 _0041_
rlabel metal2 51912 33544 51912 33544 0 _0042_
rlabel metal2 52080 31080 52080 31080 0 _0043_
rlabel metal2 61656 32928 61656 32928 0 _0044_
rlabel metal3 60592 32760 60592 32760 0 _0045_
rlabel metal2 60984 32200 60984 32200 0 _0046_
rlabel metal2 53480 33320 53480 33320 0 _0047_
rlabel metal2 15400 10528 15400 10528 0 _0048_
rlabel metal2 24248 15540 24248 15540 0 _0049_
rlabel metal2 14560 16184 14560 16184 0 _0050_
rlabel metal2 14728 19992 14728 19992 0 _0051_
rlabel metal2 19656 9128 19656 9128 0 _0052_
rlabel metal2 21840 19320 21840 19320 0 _0053_
rlabel metal2 30520 10696 30520 10696 0 _0054_
rlabel metal2 39144 9464 39144 9464 0 _0055_
rlabel metal2 58576 10472 58576 10472 0 _0056_
rlabel metal2 66472 11032 66472 11032 0 _0057_
rlabel metal2 53424 19320 53424 19320 0 _0058_
rlabel metal2 51688 10920 51688 10920 0 _0059_
rlabel metal2 75712 29512 75712 29512 0 _0060_
rlabel metal2 74536 29904 74536 29904 0 _0061_
rlabel metal2 74424 22400 74424 22400 0 _0062_
rlabel metal2 77504 18536 77504 18536 0 _0063_
rlabel metal2 15400 4648 15400 4648 0 _0064_
rlabel metal2 20552 4424 20552 4424 0 _0065_
rlabel metal2 2744 19712 2744 19712 0 _0066_
rlabel metal2 3192 29736 3192 29736 0 _0067_
rlabel metal2 6328 12488 6328 12488 0 _0068_
rlabel metal2 9240 30688 9240 30688 0 _0069_
rlabel metal2 32760 5600 32760 5600 0 _0070_
rlabel metal2 39872 4536 39872 4536 0 _0071_
rlabel metal2 58072 5992 58072 5992 0 _0072_
rlabel metal2 66080 4424 66080 4424 0 _0073_
rlabel metal2 63112 17752 63112 17752 0 _0074_
rlabel metal2 48272 9912 48272 9912 0 _0075_
rlabel metal2 67368 35000 67368 35000 0 _0076_
rlabel metal2 70784 33432 70784 33432 0 _0077_
rlabel metal2 77112 12488 77112 12488 0 _0078_
rlabel metal2 72408 7896 72408 7896 0 _0079_
rlabel metal2 12824 4760 12824 4760 0 _0080_
rlabel metal2 29176 5376 29176 5376 0 _0081_
rlabel metal2 3304 16744 3304 16744 0 _0082_
rlabel metal2 2520 26600 2520 26600 0 _0083_
rlabel metal2 2688 9576 2688 9576 0 _0084_
rlabel metal2 7392 26488 7392 26488 0 _0085_
rlabel metal2 30408 4648 30408 4648 0 _0086_
rlabel metal3 48888 5992 48888 5992 0 _0087_
rlabel metal2 57400 4480 57400 4480 0 _0088_
rlabel metal3 63560 6664 63560 6664 0 _0089_
rlabel metal2 63112 21000 63112 21000 0 _0090_
rlabel metal3 48048 8344 48048 8344 0 _0091_
rlabel metal2 65408 29624 65408 29624 0 _0092_
rlabel metal2 71064 31416 71064 31416 0 _0093_
rlabel metal2 70448 12376 70448 12376 0 _0094_
rlabel metal2 70224 5208 70224 5208 0 _0095_
rlabel metal2 10360 4648 10360 4648 0 _0096_
rlabel metal2 26152 4760 26152 4760 0 _0097_
rlabel metal2 2744 15624 2744 15624 0 _0098_
rlabel metal2 2856 22624 2856 22624 0 _0099_
rlabel metal2 3864 7784 3864 7784 0 _0100_
rlabel metal2 6776 23352 6776 23352 0 _0101_
rlabel metal2 37688 4648 37688 4648 0 _0102_
rlabel metal2 48216 4760 48216 4760 0 _0103_
rlabel metal2 53088 4424 53088 4424 0 _0104_
rlabel metal2 61488 4424 61488 4424 0 _0105_
rlabel metal2 61320 18144 61320 18144 0 _0106_
rlabel metal2 45192 8260 45192 8260 0 _0107_
rlabel metal2 65520 31080 65520 31080 0 _0108_
rlabel metal2 69832 30688 69832 30688 0 _0109_
rlabel metal3 70560 14616 70560 14616 0 _0110_
rlabel metal2 68488 5488 68488 5488 0 _0111_
rlabel metal2 15624 7896 15624 7896 0 _0112_
rlabel metal2 22792 8736 22792 8736 0 _0113_
rlabel metal2 8288 13048 8288 13048 0 _0114_
rlabel metal2 10808 27216 10808 27216 0 _0115_
rlabel metal2 9520 9912 9520 9912 0 _0116_
rlabel metal2 11368 24192 11368 24192 0 _0117_
rlabel metal2 33768 10304 33768 10304 0 _0118_
rlabel metal2 43848 6216 43848 6216 0 _0119_
rlabel metal2 57624 9352 57624 9352 0 _0120_
rlabel metal2 61824 9912 61824 9912 0 _0121_
rlabel metal3 58744 20104 58744 20104 0 _0122_
rlabel metal2 46872 17248 46872 17248 0 _0123_
rlabel metal2 63896 25144 63896 25144 0 _0124_
rlabel metal2 66808 23464 66808 23464 0 _0125_
rlabel metal2 72632 18088 72632 18088 0 _0126_
rlabel metal2 69272 10192 69272 10192 0 _0127_
rlabel metal3 64568 8120 64568 8120 0 _0128_
rlabel metal2 66584 9072 66584 9072 0 _0129_
rlabel metal3 52472 20552 52472 20552 0 _0130_
rlabel metal3 58240 23688 58240 23688 0 _0131_
rlabel metal2 54488 34384 54488 34384 0 _0132_
rlabel metal2 54152 34048 54152 34048 0 _0133_
rlabel metal2 53816 32200 53816 32200 0 _0134_
rlabel metal2 51968 21784 51968 21784 0 _0135_
rlabel metal3 58240 23800 58240 23800 0 _0136_
rlabel metal2 52696 21112 52696 21112 0 _0137_
rlabel metal2 59416 19544 59416 19544 0 _0138_
rlabel metal2 65520 20104 65520 20104 0 _0139_
rlabel metal2 71064 34104 71064 34104 0 _0140_
rlabel metal3 64176 20104 64176 20104 0 _0141_
rlabel metal2 50736 20552 50736 20552 0 _0142_
rlabel metal2 55496 33712 55496 33712 0 _0143_
rlabel metal2 54824 30968 54824 30968 0 _0144_
rlabel metal2 51240 23016 51240 23016 0 _0145_
rlabel metal2 50792 21112 50792 21112 0 _0146_
rlabel metal2 48664 17920 48664 17920 0 _0147_
rlabel metal2 45976 10304 45976 10304 0 _0148_
rlabel metal2 45416 13440 45416 13440 0 _0149_
rlabel metal2 60368 23352 60368 23352 0 _0150_
rlabel metal3 57232 33320 57232 33320 0 _0151_
rlabel metal2 59640 28896 59640 28896 0 _0152_
rlabel metal2 62664 28392 62664 28392 0 _0153_
rlabel metal2 58744 24360 58744 24360 0 _0154_
rlabel metal2 68544 30184 68544 30184 0 _0155_
rlabel metal2 67256 29008 67256 29008 0 _0156_
rlabel metal3 65800 33544 65800 33544 0 _0157_
rlabel metal2 59752 23464 59752 23464 0 _0158_
rlabel metal2 57848 30912 57848 30912 0 _0159_
rlabel metal2 57624 31192 57624 31192 0 _0160_
rlabel metal2 57456 26264 57456 26264 0 _0161_
rlabel metal2 57736 23408 57736 23408 0 _0162_
rlabel metal2 71960 28056 71960 28056 0 _0163_
rlabel metal2 71064 32648 71064 32648 0 _0164_
rlabel metal3 70112 34104 70112 34104 0 _0165_
rlabel metal2 60928 22232 60928 22232 0 _0166_
rlabel metal2 59864 24248 59864 24248 0 _0167_
rlabel metal3 60200 21784 60200 21784 0 _0168_
rlabel metal2 75656 22624 75656 22624 0 _0169_
rlabel metal2 74200 15680 74200 15680 0 _0170_
rlabel metal2 73640 14728 73640 14728 0 _0171_
rlabel metal2 57176 33768 57176 33768 0 _0172_
rlabel metal2 52920 25760 52920 25760 0 _0173_
rlabel metal2 51688 22008 51688 22008 0 _0174_
rlabel metal2 68152 11144 68152 11144 0 _0175_
rlabel metal2 76440 17752 76440 17752 0 _0176_
rlabel metal2 72856 10472 72856 10472 0 _0177_
rlabel metal2 44296 17976 44296 17976 0 _0178_
rlabel metal2 41832 16520 41832 16520 0 _0179_
rlabel metal2 76328 20356 76328 20356 0 _0180_
rlabel metal2 41328 15400 41328 15400 0 _0181_
rlabel metal3 11480 7560 11480 7560 0 _0182_
rlabel metal2 26544 8456 26544 8456 0 _0183_
rlabel metal2 7784 16912 7784 16912 0 _0184_
rlabel metal3 5432 20664 5432 20664 0 _0185_
rlabel metal2 40768 16744 40768 16744 0 _0186_
rlabel metal2 7560 6160 7560 6160 0 _0187_
rlabel metal2 7840 20216 7840 20216 0 _0188_
rlabel metal2 31080 8344 31080 8344 0 _0189_
rlabel metal2 39368 7224 39368 7224 0 _0190_
rlabel metal2 62440 18088 62440 18088 0 _0191_
rlabel metal2 54880 10808 54880 10808 0 _0192_
rlabel metal2 62216 13048 62216 13048 0 _0193_
rlabel metal3 52080 17528 52080 17528 0 _0194_
rlabel metal2 52920 9688 52920 9688 0 _0195_
rlabel metal2 76888 25424 76888 25424 0 _0196_
rlabel metal2 76384 25704 76384 25704 0 _0197_
rlabel metal2 74424 27552 74424 27552 0 _0198_
rlabel metal2 78120 22624 78120 22624 0 _0199_
rlabel metal2 75936 17416 75936 17416 0 _0200_
rlabel metal2 76888 17640 76888 17640 0 _0201_
rlabel metal2 13720 30660 13720 30660 0 _0202_
rlabel metal2 20664 33432 20664 33432 0 _0203_
rlabel metal2 15456 33544 15456 33544 0 _0204_
rlabel metal2 16744 32704 16744 32704 0 _0205_
rlabel metal3 19152 33992 19152 33992 0 _0206_
rlabel metal2 23576 33376 23576 33376 0 _0207_
rlabel metal2 26376 32872 26376 32872 0 _0208_
rlabel metal2 23688 33768 23688 33768 0 _0209_
rlabel metal2 18984 33264 18984 33264 0 _0210_
rlabel metal2 14952 32228 14952 32228 0 _0211_
rlabel metal3 16128 33208 16128 33208 0 _0212_
rlabel metal3 14896 32536 14896 32536 0 _0213_
rlabel metal2 12712 32984 12712 32984 0 _0214_
rlabel metal2 25368 32872 25368 32872 0 _0215_
rlabel metal2 25480 34104 25480 34104 0 _0216_
rlabel metal2 20496 33096 20496 33096 0 _0217_
rlabel metal3 21000 34104 21000 34104 0 _0218_
rlabel metal2 43176 31808 43176 31808 0 _0219_
rlabel metal2 43064 29400 43064 29400 0 _0220_
rlabel metal2 23464 30240 23464 30240 0 _0221_
rlabel metal2 37576 25592 37576 25592 0 _0222_
rlabel metal2 37128 25032 37128 25032 0 _0223_
rlabel metal2 37520 31528 37520 31528 0 _0224_
rlabel metal3 35392 29400 35392 29400 0 _0225_
rlabel metal2 36792 26628 36792 26628 0 _0226_
rlabel metal3 44856 26544 44856 26544 0 _0227_
rlabel metal2 45416 27552 45416 27552 0 _0228_
rlabel metal2 44184 28728 44184 28728 0 _0229_
rlabel metal2 43008 29624 43008 29624 0 _0230_
rlabel metal2 44968 32648 44968 32648 0 _0231_
rlabel metal2 46200 28168 46200 28168 0 _0232_
rlabel metal2 45416 25872 45416 25872 0 _0233_
rlabel metal2 45024 25256 45024 25256 0 _0234_
rlabel metal2 46368 26040 46368 26040 0 _0235_
rlabel metal2 46200 26600 46200 26600 0 _0236_
rlabel metal2 47320 28672 47320 28672 0 _0237_
rlabel metal2 46424 28560 46424 28560 0 _0238_
rlabel metal2 46088 29344 46088 29344 0 _0239_
rlabel metal2 44072 30296 44072 30296 0 _0240_
rlabel metal2 57624 34104 57624 34104 0 _0241_
rlabel metal2 49448 31360 49448 31360 0 _0242_
rlabel metal2 49728 31192 49728 31192 0 _0243_
rlabel metal2 49224 27384 49224 27384 0 _0244_
rlabel metal2 48664 24640 48664 24640 0 _0245_
rlabel metal2 50904 25144 50904 25144 0 _0246_
rlabel metal2 52584 26572 52584 26572 0 _0247_
rlabel metal2 50344 30296 50344 30296 0 _0248_
rlabel metal2 48216 25480 48216 25480 0 _0249_
rlabel metal2 49448 25536 49448 25536 0 _0250_
rlabel metal2 48664 29008 48664 29008 0 _0251_
rlabel metal2 47768 29568 47768 29568 0 _0252_
rlabel metal2 46872 30632 46872 30632 0 _0253_
rlabel metal2 43792 31192 43792 31192 0 _0254_
rlabel metal2 44296 33432 44296 33432 0 _0255_
rlabel metal2 51688 31864 51688 31864 0 _0256_
rlabel metal2 48328 29176 48328 29176 0 _0257_
rlabel metal2 49672 29624 49672 29624 0 _0258_
rlabel metal2 51464 28896 51464 28896 0 _0259_
rlabel metal2 52024 28896 52024 28896 0 _0260_
rlabel metal2 51912 30464 51912 30464 0 _0261_
rlabel metal2 51800 31248 51800 31248 0 _0262_
rlabel metal2 53704 29512 53704 29512 0 _0263_
rlabel metal2 54264 29680 54264 29680 0 _0264_
rlabel metal2 53816 27832 53816 27832 0 _0265_
rlabel metal2 53592 28000 53592 28000 0 _0266_
rlabel metal2 53032 29344 53032 29344 0 _0267_
rlabel metal2 46648 32200 46648 32200 0 _0268_
rlabel metal2 55048 27776 55048 27776 0 _0269_
rlabel metal3 55440 28504 55440 28504 0 _0270_
rlabel metal2 62776 29456 62776 29456 0 _0271_
rlabel metal2 62104 29008 62104 29008 0 _0272_
rlabel metal2 63000 28952 63000 28952 0 _0273_
rlabel metal2 62664 29904 62664 29904 0 _0274_
rlabel metal2 61320 30968 61320 30968 0 _0275_
rlabel metal2 58296 28896 58296 28896 0 _0276_
rlabel metal2 57064 26600 57064 26600 0 _0277_
rlabel metal3 60480 28840 60480 28840 0 _0278_
rlabel metal2 62328 29008 62328 29008 0 _0279_
rlabel metal2 59304 29008 59304 29008 0 _0280_
rlabel metal2 58128 28728 58128 28728 0 _0281_
rlabel metal2 57624 28448 57624 28448 0 _0282_
rlabel metal2 57512 29008 57512 29008 0 _0283_
rlabel metal2 59752 29848 59752 29848 0 _0284_
rlabel metal2 60088 30352 60088 30352 0 _0285_
rlabel metal2 59808 26264 59808 26264 0 _0286_
rlabel metal2 58856 27552 58856 27552 0 _0287_
rlabel metal2 59360 26376 59360 26376 0 _0288_
rlabel metal2 59696 26488 59696 26488 0 _0289_
rlabel metal2 59472 27160 59472 27160 0 _0290_
rlabel metal2 60088 31416 60088 31416 0 _0291_
rlabel metal3 52472 30968 52472 30968 0 _0292_
rlabel metal2 58408 24864 58408 24864 0 _0293_
rlabel metal3 57120 24808 57120 24808 0 _0294_
rlabel metal2 55608 25928 55608 25928 0 _0295_
rlabel metal2 52808 26684 52808 26684 0 _0296_
rlabel metal2 41608 19768 41608 19768 0 _0297_
rlabel metal2 24136 17360 24136 17360 0 _0298_
rlabel metal2 23576 16464 23576 16464 0 _0299_
rlabel metal2 74200 20356 74200 20356 0 _0300_
rlabel metal2 24248 18928 24248 18928 0 _0301_
rlabel metal3 16632 10808 16632 10808 0 _0302_
rlabel metal3 25144 16968 25144 16968 0 _0303_
rlabel metal2 24136 16072 24136 16072 0 _0304_
rlabel metal2 14952 15736 14952 15736 0 _0305_
rlabel metal2 15288 19600 15288 19600 0 _0306_
rlabel metal2 20328 9800 20328 9800 0 _0307_
rlabel metal2 22232 19880 22232 19880 0 _0308_
rlabel metal2 31192 10584 31192 10584 0 _0309_
rlabel metal2 39368 9688 39368 9688 0 _0310_
rlabel metal2 65688 18424 65688 18424 0 _0311_
rlabel metal2 58072 11368 58072 11368 0 _0312_
rlabel metal3 66416 10584 66416 10584 0 _0313_
rlabel metal2 53816 18536 53816 18536 0 _0314_
rlabel metal3 52472 11256 52472 11256 0 _0315_
rlabel metal2 77000 27832 77000 27832 0 _0316_
rlabel metal3 75880 30072 75880 30072 0 _0317_
rlabel metal2 74312 29680 74312 29680 0 _0318_
rlabel metal2 74760 21728 74760 21728 0 _0319_
rlabel metal3 76664 19096 76664 19096 0 _0320_
rlabel metal3 76272 18984 76272 18984 0 _0321_
rlabel metal2 46984 17136 46984 17136 0 _0322_
rlabel metal2 46536 15932 46536 15932 0 _0323_
rlabel metal3 48272 2520 48272 2520 0 _0324_
rlabel metal2 15736 5376 15736 5376 0 _0325_
rlabel metal2 20776 5376 20776 5376 0 _0326_
rlabel metal3 7000 29288 7000 29288 0 _0327_
rlabel metal2 4760 19376 4760 19376 0 _0328_
rlabel metal2 5768 29848 5768 29848 0 _0329_
rlabel metal2 6608 11592 6608 11592 0 _0330_
rlabel metal2 9688 30296 9688 30296 0 _0331_
rlabel metal2 42840 5376 42840 5376 0 _0332_
rlabel metal3 33992 5880 33992 5880 0 _0333_
rlabel metal3 40712 4312 40712 4312 0 _0334_
rlabel metal3 58240 6664 58240 6664 0 _0335_
rlabel metal2 66696 5600 66696 5600 0 _0336_
rlabel metal2 70504 32480 70504 32480 0 _0337_
rlabel metal2 63896 18144 63896 18144 0 _0338_
rlabel metal2 47880 10920 47880 10920 0 _0339_
rlabel metal2 67816 34020 67816 34020 0 _0340_
rlabel metal2 71624 34216 71624 34216 0 _0341_
rlabel metal2 75096 12824 75096 12824 0 _0342_
rlabel metal2 72744 8344 72744 8344 0 _0343_
rlabel metal3 46760 15512 46760 15512 0 _0344_
rlabel metal3 28392 2968 28392 2968 0 _0345_
rlabel metal3 49672 2632 49672 2632 0 _0346_
rlabel metal2 13160 4648 13160 4648 0 _0347_
rlabel metal2 29512 5376 29512 5376 0 _0348_
rlabel metal2 8064 17416 8064 17416 0 _0349_
rlabel metal3 4760 16072 4760 16072 0 _0350_
rlabel metal2 3304 26376 3304 26376 0 _0351_
rlabel metal3 3528 9688 3528 9688 0 _0352_
rlabel metal2 7448 26264 7448 26264 0 _0353_
rlabel metal2 49224 6496 49224 6496 0 _0354_
rlabel metal2 33320 4760 33320 4760 0 _0355_
rlabel metal2 47992 6160 47992 6160 0 _0356_
rlabel metal3 58520 5096 58520 5096 0 _0357_
rlabel metal2 62664 6776 62664 6776 0 _0358_
rlabel metal2 72856 29680 72856 29680 0 _0359_
rlabel metal2 61768 20776 61768 20776 0 _0360_
rlabel metal3 48552 9016 48552 9016 0 _0361_
rlabel metal2 66024 29400 66024 29400 0 _0362_
rlabel metal3 72576 30184 72576 30184 0 _0363_
rlabel metal3 71624 12264 71624 12264 0 _0364_
rlabel metal2 72184 6384 72184 6384 0 _0365_
rlabel metal2 44968 16800 44968 16800 0 _0366_
rlabel metal3 30576 2744 30576 2744 0 _0367_
rlabel metal3 50120 2856 50120 2856 0 _0368_
rlabel metal2 9016 5376 9016 5376 0 _0369_
rlabel metal2 26712 4312 26712 4312 0 _0370_
rlabel metal3 9184 23352 9184 23352 0 _0371_
rlabel metal2 5320 15736 5320 15736 0 _0372_
rlabel metal3 3528 22232 3528 22232 0 _0373_
rlabel metal2 5992 8512 5992 8512 0 _0374_
rlabel metal3 8176 23240 8176 23240 0 _0375_
rlabel metal2 38696 5432 38696 5432 0 _0376_
rlabel metal3 36288 5096 36288 5096 0 _0377_
rlabel metal3 48440 4312 48440 4312 0 _0378_
rlabel metal3 53928 5096 53928 5096 0 _0379_
rlabel metal2 62216 5600 62216 5600 0 _0380_
rlabel metal2 69720 28952 69720 28952 0 _0381_
rlabel metal2 60536 18368 60536 18368 0 _0382_
rlabel metal2 44968 8904 44968 8904 0 _0383_
rlabel metal2 66360 29400 66360 29400 0 _0384_
rlabel metal2 70168 30296 70168 30296 0 _0385_
rlabel metal2 69832 15204 69832 15204 0 _0386_
rlabel metal3 68488 5096 68488 5096 0 _0387_
rlabel metal3 46760 17640 46760 17640 0 _0388_
rlabel metal2 45528 17416 45528 17416 0 _0389_
rlabel metal2 19544 7952 19544 7952 0 _0390_
rlabel metal2 15960 7784 15960 7784 0 _0391_
rlabel metal2 23464 8344 23464 8344 0 _0392_
rlabel metal2 13608 23296 13608 23296 0 _0393_
rlabel metal2 9240 13720 9240 13720 0 _0394_
rlabel metal2 11704 26768 11704 26768 0 _0395_
rlabel metal2 9688 9464 9688 9464 0 _0396_
rlabel metal2 11704 24192 11704 24192 0 _0397_
rlabel metal2 44072 7840 44072 7840 0 _0398_
rlabel metal2 34552 9912 34552 9912 0 _0399_
rlabel metal2 43232 6664 43232 6664 0 _0400_
rlabel metal2 57848 9072 57848 9072 0 _0401_
rlabel metal2 61992 9912 61992 9912 0 _0402_
rlabel metal2 49280 17752 49280 17752 0 _0403_
rlabel metal2 58240 19432 58240 19432 0 _0404_
rlabel metal2 47432 17528 47432 17528 0 _0405_
rlabel metal3 64288 24696 64288 24696 0 _0406_
rlabel metal2 66472 23184 66472 23184 0 _0407_
rlabel metal3 71960 16968 71960 16968 0 _0408_
rlabel metal2 69608 9968 69608 9968 0 _0409_
rlabel via2 27496 19992 27496 19992 0 _0410_
rlabel metal3 31472 19208 31472 19208 0 _0411_
rlabel metal2 33768 20440 33768 20440 0 _0412_
rlabel metal2 37352 18760 37352 18760 0 _0413_
rlabel metal2 16912 10024 16912 10024 0 _0414_
rlabel metal2 40264 20776 40264 20776 0 _0415_
rlabel metal3 26628 23800 26628 23800 0 _0416_
rlabel metal2 33656 22064 33656 22064 0 _0417_
rlabel metal3 35840 22232 35840 22232 0 _0418_
rlabel metal2 42728 20944 42728 20944 0 _0419_
rlabel metal2 37240 17528 37240 17528 0 _0420_
rlabel metal2 39368 23352 39368 23352 0 _0421_
rlabel metal2 30296 21392 30296 21392 0 _0422_
rlabel metal2 37576 20160 37576 20160 0 _0423_
rlabel metal2 40600 19376 40600 19376 0 _0424_
rlabel metal2 38584 18704 38584 18704 0 _0425_
rlabel metal2 33544 16800 33544 16800 0 _0426_
rlabel metal3 20328 17360 20328 17360 0 _0427_
rlabel metal2 26544 16072 26544 16072 0 _0428_
rlabel metal2 38752 17528 38752 17528 0 _0429_
rlabel metal2 34328 17752 34328 17752 0 _0430_
rlabel metal2 43288 17416 43288 17416 0 _0431_
rlabel metal2 40264 17752 40264 17752 0 _0432_
rlabel metal3 39396 20664 39396 20664 0 _0433_
rlabel metal2 36232 17584 36232 17584 0 _0434_
rlabel metal2 37632 17752 37632 17752 0 _0435_
rlabel metal2 18760 16408 18760 16408 0 _0436_
rlabel metal2 41104 15288 41104 15288 0 _0437_
rlabel metal3 21896 15512 21896 15512 0 _0438_
rlabel metal2 20216 12544 20216 12544 0 _0439_
rlabel metal3 32144 17080 32144 17080 0 _0440_
rlabel metal2 23688 16744 23688 16744 0 _0441_
rlabel metal2 18088 12712 18088 12712 0 _0442_
rlabel metal2 16520 11424 16520 11424 0 _0443_
rlabel metal2 17304 11536 17304 11536 0 _0444_
rlabel metal2 12936 12376 12936 12376 0 _0445_
rlabel metal3 40488 14504 40488 14504 0 _0446_
rlabel metal2 29624 15232 29624 15232 0 _0447_
rlabel metal2 38920 18872 38920 18872 0 _0448_
rlabel metal3 38892 16072 38892 16072 0 _0449_
rlabel metal3 20440 15848 20440 15848 0 _0450_
rlabel metal2 15400 18032 15400 18032 0 _0451_
rlabel metal2 18088 10976 18088 10976 0 _0452_
rlabel metal3 37296 15176 37296 15176 0 _0453_
rlabel metal2 39480 20720 39480 20720 0 _0454_
rlabel metal2 35672 16464 35672 16464 0 _0455_
rlabel metal3 36288 16744 36288 16744 0 _0456_
rlabel metal3 32480 17528 32480 17528 0 _0457_
rlabel metal2 30296 16016 30296 16016 0 _0458_
rlabel metal2 29400 16968 29400 16968 0 _0459_
rlabel metal2 13608 17808 13608 17808 0 _0460_
rlabel metal2 11928 12432 11928 12432 0 _0461_
rlabel metal2 25032 17808 25032 17808 0 _0462_
rlabel metal2 25480 13552 25480 13552 0 _0463_
rlabel metal2 14280 12432 14280 12432 0 _0464_
rlabel metal2 18648 12096 18648 12096 0 _0465_
rlabel metal2 21560 13328 21560 13328 0 _0466_
rlabel metal2 18984 12992 18984 12992 0 _0467_
rlabel metal2 17976 15624 17976 15624 0 _0468_
rlabel metal3 18368 12824 18368 12824 0 _0469_
rlabel metal2 18872 12040 18872 12040 0 _0470_
rlabel metal3 19768 9856 19768 9856 0 _0471_
rlabel metal3 62636 22344 62636 22344 0 _0472_
rlabel metal2 54432 23912 54432 23912 0 _0473_
rlabel metal2 58296 22176 58296 22176 0 _0474_
rlabel metal2 55440 23240 55440 23240 0 _0475_
rlabel metal3 41328 13832 41328 13832 0 _0476_
rlabel metal2 25032 19824 25032 19824 0 _0477_
rlabel metal2 53592 23520 53592 23520 0 _0478_
rlabel metal3 55216 24024 55216 24024 0 _0479_
rlabel metal2 58184 22344 58184 22344 0 _0480_
rlabel metal2 57176 23744 57176 23744 0 _0481_
rlabel metal3 40152 13944 40152 13944 0 _0482_
rlabel metal3 26152 20608 26152 20608 0 _0483_
rlabel metal3 16016 12712 16016 12712 0 _0484_
rlabel metal3 18200 22176 18200 22176 0 _0485_
rlabel metal2 12880 14280 12880 14280 0 _0486_
rlabel metal3 47320 9744 47320 9744 0 _0487_
rlabel metal2 10920 16744 10920 16744 0 _0488_
rlabel metal3 21000 14728 21000 14728 0 _0489_
rlabel metal2 10584 16576 10584 16576 0 _0490_
rlabel metal3 15512 14056 15512 14056 0 _0491_
rlabel metal2 57176 24640 57176 24640 0 _0492_
rlabel metal2 21112 21224 21112 21224 0 _0493_
rlabel metal2 17416 14112 17416 14112 0 _0494_
rlabel metal2 19376 20552 19376 20552 0 _0495_
rlabel metal3 17416 13944 17416 13944 0 _0496_
rlabel metal3 16912 13720 16912 13720 0 _0497_
rlabel metal2 15848 24136 15848 24136 0 _0498_
rlabel metal2 26264 21000 26264 21000 0 _0499_
rlabel metal2 25592 22568 25592 22568 0 _0500_
rlabel metal2 26824 20888 26824 20888 0 _0501_
rlabel metal3 30128 23912 30128 23912 0 _0502_
rlabel metal3 26572 26376 26572 26376 0 _0503_
rlabel metal2 24472 27720 24472 27720 0 _0504_
rlabel metal2 14280 28336 14280 28336 0 _0505_
rlabel metal3 18648 23912 18648 23912 0 _0506_
rlabel metal2 27496 21952 27496 21952 0 _0507_
rlabel metal2 28168 25368 28168 25368 0 _0508_
rlabel metal2 24248 25872 24248 25872 0 _0509_
rlabel metal2 25480 31920 25480 31920 0 _0510_
rlabel metal2 29960 19656 29960 19656 0 _0511_
rlabel metal3 31024 18424 31024 18424 0 _0512_
rlabel metal2 26376 25536 26376 25536 0 _0513_
rlabel metal2 21896 25368 21896 25368 0 _0514_
rlabel metal2 16632 25368 16632 25368 0 _0515_
rlabel metal3 28672 18424 28672 18424 0 _0516_
rlabel metal2 41496 21280 41496 21280 0 _0517_
rlabel metal2 19656 24696 19656 24696 0 _0518_
rlabel metal2 44464 37240 44464 37240 0 _0519_
rlabel metal2 28056 21560 28056 21560 0 _0520_
rlabel metal2 31304 23576 31304 23576 0 _0521_
rlabel metal2 26600 28392 26600 28392 0 _0522_
rlabel metal2 47096 22568 47096 22568 0 _0523_
rlabel metal2 19768 24864 19768 24864 0 _0524_
rlabel metal3 19096 24696 19096 24696 0 _0525_
rlabel metal2 26712 26208 26712 26208 0 _0526_
rlabel metal2 18088 24696 18088 24696 0 _0527_
rlabel metal3 18648 26040 18648 26040 0 _0528_
rlabel metal2 19208 25424 19208 25424 0 _0529_
rlabel metal2 19096 24192 19096 24192 0 _0530_
rlabel metal2 27888 10808 27888 10808 0 _0531_
rlabel metal2 26824 12712 26824 12712 0 _0532_
rlabel metal2 27048 12432 27048 12432 0 _0533_
rlabel metal3 28448 12264 28448 12264 0 _0534_
rlabel metal3 27272 13608 27272 13608 0 _0535_
rlabel metal3 16352 17528 16352 17528 0 _0536_
rlabel metal3 23240 13832 23240 13832 0 _0537_
rlabel metal3 25256 13496 25256 13496 0 _0538_
rlabel metal2 25536 13944 25536 13944 0 _0539_
rlabel metal2 20440 16016 20440 16016 0 _0540_
rlabel metal2 26488 15456 26488 15456 0 _0541_
rlabel metal2 25760 15288 25760 15288 0 _0542_
rlabel metal3 24136 15288 24136 15288 0 _0543_
rlabel metal2 26712 14784 26712 14784 0 _0544_
rlabel metal2 27608 13272 27608 13272 0 _0545_
rlabel metal2 29288 11760 29288 11760 0 _0546_
rlabel metal2 41440 12376 41440 12376 0 _0547_
rlabel metal2 25424 11368 25424 11368 0 _0548_
rlabel metal2 26040 12320 26040 12320 0 _0549_
rlabel metal2 25816 10080 25816 10080 0 _0550_
rlabel metal2 24472 11480 24472 11480 0 _0551_
rlabel metal2 25480 10864 25480 10864 0 _0552_
rlabel metal2 25816 11816 25816 11816 0 _0553_
rlabel metal2 24696 12320 24696 12320 0 _0554_
rlabel metal2 24248 11928 24248 11928 0 _0555_
rlabel metal3 25032 12152 25032 12152 0 _0556_
rlabel metal2 23800 23632 23800 23632 0 _0557_
rlabel metal2 22456 23520 22456 23520 0 _0558_
rlabel metal2 22904 25088 22904 25088 0 _0559_
rlabel metal3 23184 23800 23184 23800 0 _0560_
rlabel metal2 44072 24304 44072 24304 0 _0561_
rlabel metal2 23464 24192 23464 24192 0 _0562_
rlabel metal3 22064 26936 22064 26936 0 _0563_
rlabel metal2 22680 25816 22680 25816 0 _0564_
rlabel metal2 27776 27048 27776 27048 0 _0565_
rlabel metal2 25928 25144 25928 25144 0 _0566_
rlabel metal2 22456 25536 22456 25536 0 _0567_
rlabel metal2 19824 25592 19824 25592 0 _0568_
rlabel metal3 21224 25480 21224 25480 0 _0569_
rlabel metal3 22624 27048 22624 27048 0 _0570_
rlabel metal2 3080 34552 3080 34552 0 _0571_
rlabel metal2 15624 16464 15624 16464 0 _0572_
rlabel metal2 21448 17976 21448 17976 0 _0573_
rlabel metal2 17080 16744 17080 16744 0 _0574_
rlabel metal2 17528 16240 17528 16240 0 _0575_
rlabel metal3 13384 15176 13384 15176 0 _0576_
rlabel metal2 10472 15568 10472 15568 0 _0577_
rlabel metal2 33096 16464 33096 16464 0 _0578_
rlabel metal2 15176 9520 15176 9520 0 _0579_
rlabel metal2 13608 16240 13608 16240 0 _0580_
rlabel metal2 12264 15624 12264 15624 0 _0581_
rlabel metal2 18088 16576 18088 16576 0 _0582_
rlabel metal2 18872 14504 18872 14504 0 _0583_
rlabel metal2 17752 14784 17752 14784 0 _0584_
rlabel metal2 18760 16744 18760 16744 0 _0585_
rlabel metal3 22512 13944 22512 13944 0 _0586_
rlabel metal2 23128 23856 23128 23856 0 _0587_
rlabel metal3 20888 30072 20888 30072 0 _0588_
rlabel metal2 26040 25648 26040 25648 0 _0589_
rlabel metal2 16184 16520 16184 16520 0 _0590_
rlabel metal3 16296 17024 16296 17024 0 _0591_
rlabel metal3 16800 16856 16800 16856 0 _0592_
rlabel metal2 16856 17584 16856 17584 0 _0593_
rlabel metal3 18480 27832 18480 27832 0 _0594_
rlabel metal2 19208 17472 19208 17472 0 _0595_
rlabel metal2 18760 27216 18760 27216 0 _0596_
rlabel metal2 47880 25536 47880 25536 0 _0597_
rlabel metal2 20216 27608 20216 27608 0 _0598_
rlabel metal2 19880 28336 19880 28336 0 _0599_
rlabel metal3 21224 30184 21224 30184 0 _0600_
rlabel metal2 19208 29848 19208 29848 0 _0601_
rlabel metal2 20776 30688 20776 30688 0 _0602_
rlabel metal3 19992 31080 19992 31080 0 _0603_
rlabel metal2 20440 31528 20440 31528 0 _0604_
rlabel metal2 18536 29064 18536 29064 0 _0605_
rlabel metal2 25872 28616 25872 28616 0 _0606_
rlabel metal2 17920 31192 17920 31192 0 _0607_
rlabel metal2 17640 28728 17640 28728 0 _0608_
rlabel metal2 18088 30912 18088 30912 0 _0609_
rlabel metal2 18872 32144 18872 32144 0 _0610_
rlabel metal2 16856 19152 16856 19152 0 _0611_
rlabel metal2 22120 16968 22120 16968 0 _0612_
rlabel metal2 17416 18648 17416 18648 0 _0613_
rlabel metal2 17752 18816 17752 18816 0 _0614_
rlabel metal2 14728 18424 14728 18424 0 _0615_
rlabel metal3 10136 20328 10136 20328 0 _0616_
rlabel metal2 12376 18760 12376 18760 0 _0617_
rlabel metal3 17360 17864 17360 17864 0 _0618_
rlabel metal2 18872 18368 18872 18368 0 _0619_
rlabel metal2 16744 18200 16744 18200 0 _0620_
rlabel metal2 18312 19432 18312 19432 0 _0621_
rlabel metal2 76664 9800 76664 9800 0 _0622_
rlabel metal2 14952 29064 14952 29064 0 _0623_
rlabel metal2 17304 21224 17304 21224 0 _0624_
rlabel metal2 15736 21056 15736 21056 0 _0625_
rlabel metal3 16296 21672 16296 21672 0 _0626_
rlabel metal2 15176 22960 15176 22960 0 _0627_
rlabel metal2 14392 30128 14392 30128 0 _0628_
rlabel metal2 13664 28840 13664 28840 0 _0629_
rlabel metal2 16968 19880 16968 19880 0 _0630_
rlabel metal3 21616 29400 21616 29400 0 _0631_
rlabel metal2 13160 29848 13160 29848 0 _0632_
rlabel metal2 15736 28840 15736 28840 0 _0633_
rlabel metal2 14504 30800 14504 30800 0 _0634_
rlabel metal2 14840 31248 14840 31248 0 _0635_
rlabel metal2 17080 29736 17080 29736 0 _0636_
rlabel metal2 18536 26236 18536 26236 0 _0637_
rlabel metal2 19880 9912 19880 9912 0 _0638_
rlabel metal2 20664 12320 20664 12320 0 _0639_
rlabel metal2 20888 12264 20888 12264 0 _0640_
rlabel metal2 12936 10808 12936 10808 0 _0641_
rlabel metal2 12152 10752 12152 10752 0 _0642_
rlabel metal2 14280 10864 14280 10864 0 _0643_
rlabel metal2 21336 11900 21336 11900 0 _0644_
rlabel metal2 21168 12712 21168 12712 0 _0645_
rlabel metal2 20720 10584 20720 10584 0 _0646_
rlabel metal2 21784 11816 21784 11816 0 _0647_
rlabel metal2 76440 10976 76440 10976 0 _0648_
rlabel metal2 38808 21000 38808 21000 0 _0649_
rlabel metal2 39144 30856 39144 30856 0 _0650_
rlabel metal2 23912 10472 23912 10472 0 _0651_
rlabel metal3 24136 10752 24136 10752 0 _0652_
rlabel metal2 24248 10892 24248 10892 0 _0653_
rlabel metal2 24752 10808 24752 10808 0 _0654_
rlabel metal3 25480 27160 25480 27160 0 _0655_
rlabel metal2 22736 17752 22736 17752 0 _0656_
rlabel metal2 26376 27944 26376 27944 0 _0657_
rlabel metal2 26768 28392 26768 28392 0 _0658_
rlabel metal3 26488 29512 26488 29512 0 _0659_
rlabel metal2 24696 30912 24696 30912 0 _0660_
rlabel metal2 16520 30632 16520 30632 0 _0661_
rlabel metal2 17864 29400 17864 29400 0 _0662_
rlabel metal2 23576 31360 23576 31360 0 _0663_
rlabel metal2 25032 31360 25032 31360 0 _0664_
rlabel metal2 23912 31248 23912 31248 0 _0665_
rlabel metal3 25088 28056 25088 28056 0 _0666_
rlabel metal2 24024 31416 24024 31416 0 _0667_
rlabel metal2 25816 29568 25816 29568 0 _0668_
rlabel metal2 25928 30688 25928 30688 0 _0669_
rlabel metal3 22680 18984 22680 18984 0 _0670_
rlabel metal2 22568 18032 22568 18032 0 _0671_
rlabel metal2 22568 18480 22568 18480 0 _0672_
rlabel metal2 14840 19656 14840 19656 0 _0673_
rlabel metal3 10920 19992 10920 19992 0 _0674_
rlabel metal3 13048 17752 13048 17752 0 _0675_
rlabel metal2 23464 18592 23464 18592 0 _0676_
rlabel metal2 20104 18144 20104 18144 0 _0677_
rlabel metal2 20776 18424 20776 18424 0 _0678_
rlabel metal2 22680 18256 22680 18256 0 _0679_
rlabel metal3 26684 9464 26684 9464 0 _0680_
rlabel metal2 21448 21224 21448 21224 0 _0681_
rlabel metal2 19432 21504 19432 21504 0 _0682_
rlabel metal2 19544 21728 19544 21728 0 _0683_
rlabel metal2 20048 21784 20048 21784 0 _0684_
rlabel metal2 21896 29064 21896 29064 0 _0685_
rlabel metal2 21672 28056 21672 28056 0 _0686_
rlabel metal2 23800 18424 23800 18424 0 _0687_
rlabel metal2 23352 27832 23352 27832 0 _0688_
rlabel metal3 21280 29624 21280 29624 0 _0689_
rlabel metal3 21392 29512 21392 29512 0 _0690_
rlabel metal2 26712 31080 26712 31080 0 _0691_
rlabel metal2 23688 32088 23688 32088 0 _0692_
rlabel metal2 22960 31640 22960 31640 0 _0693_
rlabel metal2 22792 29120 22792 29120 0 _0694_
rlabel metal2 30688 11368 30688 11368 0 _0695_
rlabel metal2 32088 14392 32088 14392 0 _0696_
rlabel metal2 32536 16016 32536 16016 0 _0697_
rlabel metal2 31864 13328 31864 13328 0 _0698_
rlabel metal2 31304 13832 31304 13832 0 _0699_
rlabel metal2 32368 15960 32368 15960 0 _0700_
rlabel metal2 32760 16576 32760 16576 0 _0701_
rlabel metal3 33656 13608 33656 13608 0 _0702_
rlabel metal2 33320 15204 33320 15204 0 _0703_
rlabel metal3 32648 16296 32648 16296 0 _0704_
rlabel metal2 77000 16128 77000 16128 0 _0705_
rlabel metal2 46648 25592 46648 25592 0 _0706_
rlabel metal3 35000 12936 35000 12936 0 _0707_
rlabel metal2 32760 12992 32760 12992 0 _0708_
rlabel metal2 34552 13496 34552 13496 0 _0709_
rlabel metal2 33320 12768 33320 12768 0 _0710_
rlabel metal3 33488 20216 33488 20216 0 _0711_
rlabel metal2 34104 28168 34104 28168 0 _0712_
rlabel metal2 41384 27608 41384 27608 0 _0713_
rlabel metal2 30912 16632 30912 16632 0 _0714_
rlabel metal2 30240 27272 30240 27272 0 _0715_
rlabel metal2 29960 30576 29960 30576 0 _0716_
rlabel metal2 31640 31360 31640 31360 0 _0717_
rlabel metal2 23352 28280 23352 28280 0 _0718_
rlabel metal2 24752 28840 24752 28840 0 _0719_
rlabel metal3 29680 29624 29680 29624 0 _0720_
rlabel metal2 30520 31248 30520 31248 0 _0721_
rlabel metal2 30072 29400 30072 29400 0 _0722_
rlabel metal2 33208 31752 33208 31752 0 _0723_
rlabel metal2 31864 29512 31864 29512 0 _0724_
rlabel metal2 32424 29120 32424 29120 0 _0725_
rlabel metal2 34104 31080 34104 31080 0 _0726_
rlabel metal2 34888 28000 34888 28000 0 _0727_
rlabel metal2 33992 29680 33992 29680 0 _0728_
rlabel metal2 32200 23464 32200 23464 0 _0729_
rlabel metal2 52920 14728 52920 14728 0 _0730_
rlabel metal2 68712 15792 68712 15792 0 _0731_
rlabel metal2 46760 12096 46760 12096 0 _0732_
rlabel metal2 65576 16464 65576 16464 0 _0733_
rlabel metal2 48328 13272 48328 13272 0 _0734_
rlabel metal3 63952 15848 63952 15848 0 _0735_
rlabel metal2 49000 20440 49000 20440 0 _0736_
rlabel metal2 39704 13720 39704 13720 0 _0737_
rlabel metal3 43680 15176 43680 15176 0 _0738_
rlabel metal2 69216 15512 69216 15512 0 _0739_
rlabel metal3 48328 15736 48328 15736 0 _0740_
rlabel metal2 65576 15848 65576 15848 0 _0741_
rlabel metal2 40264 13496 40264 13496 0 _0742_
rlabel metal2 39480 12656 39480 12656 0 _0743_
rlabel metal2 41944 13776 41944 13776 0 _0744_
rlabel metal2 48776 19096 48776 19096 0 _0745_
rlabel metal2 32088 23240 32088 23240 0 _0746_
rlabel metal2 33656 24528 33656 24528 0 _0747_
rlabel metal2 47096 21000 47096 21000 0 _0748_
rlabel metal2 41720 10864 41720 10864 0 _0749_
rlabel metal2 41944 10752 41944 10752 0 _0750_
rlabel metal2 42280 10472 42280 10472 0 _0751_
rlabel metal2 37128 23632 37128 23632 0 _0752_
rlabel metal2 34104 24752 34104 24752 0 _0753_
rlabel metal3 35448 28392 35448 28392 0 _0754_
rlabel metal2 41048 22736 41048 22736 0 _0755_
rlabel metal2 33768 23436 33768 23436 0 _0756_
rlabel metal2 33320 28336 33320 28336 0 _0757_
rlabel metal2 31528 28336 31528 28336 0 _0758_
rlabel metal2 32312 27440 32312 27440 0 _0759_
rlabel metal3 31528 27608 31528 27608 0 _0760_
rlabel metal2 32536 26600 32536 26600 0 _0761_
rlabel metal2 33432 25424 33432 25424 0 _0762_
rlabel metal2 33992 26376 33992 26376 0 _0763_
rlabel metal2 2072 22680 2072 22680 0 _0764_
rlabel metal2 49672 15736 49672 15736 0 _0765_
rlabel metal2 66360 16128 66360 16128 0 _0766_
rlabel metal2 48888 15064 48888 15064 0 _0767_
rlabel metal2 63896 15568 63896 15568 0 _0768_
rlabel metal2 60256 12376 60256 12376 0 _0769_
rlabel metal2 59752 14616 59752 14616 0 _0770_
rlabel metal3 58912 15400 58912 15400 0 _0771_
rlabel metal2 49560 26432 49560 26432 0 _0772_
rlabel metal3 65912 17080 65912 17080 0 _0773_
rlabel metal3 65128 17416 65128 17416 0 _0774_
rlabel metal2 58856 14616 58856 14616 0 _0775_
rlabel metal2 67536 18424 67536 18424 0 _0776_
rlabel metal2 67872 18984 67872 18984 0 _0777_
rlabel metal2 57960 13888 57960 13888 0 _0778_
rlabel metal2 65744 15624 65744 15624 0 _0779_
rlabel metal3 57288 14392 57288 14392 0 _0780_
rlabel metal3 64624 15736 64624 15736 0 _0781_
rlabel metal2 64120 14784 64120 14784 0 _0782_
rlabel metal3 57232 13048 57232 13048 0 _0783_
rlabel metal2 52192 20776 52192 20776 0 _0784_
rlabel metal2 48552 30240 48552 30240 0 _0785_
rlabel metal3 41104 23240 41104 23240 0 _0786_
rlabel metal2 35728 24472 35728 24472 0 _0787_
rlabel metal2 31528 34048 31528 34048 0 _0788_
rlabel metal3 18088 29624 18088 29624 0 _0789_
rlabel metal3 24808 28448 24808 28448 0 _0790_
rlabel metal2 31192 29288 31192 29288 0 _0791_
rlabel metal2 31640 28896 31640 28896 0 _0792_
rlabel metal2 34664 28112 34664 28112 0 _0793_
rlabel metal2 33992 28672 33992 28672 0 _0794_
rlabel metal2 32424 34944 32424 34944 0 _0795_
rlabel metal2 31248 34888 31248 34888 0 _0796_
rlabel metal2 32872 34048 32872 34048 0 _0797_
rlabel metal2 32200 35840 32200 35840 0 _0798_
rlabel metal3 32592 31864 32592 31864 0 _0799_
rlabel metal2 31864 33320 31864 33320 0 _0800_
rlabel metal2 33320 32928 33320 32928 0 _0801_
rlabel metal2 66920 14840 66920 14840 0 _0802_
rlabel metal2 66136 14224 66136 14224 0 _0803_
rlabel metal2 65912 13384 65912 13384 0 _0804_
rlabel metal3 45752 29512 45752 29512 0 _0805_
rlabel metal2 65184 14616 65184 14616 0 _0806_
rlabel metal3 64568 13944 64568 13944 0 _0807_
rlabel metal2 64792 15204 64792 15204 0 _0808_
rlabel metal2 63112 24416 63112 24416 0 _0809_
rlabel metal2 46928 27832 46928 27832 0 _0810_
rlabel metal2 31472 24136 31472 24136 0 _0811_
rlabel metal2 28280 32760 28280 32760 0 _0812_
rlabel metal2 29400 33432 29400 33432 0 _0813_
rlabel metal3 30632 35672 30632 35672 0 _0814_
rlabel metal2 30968 34888 30968 34888 0 _0815_
rlabel metal2 30408 36120 30408 36120 0 _0816_
rlabel metal3 30072 34888 30072 34888 0 _0817_
rlabel metal2 29568 34104 29568 34104 0 _0818_
rlabel metal2 29400 34104 29400 34104 0 _0819_
rlabel metal3 44800 21560 44800 21560 0 _0820_
rlabel metal2 56952 17360 56952 17360 0 _0821_
rlabel metal2 55944 16912 55944 16912 0 _0822_
rlabel metal2 55496 17304 55496 17304 0 _0823_
rlabel metal2 50344 28280 50344 28280 0 _0824_
rlabel metal2 58856 18088 58856 18088 0 _0825_
rlabel metal3 56504 18424 56504 18424 0 _0826_
rlabel metal2 56952 18760 56952 18760 0 _0827_
rlabel metal2 57848 18032 57848 18032 0 _0828_
rlabel metal2 54208 24248 54208 24248 0 _0829_
rlabel metal2 41160 34272 41160 34272 0 _0830_
rlabel metal2 40264 23800 40264 23800 0 _0831_
rlabel metal2 40600 35336 40600 35336 0 _0832_
rlabel metal2 37744 35784 37744 35784 0 _0833_
rlabel metal2 37240 33096 37240 33096 0 _0834_
rlabel metal3 30016 33992 30016 33992 0 _0835_
rlabel metal2 33880 34440 33880 34440 0 _0836_
rlabel metal3 34888 33432 34888 33432 0 _0837_
rlabel metal3 37352 34888 37352 34888 0 _0838_
rlabel metal2 35896 34216 35896 34216 0 _0839_
rlabel metal2 37016 33208 37016 33208 0 _0840_
rlabel metal2 37912 32480 37912 32480 0 _0841_
rlabel metal2 49112 14616 49112 14616 0 _0842_
rlabel metal2 50232 13384 50232 13384 0 _0843_
rlabel metal2 47880 13888 47880 13888 0 _0844_
rlabel metal2 38584 35000 38584 35000 0 _0845_
rlabel metal2 41160 24500 41160 24500 0 _0846_
rlabel metal2 43400 27664 43400 27664 0 _0847_
rlabel metal2 43624 13104 43624 13104 0 _0848_
rlabel metal3 43400 13720 43400 13720 0 _0849_
rlabel metal2 43680 11480 43680 11480 0 _0850_
rlabel metal2 42336 19544 42336 19544 0 _0851_
rlabel metal2 39480 30800 39480 30800 0 _0852_
rlabel metal2 38920 33600 38920 33600 0 _0853_
rlabel metal2 39032 33824 39032 33824 0 _0854_
rlabel metal2 39312 34664 39312 34664 0 _0855_
rlabel metal2 38360 32592 38360 32592 0 _0856_
rlabel metal2 41272 34608 41272 34608 0 _0857_
rlabel metal2 39928 32592 39928 32592 0 _0858_
rlabel metal2 40936 22456 40936 22456 0 _0859_
rlabel metal3 40656 31192 40656 31192 0 _0860_
rlabel metal2 73136 27160 73136 27160 0 _0861_
rlabel metal2 69832 25368 69832 25368 0 _0862_
rlabel metal2 69216 25704 69216 25704 0 _0863_
rlabel metal2 73976 25872 73976 25872 0 _0864_
rlabel metal2 71512 17584 71512 17584 0 _0865_
rlabel metal2 67704 16856 67704 16856 0 _0866_
rlabel metal2 70056 26544 70056 26544 0 _0867_
rlabel metal2 69272 25536 69272 25536 0 _0868_
rlabel metal2 71512 16856 71512 16856 0 _0869_
rlabel metal2 69720 26264 69720 26264 0 _0870_
rlabel metal2 62552 28112 62552 28112 0 _0871_
rlabel metal3 64400 23240 64400 23240 0 _0872_
rlabel metal3 62552 24584 62552 24584 0 _0873_
rlabel metal2 69440 20216 69440 20216 0 _0874_
rlabel metal2 67032 18312 67032 18312 0 _0875_
rlabel metal2 67536 27048 67536 27048 0 _0876_
rlabel metal3 69048 27832 69048 27832 0 _0877_
rlabel metal3 69664 27720 69664 27720 0 _0878_
rlabel metal2 67032 27384 67032 27384 0 _0879_
rlabel metal2 70896 27832 70896 27832 0 _0880_
rlabel metal3 65968 26936 65968 26936 0 _0881_
rlabel metal2 74312 24192 74312 24192 0 _0882_
rlabel metal2 69720 22848 69720 22848 0 _0883_
rlabel metal2 66360 26964 66360 26964 0 _0884_
rlabel metal2 63448 27552 63448 27552 0 _0885_
rlabel metal2 62328 27440 62328 27440 0 _0886_
rlabel metal2 36568 35504 36568 35504 0 _0887_
rlabel metal2 33992 34776 33992 34776 0 _0888_
rlabel metal3 40544 32536 40544 32536 0 _0889_
rlabel metal2 39368 33432 39368 33432 0 _0890_
rlabel metal2 36120 32536 36120 32536 0 _0891_
rlabel metal2 42784 26264 42784 26264 0 _0892_
rlabel metal3 40040 27720 40040 27720 0 _0893_
rlabel metal2 38696 28560 38696 28560 0 _0894_
rlabel metal2 37688 30016 37688 30016 0 _0895_
rlabel metal2 36512 30408 36512 30408 0 _0896_
rlabel metal3 36288 29512 36288 29512 0 _0897_
rlabel metal2 38808 28224 38808 28224 0 _0898_
rlabel metal2 36120 28728 36120 28728 0 _0899_
rlabel metal2 37016 28952 37016 28952 0 _0900_
rlabel metal3 72408 27048 72408 27048 0 _0901_
rlabel metal2 73752 26320 73752 26320 0 _0902_
rlabel metal2 73192 26712 73192 26712 0 _0903_
rlabel metal3 42000 27832 42000 27832 0 _0904_
rlabel metal2 40936 28784 40936 28784 0 _0905_
rlabel metal3 71176 25256 71176 25256 0 _0906_
rlabel metal3 70840 27832 70840 27832 0 _0907_
rlabel metal2 72352 24024 72352 24024 0 _0908_
rlabel metal3 66808 27608 66808 27608 0 _0909_
rlabel metal2 62944 27048 62944 27048 0 _0910_
rlabel metal2 42392 28784 42392 28784 0 _0911_
rlabel metal2 39816 28672 39816 28672 0 _0912_
rlabel metal2 39368 29008 39368 29008 0 _0913_
rlabel metal2 38136 30576 38136 30576 0 _0914_
rlabel metal2 39480 30240 39480 30240 0 _0915_
rlabel metal2 38696 30464 38696 30464 0 _0916_
rlabel metal3 40768 29624 40768 29624 0 _0917_
rlabel metal2 71400 21112 71400 21112 0 _0918_
rlabel metal2 75096 21448 75096 21448 0 _0919_
rlabel metal3 72184 20664 72184 20664 0 _0920_
rlabel metal2 40264 28168 40264 28168 0 _0921_
rlabel metal2 38584 27328 38584 27328 0 _0922_
rlabel metal2 43064 24192 43064 24192 0 _0923_
rlabel metal2 68488 22568 68488 22568 0 _0924_
rlabel metal3 70672 21784 70672 21784 0 _0925_
rlabel metal2 69048 22400 69048 22400 0 _0926_
rlabel metal2 68376 22848 68376 22848 0 _0927_
rlabel metal2 63000 23632 63000 23632 0 _0928_
rlabel metal2 43288 24416 43288 24416 0 _0929_
rlabel metal2 37912 24584 37912 24584 0 _0930_
rlabel metal2 39368 27272 39368 27272 0 _0931_
rlabel metal3 39648 26936 39648 26936 0 _0932_
rlabel metal2 38024 26208 38024 26208 0 _0933_
rlabel metal2 38472 26544 38472 26544 0 _0934_
rlabel metal2 38696 27104 38696 27104 0 _0935_
rlabel metal2 38808 26600 38808 26600 0 _0936_
rlabel metal3 42448 23800 42448 23800 0 _0937_
rlabel metal3 39256 24808 39256 24808 0 _0938_
rlabel metal2 40264 25704 40264 25704 0 _0939_
rlabel metal2 40152 26376 40152 26376 0 _0940_
rlabel metal2 73976 18536 73976 18536 0 _0941_
rlabel metal2 73080 18088 73080 18088 0 _0942_
rlabel metal3 72128 17080 72128 17080 0 _0943_
rlabel metal3 38976 24696 38976 24696 0 _0944_
rlabel metal2 69720 19208 69720 19208 0 _0945_
rlabel metal2 69608 18872 69608 18872 0 _0946_
rlabel metal3 67592 18984 67592 18984 0 _0947_
rlabel metal3 66584 21784 66584 21784 0 _0948_
rlabel metal2 69720 20832 69720 20832 0 _0949_
rlabel metal2 65352 22064 65352 22064 0 _0950_
rlabel metal2 41944 21840 41944 21840 0 _0951_
rlabel metal3 41160 23352 41160 23352 0 _0952_
rlabel metal2 39256 23184 39256 23184 0 _0953_
rlabel metal2 39816 24304 39816 24304 0 _0954_
rlabel metal3 38248 23912 38248 23912 0 _0955_
rlabel metal2 41384 22344 41384 22344 0 _0956_
rlabel metal3 39592 21784 39592 21784 0 _0957_
rlabel metal2 40488 23240 40488 23240 0 _0958_
rlabel metal2 16296 25452 16296 25452 0 _0959_
rlabel metal2 26600 22400 26600 22400 0 _0960_
rlabel metal2 26488 21952 26488 21952 0 _0961_
rlabel metal2 18536 23968 18536 23968 0 _0962_
rlabel metal2 49280 21560 49280 21560 0 _0963_
rlabel metal2 15960 22736 15960 22736 0 _0964_
rlabel metal3 16912 23352 16912 23352 0 _0965_
rlabel metal2 19768 17304 19768 17304 0 _0966_
rlabel metal2 18536 4592 18536 4592 0 _0967_
rlabel metal2 43512 18872 43512 18872 0 _0968_
rlabel metal2 43680 15512 43680 15512 0 _0969_
rlabel metal2 41496 19600 41496 19600 0 _0970_
rlabel metal3 43176 16072 43176 16072 0 _0971_
rlabel metal2 44744 15568 44744 15568 0 _0972_
rlabel metal2 45192 15148 45192 15148 0 _0973_
rlabel metal3 19096 4312 19096 4312 0 _0974_
rlabel metal3 17136 4536 17136 4536 0 _0975_
rlabel metal2 25032 22176 25032 22176 0 _0976_
rlabel metal2 23800 21224 23800 21224 0 _0977_
rlabel metal2 23016 22512 23016 22512 0 _0978_
rlabel metal2 24248 21280 24248 21280 0 _0979_
rlabel metal2 24024 22064 24024 22064 0 _0980_
rlabel metal2 24304 7560 24304 7560 0 _0981_
rlabel metal2 24472 4536 24472 4536 0 _0982_
rlabel metal3 22568 4536 22568 4536 0 _0983_
rlabel metal2 47488 21560 47488 21560 0 _0984_
rlabel metal2 13272 11536 13272 11536 0 _0985_
rlabel metal2 26768 23128 26768 23128 0 _0986_
rlabel metal2 20328 22680 20328 22680 0 _0987_
rlabel metal2 17752 35224 17752 35224 0 _0988_
rlabel metal2 18536 22624 18536 22624 0 _0989_
rlabel metal3 46872 23352 46872 23352 0 _0990_
rlabel metal2 25704 23352 25704 23352 0 _0991_
rlabel metal3 18424 22064 18424 22064 0 _0992_
rlabel metal2 15176 15176 15176 15176 0 _0993_
rlabel metal3 6272 17528 6272 17528 0 _0994_
rlabel metal2 6944 27720 6944 27720 0 _0995_
rlabel metal3 4704 12936 4704 12936 0 _0996_
rlabel metal2 15456 34104 15456 34104 0 _0997_
rlabel metal2 15512 31864 15512 31864 0 _0998_
rlabel metal2 15680 23352 15680 23352 0 _0999_
rlabel metal3 15512 25536 15512 25536 0 _1000_
rlabel metal2 4984 28728 4984 28728 0 _1001_
rlabel metal2 5880 28336 5880 28336 0 _1002_
rlabel metal2 20328 8120 20328 8120 0 _1003_
rlabel metal2 26824 34608 26824 34608 0 _1004_
rlabel metal2 25760 33096 25760 33096 0 _1005_
rlabel metal3 23632 23016 23632 23016 0 _1006_
rlabel metal2 19880 8904 19880 8904 0 _1007_
rlabel metal2 7560 10248 7560 10248 0 _1008_
rlabel metal2 3192 11480 3192 11480 0 _1009_
rlabel metal2 23464 34272 23464 34272 0 _1010_
rlabel metal2 20832 33208 20832 33208 0 _1011_
rlabel metal2 22288 22568 22288 22568 0 _1012_
rlabel metal2 15400 23912 15400 23912 0 _1013_
rlabel metal2 10584 28728 10584 28728 0 _1014_
rlabel metal2 8344 28728 8344 28728 0 _1015_
rlabel metal2 44408 35168 44408 35168 0 _1016_
rlabel metal2 45360 31976 45360 31976 0 _1017_
rlabel metal2 44296 25872 44296 25872 0 _1018_
rlabel metal2 31136 22456 31136 22456 0 _1019_
rlabel metal2 32256 15288 32256 15288 0 _1020_
rlabel metal2 38136 6552 38136 6552 0 _1021_
rlabel metal2 38808 7952 38808 7952 0 _1022_
rlabel metal2 35672 8176 35672 8176 0 _1023_
rlabel metal2 47656 34944 47656 34944 0 _1024_
rlabel metal2 46648 29904 46648 29904 0 _1025_
rlabel metal2 44744 22008 44744 22008 0 _1026_
rlabel metal2 44632 8120 44632 8120 0 _1027_
rlabel metal2 49896 5488 49896 5488 0 _1028_
rlabel metal3 43848 5096 43848 5096 0 _1029_
rlabel metal2 48776 20328 48776 20328 0 _1030_
rlabel metal2 49112 20440 49112 20440 0 _1031_
rlabel metal2 49280 33992 49280 33992 0 _1032_
rlabel metal3 48328 33544 48328 33544 0 _1033_
rlabel metal2 50120 26264 50120 26264 0 _1034_
rlabel metal2 47768 25312 47768 25312 0 _1035_
rlabel metal2 48104 22400 48104 22400 0 _1036_
rlabel metal2 47880 21112 47880 21112 0 _1037_
rlabel metal2 55160 10304 55160 10304 0 _1038_
rlabel metal2 57288 5544 57288 5544 0 _1039_
rlabel metal3 54040 6552 54040 6552 0 _1040_
rlabel metal3 48440 30184 48440 30184 0 _1041_
rlabel metal2 45304 21448 45304 21448 0 _1042_
rlabel metal2 45192 21224 45192 21224 0 _1043_
rlabel metal3 64792 10472 64792 10472 0 _1044_
rlabel metal3 72408 3528 72408 3528 0 clk
rlabel metal3 2086 38360 2086 38360 0 dmem_addr[0]
rlabel metal3 1358 13720 1358 13720 0 dmem_addr[10]
rlabel metal3 1358 11256 1358 11256 0 dmem_addr[11]
rlabel metal3 1358 8792 1358 8792 0 dmem_addr[12]
rlabel metal3 1638 6328 1638 6328 0 dmem_addr[13]
rlabel metal3 1358 3864 1358 3864 0 dmem_addr[14]
rlabel metal3 1358 1400 1358 1400 0 dmem_addr[15]
rlabel metal3 1358 35896 1358 35896 0 dmem_addr[1]
rlabel metal3 1358 33432 1358 33432 0 dmem_addr[2]
rlabel metal3 1358 30968 1358 30968 0 dmem_addr[3]
rlabel metal3 1358 28504 1358 28504 0 dmem_addr[4]
rlabel metal2 1960 25872 1960 25872 0 dmem_addr[5]
rlabel metal3 1358 23576 1358 23576 0 dmem_addr[6]
rlabel metal3 1750 21112 1750 21112 0 dmem_addr[7]
rlabel metal3 1358 18648 1358 18648 0 dmem_addr[8]
rlabel metal3 1358 16184 1358 16184 0 dmem_addr[9]
rlabel metal3 77378 1400 77378 1400 0 dmem_data_in[0]
rlabel metal2 78008 26824 78008 26824 0 dmem_data_in[10]
rlabel metal2 75432 28616 75432 28616 0 dmem_data_in[11]
rlabel metal3 78610 30968 78610 30968 0 dmem_data_in[12]
rlabel metal2 78008 33656 78008 33656 0 dmem_data_in[13]
rlabel metal2 75096 35672 75096 35672 0 dmem_data_in[14]
rlabel metal3 76594 38360 76594 38360 0 dmem_data_in[15]
rlabel metal2 78008 3976 78008 3976 0 dmem_data_in[1]
rlabel metal2 78008 5936 78008 5936 0 dmem_data_in[2]
rlabel metal3 78610 8792 78610 8792 0 dmem_data_in[3]
rlabel metal3 76930 11256 76930 11256 0 dmem_data_in[4]
rlabel metal3 78162 13720 78162 13720 0 dmem_data_in[5]
rlabel metal2 78008 15680 78008 15680 0 dmem_data_in[6]
rlabel metal2 75096 19208 75096 19208 0 dmem_data_in[7]
rlabel metal3 78610 21112 78610 21112 0 dmem_data_in[8]
rlabel metal2 75432 23856 75432 23856 0 dmem_data_in[9]
rlabel metal2 4312 728 4312 728 0 dmem_data_out[0]
rlabel metal2 44072 3416 44072 3416 0 dmem_data_out[10]
rlabel metal2 48104 3416 48104 3416 0 dmem_data_out[11]
rlabel metal2 52136 3416 52136 3416 0 dmem_data_out[12]
rlabel metal2 56168 3416 56168 3416 0 dmem_data_out[13]
rlabel metal2 60200 3416 60200 3416 0 dmem_data_out[14]
rlabel metal2 64232 3416 64232 3416 0 dmem_data_out[15]
rlabel metal2 7784 3416 7784 3416 0 dmem_data_out[1]
rlabel metal2 11816 3416 11816 3416 0 dmem_data_out[2]
rlabel metal2 15848 3416 15848 3416 0 dmem_data_out[3]
rlabel metal3 20664 3528 20664 3528 0 dmem_data_out[4]
rlabel metal2 23968 2184 23968 2184 0 dmem_data_out[5]
rlabel metal2 28168 3416 28168 3416 0 dmem_data_out[6]
rlabel metal2 32032 3416 32032 3416 0 dmem_data_out[7]
rlabel metal2 35728 3416 35728 3416 0 dmem_data_out[8]
rlabel metal2 40096 2296 40096 2296 0 dmem_data_out[9]
rlabel metal2 68152 1414 68152 1414 0 dmem_we
rlabel metal2 38696 36512 38696 36512 0 instr[0]
rlabel metal2 13944 37898 13944 37898 0 instr[10]
rlabel metal2 11480 37898 11480 37898 0 instr[11]
rlabel metal2 8960 36568 8960 36568 0 instr[12]
rlabel metal2 6552 37898 6552 37898 0 instr[13]
rlabel metal2 4368 35896 4368 35896 0 instr[14]
rlabel metal2 1848 35056 1848 35056 0 instr[15]
rlabel metal2 35560 37912 35560 37912 0 instr[1]
rlabel metal2 33880 36848 33880 36848 0 instr[2]
rlabel metal2 31640 36904 31640 36904 0 instr[3]
rlabel metal2 29176 36848 29176 36848 0 instr[4]
rlabel metal2 24808 36176 24808 36176 0 instr[5]
rlabel metal2 23744 36568 23744 36568 0 instr[6]
rlabel metal2 21336 37898 21336 37898 0 instr[7]
rlabel metal2 18872 37898 18872 37898 0 instr[8]
rlabel metal2 16408 37898 16408 37898 0 instr[9]
rlabel metal3 71624 5432 71624 5432 0 net1
rlabel metal2 12264 3696 12264 3696 0 net10
rlabel metal2 13832 35952 13832 35952 0 net100
rlabel metal2 9464 31472 9464 31472 0 net101
rlabel metal2 20664 5824 20664 5824 0 net102
rlabel metal2 22008 7896 22008 7896 0 net103
rlabel metal3 25592 6104 25592 6104 0 net104
rlabel metal2 29736 9408 29736 9408 0 net105
rlabel metal2 37352 7952 37352 7952 0 net106
rlabel metal2 38696 8708 38696 8708 0 net107
rlabel metal3 26628 5880 26628 5880 0 net108
rlabel metal2 26320 11704 26320 11704 0 net109
rlabel metal2 15512 22568 15512 22568 0 net11
rlabel metal2 36232 6328 36232 6328 0 net110
rlabel via2 39032 5880 39032 5880 0 net111
rlabel metal2 47096 9744 47096 9744 0 net112
rlabel metal2 45416 16772 45416 16772 0 net113
rlabel metal2 47880 5488 47880 5488 0 net114
rlabel metal2 56056 4368 56056 4368 0 net115
rlabel metal3 50120 16912 50120 16912 0 net116
rlabel metal2 44296 5712 44296 5712 0 net117
rlabel metal2 49224 34776 49224 34776 0 net118
rlabel metal2 54376 34944 54376 34944 0 net119
rlabel metal2 20832 3416 20832 3416 0 net12
rlabel metal2 55384 7168 55384 7168 0 net120
rlabel metal2 61096 9856 61096 9856 0 net121
rlabel metal2 65128 10192 65128 10192 0 net122
rlabel metal2 65128 5152 65128 5152 0 net123
rlabel metal2 60648 17864 60648 17864 0 net124
rlabel metal2 70728 9016 70728 9016 0 net125
rlabel metal2 77896 17640 77896 17640 0 net126
rlabel metal2 73976 16856 73976 16856 0 net127
rlabel metal2 72632 10640 72632 10640 0 net128
rlabel metal3 65688 5880 65688 5880 0 net129
rlabel metal2 23184 4984 23184 4984 0 net13
rlabel metal2 60760 33320 60760 33320 0 net130
rlabel metal2 64680 30576 64680 30576 0 net131
rlabel metal2 63896 22064 63896 22064 0 net132
rlabel metal2 64904 31752 64904 31752 0 net133
rlabel metal2 70168 34384 70168 34384 0 net134
rlabel metal2 74872 30184 74872 30184 0 net135
rlabel metal2 75096 24696 75096 24696 0 net136
rlabel metal2 69832 31472 69832 31472 0 net137
rlabel metal2 69832 32172 69832 32172 0 net138
rlabel metal2 71288 7448 71288 7448 0 net139
rlabel metal2 30856 9240 30856 9240 0 net14
rlabel metal2 69776 7560 69776 7560 0 net140
rlabel metal2 48776 6664 48776 6664 0 net141
rlabel metal2 45080 22512 45080 22512 0 net15
rlabel metal2 47656 19376 47656 19376 0 net16
rlabel metal2 45136 20552 45136 20552 0 net17
rlabel metal2 39256 35896 39256 35896 0 net18
rlabel metal2 14504 36960 14504 36960 0 net19
rlabel metal3 15596 23240 15596 23240 0 net2
rlabel metal2 12264 35840 12264 35840 0 net20
rlabel metal2 9912 35672 9912 35672 0 net21
rlabel metal2 25256 24136 25256 24136 0 net22
rlabel metal2 5208 33320 5208 33320 0 net23
rlabel metal2 2408 29120 2408 29120 0 net24
rlabel metal2 36120 23744 36120 23744 0 net25
rlabel metal2 36568 22568 36568 22568 0 net26
rlabel metal2 44968 29568 44968 29568 0 net27
rlabel metal3 48384 28056 48384 28056 0 net28
rlabel metal2 27608 32816 27608 32816 0 net29
rlabel metal2 47432 5600 47432 5600 0 net3
rlabel metal2 25144 34664 25144 34664 0 net30
rlabel metal2 22120 36736 22120 36736 0 net31
rlabel metal2 19656 36624 19656 36624 0 net32
rlabel metal2 17304 36064 17304 36064 0 net33
rlabel metal2 73976 30128 73976 30128 0 net34
rlabel metal2 4760 33992 4760 33992 0 net35
rlabel metal2 49896 32928 49896 32928 0 net36
rlabel metal2 49952 20776 49952 20776 0 net37
rlabel metal2 34944 21784 34944 21784 0 net38
rlabel metal2 38920 9968 38920 9968 0 net39
rlabel metal2 51128 21560 51128 21560 0 net4
rlabel metal2 39088 20664 39088 20664 0 net40
rlabel metal2 41664 20664 41664 20664 0 net41
rlabel metal3 3472 35112 3472 35112 0 net42
rlabel metal2 4312 34048 4312 34048 0 net43
rlabel metal3 14616 31752 14616 31752 0 net44
rlabel metal2 4312 27888 4312 27888 0 net45
rlabel metal2 4312 25368 4312 25368 0 net46
rlabel metal2 42280 31248 42280 31248 0 net47
rlabel metal2 1848 21056 1848 21056 0 net48
rlabel metal2 4032 31192 4032 31192 0 net49
rlabel metal2 58632 22008 58632 22008 0 net5
rlabel metal2 3864 19208 3864 19208 0 net50
rlabel metal2 77224 5320 77224 5320 0 net51
rlabel metal2 75656 27160 75656 27160 0 net52
rlabel metal2 72744 29008 72744 29008 0 net53
rlabel metal2 75656 32816 75656 32816 0 net54
rlabel metal2 75544 34104 75544 34104 0 net55
rlabel metal2 73696 34440 73696 34440 0 net56
rlabel metal3 74760 33208 74760 33208 0 net57
rlabel metal2 75656 7336 75656 7336 0 net58
rlabel metal2 76104 6720 76104 6720 0 net59
rlabel metal2 57848 22400 57848 22400 0 net6
rlabel metal2 76104 9128 76104 9128 0 net60
rlabel metal2 76776 11312 76776 11312 0 net61
rlabel metal2 76888 14448 76888 14448 0 net62
rlabel metal2 76104 15400 76104 15400 0 net63
rlabel metal2 49448 18592 49448 18592 0 net64
rlabel metal2 75320 20384 75320 20384 0 net65
rlabel metal3 41608 24696 41608 24696 0 net66
rlabel metal2 40712 19096 40712 19096 0 net67
rlabel metal2 72744 32648 72744 32648 0 net68
rlabel metal2 54264 36008 54264 36008 0 net69
rlabel metal2 60648 20832 60648 20832 0 net7
rlabel metal3 54320 33320 54320 33320 0 net70
rlabel metal2 58856 34328 58856 34328 0 net71
rlabel metal2 63560 34496 63560 34496 0 net72
rlabel metal2 63672 32256 63672 32256 0 net73
rlabel metal3 44464 36456 44464 36456 0 net74
rlabel metal2 76328 34608 76328 34608 0 net75
rlabel metal2 74088 36680 74088 36680 0 net76
rlabel metal2 70840 36344 70840 36344 0 net77
rlabel metal2 68600 35140 68600 35140 0 net78
rlabel metal2 65912 35952 65912 35952 0 net79
rlabel metal3 63616 3640 63616 3640 0 net8
rlabel metal2 64456 35728 64456 35728 0 net80
rlabel metal2 48888 35560 48888 35560 0 net81
rlabel metal3 48608 35784 48608 35784 0 net82
rlabel metal2 49448 34272 49448 34272 0 net83
rlabel metal2 26600 35560 26600 35560 0 net84
rlabel metal2 18312 34160 18312 34160 0 net85
rlabel metal2 10080 6104 10080 6104 0 net86
rlabel metal2 2408 7448 2408 7448 0 net87
rlabel metal2 10360 7840 10360 7840 0 net88
rlabel metal2 2184 18424 2184 18424 0 net89
rlabel metal2 22400 21448 22400 21448 0 net9
rlabel metal3 6888 15960 6888 15960 0 net90
rlabel metal2 2744 7616 2744 7616 0 net91
rlabel metal2 16240 5992 16240 5992 0 net92
rlabel metal2 20048 6552 20048 6552 0 net93
rlabel metal2 15848 7196 15848 7196 0 net94
rlabel metal2 19992 5936 19992 5936 0 net95
rlabel metal2 1848 24696 1848 24696 0 net96
rlabel metal3 8456 27048 8456 27048 0 net97
rlabel metal2 2296 25088 2296 25088 0 net98
rlabel metal2 8568 30856 8568 30856 0 net99
rlabel metal2 75096 33264 75096 33264 0 pc[0]
rlabel metal2 53368 37954 53368 37954 0 pc[10]
rlabel metal2 50904 36610 50904 36610 0 pc[11]
rlabel metal2 48440 37170 48440 37170 0 pc[12]
rlabel metal2 47656 36792 47656 36792 0 pc[13]
rlabel metal2 43736 36680 43736 36680 0 pc[14]
rlabel metal2 41048 37898 41048 37898 0 pc[15]
rlabel metal2 75544 37562 75544 37562 0 pc[1]
rlabel metal2 73080 37954 73080 37954 0 pc[2]
rlabel metal2 71232 36680 71232 36680 0 pc[3]
rlabel metal3 68768 35112 68768 35112 0 pc[4]
rlabel metal2 67480 35784 67480 35784 0 pc[5]
rlabel metal2 63224 37562 63224 37562 0 pc[6]
rlabel metal3 61432 33544 61432 33544 0 pc[7]
rlabel metal2 64120 35896 64120 35896 0 pc[8]
rlabel metal2 55832 37226 55832 37226 0 pc[9]
rlabel metal2 18536 12768 18536 12768 0 register_file.reg_file_read\[1\]\[0\]
rlabel metal3 66080 19992 66080 19992 0 register_file.reg_file_read\[1\]\[10\]
rlabel metal2 45752 13328 45752 13328 0 register_file.reg_file_read\[1\]\[11\]
rlabel metal2 67704 34160 67704 34160 0 register_file.reg_file_read\[1\]\[12\]
rlabel metal2 73080 34664 73080 34664 0 register_file.reg_file_read\[1\]\[13\]
rlabel metal2 72520 21504 72520 21504 0 register_file.reg_file_read\[1\]\[14\]
rlabel metal3 71456 11256 71456 11256 0 register_file.reg_file_read\[1\]\[15\]
rlabel metal2 24416 5208 24416 5208 0 register_file.reg_file_read\[1\]\[1\]
rlabel metal3 17584 14280 17584 14280 0 register_file.reg_file_read\[1\]\[2\]
rlabel metal2 5992 27608 5992 27608 0 register_file.reg_file_read\[1\]\[3\]
rlabel metal2 21336 12488 21336 12488 0 register_file.reg_file_read\[1\]\[4\]
rlabel metal3 11088 27608 11088 27608 0 register_file.reg_file_read\[1\]\[5\]
rlabel metal3 35952 7336 35952 7336 0 register_file.reg_file_read\[1\]\[6\]
rlabel metal2 44296 13160 44296 13160 0 register_file.reg_file_read\[1\]\[7\]
rlabel metal3 57512 12824 57512 12824 0 register_file.reg_file_read\[1\]\[8\]
rlabel metal2 66584 12992 66584 12992 0 register_file.reg_file_read\[1\]\[9\]
rlabel metal3 13216 12824 13216 12824 0 register_file.reg_file_read\[2\]\[0\]
rlabel metal2 53928 17136 53928 17136 0 register_file.reg_file_read\[2\]\[10\]
rlabel metal2 49000 12656 49000 12656 0 register_file.reg_file_read\[2\]\[11\]
rlabel metal3 77840 25368 77840 25368 0 register_file.reg_file_read\[2\]\[12\]
rlabel metal2 75320 26208 75320 26208 0 register_file.reg_file_read\[2\]\[13\]
rlabel metal2 77000 22960 77000 22960 0 register_file.reg_file_read\[2\]\[14\]
rlabel metal2 74984 17192 74984 17192 0 register_file.reg_file_read\[2\]\[15\]
rlabel metal2 27720 11536 27720 11536 0 register_file.reg_file_read\[2\]\[1\]
rlabel metal2 11200 16856 11200 16856 0 register_file.reg_file_read\[2\]\[2\]
rlabel metal2 11256 20720 11256 20720 0 register_file.reg_file_read\[2\]\[3\]
rlabel metal3 21504 10696 21504 10696 0 register_file.reg_file_read\[2\]\[4\]
rlabel metal3 11592 21560 11592 21560 0 register_file.reg_file_read\[2\]\[5\]
rlabel metal2 32256 7560 32256 7560 0 register_file.reg_file_read\[2\]\[6\]
rlabel metal2 41272 11032 41272 11032 0 register_file.reg_file_read\[2\]\[7\]
rlabel metal2 57960 12208 57960 12208 0 register_file.reg_file_read\[2\]\[8\]
rlabel metal2 66920 13272 66920 13272 0 register_file.reg_file_read\[2\]\[9\]
rlabel metal2 16128 11256 16128 11256 0 register_file.reg_file_read\[3\]\[0\]
rlabel metal2 60984 17192 60984 17192 0 register_file.reg_file_read\[3\]\[10\]
rlabel metal2 48216 12656 48216 12656 0 register_file.reg_file_read\[3\]\[11\]
rlabel metal2 67704 32536 67704 32536 0 register_file.reg_file_read\[3\]\[12\]
rlabel metal3 73136 33432 73136 33432 0 register_file.reg_file_read\[3\]\[13\]
rlabel metal2 71736 21616 71736 21616 0 register_file.reg_file_read\[3\]\[14\]
rlabel metal2 72408 10080 72408 10080 0 register_file.reg_file_read\[3\]\[15\]
rlabel metal2 22792 4928 22792 4928 0 register_file.reg_file_read\[3\]\[1\]
rlabel metal2 16184 17696 16184 17696 0 register_file.reg_file_read\[3\]\[2\]
rlabel metal3 6440 29176 6440 29176 0 register_file.reg_file_read\[3\]\[3\]
rlabel metal2 20104 13552 20104 13552 0 register_file.reg_file_read\[3\]\[4\]
rlabel metal2 11368 28952 11368 28952 0 register_file.reg_file_read\[3\]\[5\]
rlabel metal2 35000 12992 35000 12992 0 register_file.reg_file_read\[3\]\[6\]
rlabel metal2 41216 12264 41216 12264 0 register_file.reg_file_read\[3\]\[7\]
rlabel metal3 59640 12264 59640 12264 0 register_file.reg_file_read\[3\]\[8\]
rlabel metal2 66360 4648 66360 4648 0 register_file.reg_file_read\[3\]\[9\]
rlabel metal2 16352 9912 16352 9912 0 register_file.reg_file_read\[4\]\[0\]
rlabel via2 55832 18312 55832 18312 0 register_file.reg_file_read\[4\]\[10\]
rlabel metal2 43064 12040 43064 12040 0 register_file.reg_file_read\[4\]\[11\]
rlabel metal2 68712 27384 68712 27384 0 register_file.reg_file_read\[4\]\[12\]
rlabel metal2 75320 30464 75320 30464 0 register_file.reg_file_read\[4\]\[13\]
rlabel metal2 77224 22624 77224 22624 0 register_file.reg_file_read\[4\]\[14\]
rlabel metal2 75320 18368 75320 18368 0 register_file.reg_file_read\[4\]\[15\]
rlabel metal2 24472 15792 24472 15792 0 register_file.reg_file_read\[4\]\[1\]
rlabel metal2 15736 16408 15736 16408 0 register_file.reg_file_read\[4\]\[2\]
rlabel metal2 16744 20384 16744 20384 0 register_file.reg_file_read\[4\]\[3\]
rlabel metal2 21448 9968 21448 9968 0 register_file.reg_file_read\[4\]\[4\]
rlabel metal2 21896 20328 21896 20328 0 register_file.reg_file_read\[4\]\[5\]
rlabel metal2 31976 11704 31976 11704 0 register_file.reg_file_read\[4\]\[6\]
rlabel metal3 39704 10696 39704 10696 0 register_file.reg_file_read\[4\]\[7\]
rlabel metal2 60424 11312 60424 11312 0 register_file.reg_file_read\[4\]\[8\]
rlabel metal2 66248 13048 66248 13048 0 register_file.reg_file_read\[4\]\[9\]
rlabel metal3 13440 5208 13440 5208 0 register_file.reg_file_read\[5\]\[0\]
rlabel metal2 56840 18984 56840 18984 0 register_file.reg_file_read\[5\]\[10\]
rlabel metal3 45640 9016 45640 9016 0 register_file.reg_file_read\[5\]\[11\]
rlabel metal3 69552 29960 69552 29960 0 register_file.reg_file_read\[5\]\[12\]
rlabel metal2 71176 27776 71176 27776 0 register_file.reg_file_read\[5\]\[13\]
rlabel metal2 74872 22176 74872 22176 0 register_file.reg_file_read\[5\]\[14\]
rlabel metal2 69552 17752 69552 17752 0 register_file.reg_file_read\[5\]\[15\]
rlabel metal2 28168 6272 28168 6272 0 register_file.reg_file_read\[5\]\[1\]
rlabel metal2 11872 16856 11872 16856 0 register_file.reg_file_read\[5\]\[2\]
rlabel metal2 4088 25424 4088 25424 0 register_file.reg_file_read\[5\]\[3\]
rlabel metal2 23576 11144 23576 11144 0 register_file.reg_file_read\[5\]\[4\]
rlabel metal3 8848 26264 8848 26264 0 register_file.reg_file_read\[5\]\[5\]
rlabel metal2 31696 12824 31696 12824 0 register_file.reg_file_read\[5\]\[6\]
rlabel metal3 46200 6888 46200 6888 0 register_file.reg_file_read\[5\]\[7\]
rlabel metal2 61320 14056 61320 14056 0 register_file.reg_file_read\[5\]\[8\]
rlabel metal2 64400 13720 64400 13720 0 register_file.reg_file_read\[5\]\[9\]
rlabel metal2 11928 4928 11928 4928 0 register_file.reg_file_read\[6\]\[0\]
rlabel metal2 63448 17640 63448 17640 0 register_file.reg_file_read\[6\]\[10\]
rlabel metal2 44128 11368 44128 11368 0 register_file.reg_file_read\[6\]\[11\]
rlabel metal2 67592 30520 67592 30520 0 register_file.reg_file_read\[6\]\[12\]
rlabel metal2 72072 28672 72072 28672 0 register_file.reg_file_read\[6\]\[13\]
rlabel metal2 68936 14504 68936 14504 0 register_file.reg_file_read\[6\]\[14\]
rlabel metal3 67424 21672 67424 21672 0 register_file.reg_file_read\[6\]\[15\]
rlabel metal2 28448 11368 28448 11368 0 register_file.reg_file_read\[6\]\[1\]
rlabel metal2 10360 16520 10360 16520 0 register_file.reg_file_read\[6\]\[2\]
rlabel metal3 10248 20776 10248 20776 0 register_file.reg_file_read\[6\]\[3\]
rlabel metal2 19880 10584 19880 10584 0 register_file.reg_file_read\[6\]\[4\]
rlabel metal3 10136 21560 10136 21560 0 register_file.reg_file_read\[6\]\[5\]
rlabel metal3 32368 12264 32368 12264 0 register_file.reg_file_read\[6\]\[6\]
rlabel metal2 49224 4592 49224 4592 0 register_file.reg_file_read\[6\]\[7\]
rlabel metal2 56728 13328 56728 13328 0 register_file.reg_file_read\[6\]\[8\]
rlabel metal2 64008 14448 64008 14448 0 register_file.reg_file_read\[6\]\[9\]
rlabel metal2 17752 12936 17752 12936 0 register_file.reg_file_read\[7\]\[0\]
rlabel metal2 58968 18144 58968 18144 0 register_file.reg_file_read\[7\]\[10\]
rlabel metal2 47936 17640 47936 17640 0 register_file.reg_file_read\[7\]\[11\]
rlabel metal3 67872 25480 67872 25480 0 register_file.reg_file_read\[7\]\[12\]
rlabel metal2 68936 23240 68936 23240 0 register_file.reg_file_read\[7\]\[13\]
rlabel metal3 69944 23128 69944 23128 0 register_file.reg_file_read\[7\]\[14\]
rlabel metal2 71736 18424 71736 18424 0 register_file.reg_file_read\[7\]\[15\]
rlabel metal2 24024 12936 24024 12936 0 register_file.reg_file_read\[7\]\[1\]
rlabel metal2 16744 14616 16744 14616 0 register_file.reg_file_read\[7\]\[2\]
rlabel metal3 12488 25704 12488 25704 0 register_file.reg_file_read\[7\]\[3\]
rlabel metal2 20440 10528 20440 10528 0 register_file.reg_file_read\[7\]\[4\]
rlabel metal2 18312 21168 18312 21168 0 register_file.reg_file_read\[7\]\[5\]
rlabel metal2 35448 13384 35448 13384 0 register_file.reg_file_read\[7\]\[6\]
rlabel metal2 42392 11592 42392 11592 0 register_file.reg_file_read\[7\]\[7\]
rlabel metal2 59416 12936 59416 12936 0 register_file.reg_file_read\[7\]\[8\]
rlabel metal2 64008 9464 64008 9464 0 register_file.reg_file_read\[7\]\[9\]
rlabel metal2 76216 2058 76216 2058 0 rst_n
<< properties >>
string FIXED_BBOX 0 0 80000 40000
<< end >>
