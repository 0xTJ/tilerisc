magic
tech gf180mcuD
magscale 1 5
timestamp 1702129541
<< obsm1 >>
rect 672 1538 149296 148206
<< metal2 >>
rect 2576 0 2632 400
rect 6832 0 6888 400
rect 11088 0 11144 400
rect 15344 0 15400 400
rect 19600 0 19656 400
rect 23856 0 23912 400
rect 28112 0 28168 400
rect 32368 0 32424 400
rect 36624 0 36680 400
rect 40880 0 40936 400
rect 45136 0 45192 400
rect 49392 0 49448 400
rect 53648 0 53704 400
rect 57904 0 57960 400
rect 62160 0 62216 400
rect 66416 0 66472 400
rect 70672 0 70728 400
rect 74928 0 74984 400
rect 79184 0 79240 400
rect 83440 0 83496 400
rect 87696 0 87752 400
rect 91952 0 92008 400
rect 96208 0 96264 400
rect 100464 0 100520 400
rect 104720 0 104776 400
rect 108976 0 109032 400
rect 113232 0 113288 400
rect 117488 0 117544 400
rect 121744 0 121800 400
rect 126000 0 126056 400
rect 130256 0 130312 400
rect 134512 0 134568 400
rect 138768 0 138824 400
rect 143024 0 143080 400
rect 147280 0 147336 400
<< obsm2 >>
rect 910 430 149170 148195
rect 910 350 2546 430
rect 2662 350 6802 430
rect 6918 350 11058 430
rect 11174 350 15314 430
rect 15430 350 19570 430
rect 19686 350 23826 430
rect 23942 350 28082 430
rect 28198 350 32338 430
rect 32454 350 36594 430
rect 36710 350 40850 430
rect 40966 350 45106 430
rect 45222 350 49362 430
rect 49478 350 53618 430
rect 53734 350 57874 430
rect 57990 350 62130 430
rect 62246 350 66386 430
rect 66502 350 70642 430
rect 70758 350 74898 430
rect 75014 350 79154 430
rect 79270 350 83410 430
rect 83526 350 87666 430
rect 87782 350 91922 430
rect 92038 350 96178 430
rect 96294 350 100434 430
rect 100550 350 104690 430
rect 104806 350 108946 430
rect 109062 350 113202 430
rect 113318 350 117458 430
rect 117574 350 121714 430
rect 121830 350 125970 430
rect 126086 350 130226 430
rect 130342 350 134482 430
rect 134598 350 138738 430
rect 138854 350 142994 430
rect 143110 350 147250 430
rect 147366 350 149170 430
<< metal3 >>
rect 0 145488 400 145544
rect 149600 145488 150000 145544
rect 0 143248 400 143304
rect 149600 143248 150000 143304
rect 0 141008 400 141064
rect 149600 141008 150000 141064
rect 0 138768 400 138824
rect 149600 138768 150000 138824
rect 0 136528 400 136584
rect 149600 136528 150000 136584
rect 0 134288 400 134344
rect 149600 134288 150000 134344
rect 0 132048 400 132104
rect 149600 132048 150000 132104
rect 0 129808 400 129864
rect 149600 129808 150000 129864
rect 0 127568 400 127624
rect 149600 127568 150000 127624
rect 0 125328 400 125384
rect 149600 125328 150000 125384
rect 0 123088 400 123144
rect 149600 123088 150000 123144
rect 0 120848 400 120904
rect 149600 120848 150000 120904
rect 0 118608 400 118664
rect 149600 118608 150000 118664
rect 0 116368 400 116424
rect 149600 116368 150000 116424
rect 0 114128 400 114184
rect 149600 114128 150000 114184
rect 0 111888 400 111944
rect 149600 111888 150000 111944
rect 0 109648 400 109704
rect 149600 109648 150000 109704
rect 0 107408 400 107464
rect 149600 107408 150000 107464
rect 0 105168 400 105224
rect 149600 105168 150000 105224
rect 0 102928 400 102984
rect 149600 102928 150000 102984
rect 0 100688 400 100744
rect 149600 100688 150000 100744
rect 0 98448 400 98504
rect 149600 98448 150000 98504
rect 0 96208 400 96264
rect 149600 96208 150000 96264
rect 0 93968 400 94024
rect 149600 93968 150000 94024
rect 0 91728 400 91784
rect 149600 91728 150000 91784
rect 0 89488 400 89544
rect 149600 89488 150000 89544
rect 0 87248 400 87304
rect 149600 87248 150000 87304
rect 0 85008 400 85064
rect 149600 85008 150000 85064
rect 0 82768 400 82824
rect 149600 82768 150000 82824
rect 0 80528 400 80584
rect 149600 80528 150000 80584
rect 0 78288 400 78344
rect 149600 78288 150000 78344
rect 0 76048 400 76104
rect 149600 76048 150000 76104
rect 0 73808 400 73864
rect 149600 73808 150000 73864
rect 0 71568 400 71624
rect 149600 71568 150000 71624
rect 0 69328 400 69384
rect 149600 69328 150000 69384
rect 0 67088 400 67144
rect 149600 67088 150000 67144
rect 0 64848 400 64904
rect 149600 64848 150000 64904
rect 0 62608 400 62664
rect 149600 62608 150000 62664
rect 0 60368 400 60424
rect 149600 60368 150000 60424
rect 0 58128 400 58184
rect 149600 58128 150000 58184
rect 0 55888 400 55944
rect 149600 55888 150000 55944
rect 0 53648 400 53704
rect 149600 53648 150000 53704
rect 0 51408 400 51464
rect 149600 51408 150000 51464
rect 0 49168 400 49224
rect 149600 49168 150000 49224
rect 0 46928 400 46984
rect 149600 46928 150000 46984
rect 0 44688 400 44744
rect 149600 44688 150000 44744
rect 0 42448 400 42504
rect 149600 42448 150000 42504
rect 0 40208 400 40264
rect 149600 40208 150000 40264
rect 0 37968 400 38024
rect 149600 37968 150000 38024
rect 0 35728 400 35784
rect 149600 35728 150000 35784
rect 0 33488 400 33544
rect 149600 33488 150000 33544
rect 0 31248 400 31304
rect 149600 31248 150000 31304
rect 0 29008 400 29064
rect 149600 29008 150000 29064
rect 0 26768 400 26824
rect 149600 26768 150000 26824
rect 0 24528 400 24584
rect 149600 24528 150000 24584
rect 0 22288 400 22344
rect 149600 22288 150000 22344
rect 0 20048 400 20104
rect 149600 20048 150000 20104
rect 0 17808 400 17864
rect 149600 17808 150000 17864
rect 0 15568 400 15624
rect 149600 15568 150000 15624
rect 0 13328 400 13384
rect 149600 13328 150000 13384
rect 0 11088 400 11144
rect 149600 11088 150000 11144
rect 0 8848 400 8904
rect 149600 8848 150000 8904
rect 0 6608 400 6664
rect 149600 6608 150000 6664
rect 0 4368 400 4424
rect 149600 4368 150000 4424
<< obsm3 >>
rect 400 145574 149600 148190
rect 430 145458 149570 145574
rect 400 143334 149600 145458
rect 430 143218 149570 143334
rect 400 141094 149600 143218
rect 430 140978 149570 141094
rect 400 138854 149600 140978
rect 430 138738 149570 138854
rect 400 136614 149600 138738
rect 430 136498 149570 136614
rect 400 134374 149600 136498
rect 430 134258 149570 134374
rect 400 132134 149600 134258
rect 430 132018 149570 132134
rect 400 129894 149600 132018
rect 430 129778 149570 129894
rect 400 127654 149600 129778
rect 430 127538 149570 127654
rect 400 125414 149600 127538
rect 430 125298 149570 125414
rect 400 123174 149600 125298
rect 430 123058 149570 123174
rect 400 120934 149600 123058
rect 430 120818 149570 120934
rect 400 118694 149600 120818
rect 430 118578 149570 118694
rect 400 116454 149600 118578
rect 430 116338 149570 116454
rect 400 114214 149600 116338
rect 430 114098 149570 114214
rect 400 111974 149600 114098
rect 430 111858 149570 111974
rect 400 109734 149600 111858
rect 430 109618 149570 109734
rect 400 107494 149600 109618
rect 430 107378 149570 107494
rect 400 105254 149600 107378
rect 430 105138 149570 105254
rect 400 103014 149600 105138
rect 430 102898 149570 103014
rect 400 100774 149600 102898
rect 430 100658 149570 100774
rect 400 98534 149600 100658
rect 430 98418 149570 98534
rect 400 96294 149600 98418
rect 430 96178 149570 96294
rect 400 94054 149600 96178
rect 430 93938 149570 94054
rect 400 91814 149600 93938
rect 430 91698 149570 91814
rect 400 89574 149600 91698
rect 430 89458 149570 89574
rect 400 87334 149600 89458
rect 430 87218 149570 87334
rect 400 85094 149600 87218
rect 430 84978 149570 85094
rect 400 82854 149600 84978
rect 430 82738 149570 82854
rect 400 80614 149600 82738
rect 430 80498 149570 80614
rect 400 78374 149600 80498
rect 430 78258 149570 78374
rect 400 76134 149600 78258
rect 430 76018 149570 76134
rect 400 73894 149600 76018
rect 430 73778 149570 73894
rect 400 71654 149600 73778
rect 430 71538 149570 71654
rect 400 69414 149600 71538
rect 430 69298 149570 69414
rect 400 67174 149600 69298
rect 430 67058 149570 67174
rect 400 64934 149600 67058
rect 430 64818 149570 64934
rect 400 62694 149600 64818
rect 430 62578 149570 62694
rect 400 60454 149600 62578
rect 430 60338 149570 60454
rect 400 58214 149600 60338
rect 430 58098 149570 58214
rect 400 55974 149600 58098
rect 430 55858 149570 55974
rect 400 53734 149600 55858
rect 430 53618 149570 53734
rect 400 51494 149600 53618
rect 430 51378 149570 51494
rect 400 49254 149600 51378
rect 430 49138 149570 49254
rect 400 47014 149600 49138
rect 430 46898 149570 47014
rect 400 44774 149600 46898
rect 430 44658 149570 44774
rect 400 42534 149600 44658
rect 430 42418 149570 42534
rect 400 40294 149600 42418
rect 430 40178 149570 40294
rect 400 38054 149600 40178
rect 430 37938 149570 38054
rect 400 35814 149600 37938
rect 430 35698 149570 35814
rect 400 33574 149600 35698
rect 430 33458 149570 33574
rect 400 31334 149600 33458
rect 430 31218 149570 31334
rect 400 29094 149600 31218
rect 430 28978 149570 29094
rect 400 26854 149600 28978
rect 430 26738 149570 26854
rect 400 24614 149600 26738
rect 430 24498 149570 24614
rect 400 22374 149600 24498
rect 430 22258 149570 22374
rect 400 20134 149600 22258
rect 430 20018 149570 20134
rect 400 17894 149600 20018
rect 430 17778 149570 17894
rect 400 15654 149600 17778
rect 430 15538 149570 15654
rect 400 13414 149600 15538
rect 430 13298 149570 13414
rect 400 11174 149600 13298
rect 430 11058 149570 11174
rect 400 8934 149600 11058
rect 430 8818 149570 8934
rect 400 6694 149600 8818
rect 430 6578 149570 6694
rect 400 4454 149600 6578
rect 430 4338 149570 4454
rect 400 1554 149600 4338
<< metal4 >>
rect 2224 1538 2384 148206
rect 9904 1538 10064 148206
rect 17584 1538 17744 148206
rect 25264 1538 25424 148206
rect 32944 1538 33104 148206
rect 40624 1538 40784 148206
rect 48304 1538 48464 148206
rect 55984 1538 56144 148206
rect 63664 1538 63824 148206
rect 71344 1538 71504 148206
rect 79024 1538 79184 148206
rect 86704 1538 86864 148206
rect 94384 1538 94544 148206
rect 102064 1538 102224 148206
rect 109744 1538 109904 148206
rect 117424 1538 117584 148206
rect 125104 1538 125264 148206
rect 132784 1538 132944 148206
rect 140464 1538 140624 148206
rect 148144 1538 148304 148206
<< obsm4 >>
rect 6790 26833 9874 141223
rect 10094 26833 17554 141223
rect 17774 26833 25234 141223
rect 25454 26833 32914 141223
rect 33134 26833 40594 141223
rect 40814 26833 48274 141223
rect 48494 26833 55954 141223
rect 56174 26833 63634 141223
rect 63854 26833 71314 141223
rect 71534 26833 78994 141223
rect 79214 26833 86674 141223
rect 86894 26833 94354 141223
rect 94574 26833 102034 141223
rect 102254 26833 109714 141223
rect 109934 26833 117394 141223
rect 117614 26833 125074 141223
rect 125294 26833 132754 141223
rect 132974 26833 140434 141223
rect 140654 26833 140770 141223
<< labels >>
rlabel metal2 s 11088 0 11144 400 6 ack
port 1 nsew signal output
rlabel metal2 s 2576 0 2632 400 6 clk
port 2 nsew signal input
rlabel metal2 s 15344 0 15400 400 6 command[0]
port 3 nsew signal input
rlabel metal2 s 57904 0 57960 400 6 command[10]
port 4 nsew signal input
rlabel metal2 s 62160 0 62216 400 6 command[11]
port 5 nsew signal input
rlabel metal2 s 66416 0 66472 400 6 command[12]
port 6 nsew signal input
rlabel metal2 s 70672 0 70728 400 6 command[13]
port 7 nsew signal input
rlabel metal2 s 74928 0 74984 400 6 command[14]
port 8 nsew signal input
rlabel metal2 s 79184 0 79240 400 6 command[15]
port 9 nsew signal input
rlabel metal2 s 83440 0 83496 400 6 command[16]
port 10 nsew signal input
rlabel metal2 s 87696 0 87752 400 6 command[17]
port 11 nsew signal input
rlabel metal2 s 91952 0 92008 400 6 command[18]
port 12 nsew signal input
rlabel metal2 s 96208 0 96264 400 6 command[19]
port 13 nsew signal input
rlabel metal2 s 19600 0 19656 400 6 command[1]
port 14 nsew signal input
rlabel metal2 s 100464 0 100520 400 6 command[20]
port 15 nsew signal input
rlabel metal2 s 104720 0 104776 400 6 command[21]
port 16 nsew signal input
rlabel metal2 s 108976 0 109032 400 6 command[22]
port 17 nsew signal input
rlabel metal2 s 113232 0 113288 400 6 command[23]
port 18 nsew signal input
rlabel metal2 s 117488 0 117544 400 6 command[24]
port 19 nsew signal input
rlabel metal2 s 121744 0 121800 400 6 command[25]
port 20 nsew signal input
rlabel metal2 s 126000 0 126056 400 6 command[26]
port 21 nsew signal input
rlabel metal2 s 130256 0 130312 400 6 command[27]
port 22 nsew signal input
rlabel metal2 s 134512 0 134568 400 6 command[28]
port 23 nsew signal input
rlabel metal2 s 138768 0 138824 400 6 command[29]
port 24 nsew signal input
rlabel metal2 s 23856 0 23912 400 6 command[2]
port 25 nsew signal input
rlabel metal2 s 143024 0 143080 400 6 command[30]
port 26 nsew signal input
rlabel metal2 s 147280 0 147336 400 6 command[31]
port 27 nsew signal input
rlabel metal2 s 28112 0 28168 400 6 command[3]
port 28 nsew signal input
rlabel metal2 s 32368 0 32424 400 6 command[4]
port 29 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 command[5]
port 30 nsew signal input
rlabel metal2 s 40880 0 40936 400 6 command[6]
port 31 nsew signal input
rlabel metal2 s 45136 0 45192 400 6 command[7]
port 32 nsew signal input
rlabel metal2 s 49392 0 49448 400 6 command[8]
port 33 nsew signal input
rlabel metal2 s 53648 0 53704 400 6 command[9]
port 34 nsew signal input
rlabel metal3 s 149600 4368 150000 4424 6 data_in[0]
port 35 nsew signal input
rlabel metal3 s 149600 26768 150000 26824 6 data_in[10]
port 36 nsew signal input
rlabel metal3 s 149600 29008 150000 29064 6 data_in[11]
port 37 nsew signal input
rlabel metal3 s 149600 31248 150000 31304 6 data_in[12]
port 38 nsew signal input
rlabel metal3 s 149600 33488 150000 33544 6 data_in[13]
port 39 nsew signal input
rlabel metal3 s 149600 35728 150000 35784 6 data_in[14]
port 40 nsew signal input
rlabel metal3 s 149600 37968 150000 38024 6 data_in[15]
port 41 nsew signal input
rlabel metal3 s 149600 40208 150000 40264 6 data_in[16]
port 42 nsew signal input
rlabel metal3 s 149600 42448 150000 42504 6 data_in[17]
port 43 nsew signal input
rlabel metal3 s 149600 44688 150000 44744 6 data_in[18]
port 44 nsew signal input
rlabel metal3 s 149600 46928 150000 46984 6 data_in[19]
port 45 nsew signal input
rlabel metal3 s 149600 6608 150000 6664 6 data_in[1]
port 46 nsew signal input
rlabel metal3 s 149600 49168 150000 49224 6 data_in[20]
port 47 nsew signal input
rlabel metal3 s 149600 51408 150000 51464 6 data_in[21]
port 48 nsew signal input
rlabel metal3 s 149600 53648 150000 53704 6 data_in[22]
port 49 nsew signal input
rlabel metal3 s 149600 55888 150000 55944 6 data_in[23]
port 50 nsew signal input
rlabel metal3 s 149600 58128 150000 58184 6 data_in[24]
port 51 nsew signal input
rlabel metal3 s 149600 60368 150000 60424 6 data_in[25]
port 52 nsew signal input
rlabel metal3 s 149600 62608 150000 62664 6 data_in[26]
port 53 nsew signal input
rlabel metal3 s 149600 64848 150000 64904 6 data_in[27]
port 54 nsew signal input
rlabel metal3 s 149600 67088 150000 67144 6 data_in[28]
port 55 nsew signal input
rlabel metal3 s 149600 69328 150000 69384 6 data_in[29]
port 56 nsew signal input
rlabel metal3 s 149600 8848 150000 8904 6 data_in[2]
port 57 nsew signal input
rlabel metal3 s 149600 71568 150000 71624 6 data_in[30]
port 58 nsew signal input
rlabel metal3 s 149600 73808 150000 73864 6 data_in[31]
port 59 nsew signal input
rlabel metal3 s 149600 76048 150000 76104 6 data_in[32]
port 60 nsew signal input
rlabel metal3 s 149600 78288 150000 78344 6 data_in[33]
port 61 nsew signal input
rlabel metal3 s 149600 80528 150000 80584 6 data_in[34]
port 62 nsew signal input
rlabel metal3 s 149600 82768 150000 82824 6 data_in[35]
port 63 nsew signal input
rlabel metal3 s 149600 85008 150000 85064 6 data_in[36]
port 64 nsew signal input
rlabel metal3 s 149600 87248 150000 87304 6 data_in[37]
port 65 nsew signal input
rlabel metal3 s 149600 89488 150000 89544 6 data_in[38]
port 66 nsew signal input
rlabel metal3 s 149600 91728 150000 91784 6 data_in[39]
port 67 nsew signal input
rlabel metal3 s 149600 11088 150000 11144 6 data_in[3]
port 68 nsew signal input
rlabel metal3 s 149600 93968 150000 94024 6 data_in[40]
port 69 nsew signal input
rlabel metal3 s 149600 96208 150000 96264 6 data_in[41]
port 70 nsew signal input
rlabel metal3 s 149600 98448 150000 98504 6 data_in[42]
port 71 nsew signal input
rlabel metal3 s 149600 100688 150000 100744 6 data_in[43]
port 72 nsew signal input
rlabel metal3 s 149600 102928 150000 102984 6 data_in[44]
port 73 nsew signal input
rlabel metal3 s 149600 105168 150000 105224 6 data_in[45]
port 74 nsew signal input
rlabel metal3 s 149600 107408 150000 107464 6 data_in[46]
port 75 nsew signal input
rlabel metal3 s 149600 109648 150000 109704 6 data_in[47]
port 76 nsew signal input
rlabel metal3 s 149600 111888 150000 111944 6 data_in[48]
port 77 nsew signal input
rlabel metal3 s 149600 114128 150000 114184 6 data_in[49]
port 78 nsew signal input
rlabel metal3 s 149600 13328 150000 13384 6 data_in[4]
port 79 nsew signal input
rlabel metal3 s 149600 116368 150000 116424 6 data_in[50]
port 80 nsew signal input
rlabel metal3 s 149600 118608 150000 118664 6 data_in[51]
port 81 nsew signal input
rlabel metal3 s 149600 120848 150000 120904 6 data_in[52]
port 82 nsew signal input
rlabel metal3 s 149600 123088 150000 123144 6 data_in[53]
port 83 nsew signal input
rlabel metal3 s 149600 125328 150000 125384 6 data_in[54]
port 84 nsew signal input
rlabel metal3 s 149600 127568 150000 127624 6 data_in[55]
port 85 nsew signal input
rlabel metal3 s 149600 129808 150000 129864 6 data_in[56]
port 86 nsew signal input
rlabel metal3 s 149600 132048 150000 132104 6 data_in[57]
port 87 nsew signal input
rlabel metal3 s 149600 134288 150000 134344 6 data_in[58]
port 88 nsew signal input
rlabel metal3 s 149600 136528 150000 136584 6 data_in[59]
port 89 nsew signal input
rlabel metal3 s 149600 15568 150000 15624 6 data_in[5]
port 90 nsew signal input
rlabel metal3 s 149600 138768 150000 138824 6 data_in[60]
port 91 nsew signal input
rlabel metal3 s 149600 141008 150000 141064 6 data_in[61]
port 92 nsew signal input
rlabel metal3 s 149600 143248 150000 143304 6 data_in[62]
port 93 nsew signal input
rlabel metal3 s 149600 145488 150000 145544 6 data_in[63]
port 94 nsew signal input
rlabel metal3 s 149600 17808 150000 17864 6 data_in[6]
port 95 nsew signal input
rlabel metal3 s 149600 20048 150000 20104 6 data_in[7]
port 96 nsew signal input
rlabel metal3 s 149600 22288 150000 22344 6 data_in[8]
port 97 nsew signal input
rlabel metal3 s 149600 24528 150000 24584 6 data_in[9]
port 98 nsew signal input
rlabel metal3 s 0 145488 400 145544 6 data_out[0]
port 99 nsew signal output
rlabel metal3 s 0 123088 400 123144 6 data_out[10]
port 100 nsew signal output
rlabel metal3 s 0 120848 400 120904 6 data_out[11]
port 101 nsew signal output
rlabel metal3 s 0 118608 400 118664 6 data_out[12]
port 102 nsew signal output
rlabel metal3 s 0 116368 400 116424 6 data_out[13]
port 103 nsew signal output
rlabel metal3 s 0 114128 400 114184 6 data_out[14]
port 104 nsew signal output
rlabel metal3 s 0 111888 400 111944 6 data_out[15]
port 105 nsew signal output
rlabel metal3 s 0 109648 400 109704 6 data_out[16]
port 106 nsew signal output
rlabel metal3 s 0 107408 400 107464 6 data_out[17]
port 107 nsew signal output
rlabel metal3 s 0 105168 400 105224 6 data_out[18]
port 108 nsew signal output
rlabel metal3 s 0 102928 400 102984 6 data_out[19]
port 109 nsew signal output
rlabel metal3 s 0 143248 400 143304 6 data_out[1]
port 110 nsew signal output
rlabel metal3 s 0 100688 400 100744 6 data_out[20]
port 111 nsew signal output
rlabel metal3 s 0 98448 400 98504 6 data_out[21]
port 112 nsew signal output
rlabel metal3 s 0 96208 400 96264 6 data_out[22]
port 113 nsew signal output
rlabel metal3 s 0 93968 400 94024 6 data_out[23]
port 114 nsew signal output
rlabel metal3 s 0 91728 400 91784 6 data_out[24]
port 115 nsew signal output
rlabel metal3 s 0 89488 400 89544 6 data_out[25]
port 116 nsew signal output
rlabel metal3 s 0 87248 400 87304 6 data_out[26]
port 117 nsew signal output
rlabel metal3 s 0 85008 400 85064 6 data_out[27]
port 118 nsew signal output
rlabel metal3 s 0 82768 400 82824 6 data_out[28]
port 119 nsew signal output
rlabel metal3 s 0 80528 400 80584 6 data_out[29]
port 120 nsew signal output
rlabel metal3 s 0 141008 400 141064 6 data_out[2]
port 121 nsew signal output
rlabel metal3 s 0 78288 400 78344 6 data_out[30]
port 122 nsew signal output
rlabel metal3 s 0 76048 400 76104 6 data_out[31]
port 123 nsew signal output
rlabel metal3 s 0 73808 400 73864 6 data_out[32]
port 124 nsew signal output
rlabel metal3 s 0 71568 400 71624 6 data_out[33]
port 125 nsew signal output
rlabel metal3 s 0 69328 400 69384 6 data_out[34]
port 126 nsew signal output
rlabel metal3 s 0 67088 400 67144 6 data_out[35]
port 127 nsew signal output
rlabel metal3 s 0 64848 400 64904 6 data_out[36]
port 128 nsew signal output
rlabel metal3 s 0 62608 400 62664 6 data_out[37]
port 129 nsew signal output
rlabel metal3 s 0 60368 400 60424 6 data_out[38]
port 130 nsew signal output
rlabel metal3 s 0 58128 400 58184 6 data_out[39]
port 131 nsew signal output
rlabel metal3 s 0 138768 400 138824 6 data_out[3]
port 132 nsew signal output
rlabel metal3 s 0 55888 400 55944 6 data_out[40]
port 133 nsew signal output
rlabel metal3 s 0 53648 400 53704 6 data_out[41]
port 134 nsew signal output
rlabel metal3 s 0 51408 400 51464 6 data_out[42]
port 135 nsew signal output
rlabel metal3 s 0 49168 400 49224 6 data_out[43]
port 136 nsew signal output
rlabel metal3 s 0 46928 400 46984 6 data_out[44]
port 137 nsew signal output
rlabel metal3 s 0 44688 400 44744 6 data_out[45]
port 138 nsew signal output
rlabel metal3 s 0 42448 400 42504 6 data_out[46]
port 139 nsew signal output
rlabel metal3 s 0 40208 400 40264 6 data_out[47]
port 140 nsew signal output
rlabel metal3 s 0 37968 400 38024 6 data_out[48]
port 141 nsew signal output
rlabel metal3 s 0 35728 400 35784 6 data_out[49]
port 142 nsew signal output
rlabel metal3 s 0 136528 400 136584 6 data_out[4]
port 143 nsew signal output
rlabel metal3 s 0 33488 400 33544 6 data_out[50]
port 144 nsew signal output
rlabel metal3 s 0 31248 400 31304 6 data_out[51]
port 145 nsew signal output
rlabel metal3 s 0 29008 400 29064 6 data_out[52]
port 146 nsew signal output
rlabel metal3 s 0 26768 400 26824 6 data_out[53]
port 147 nsew signal output
rlabel metal3 s 0 24528 400 24584 6 data_out[54]
port 148 nsew signal output
rlabel metal3 s 0 22288 400 22344 6 data_out[55]
port 149 nsew signal output
rlabel metal3 s 0 20048 400 20104 6 data_out[56]
port 150 nsew signal output
rlabel metal3 s 0 17808 400 17864 6 data_out[57]
port 151 nsew signal output
rlabel metal3 s 0 15568 400 15624 6 data_out[58]
port 152 nsew signal output
rlabel metal3 s 0 13328 400 13384 6 data_out[59]
port 153 nsew signal output
rlabel metal3 s 0 134288 400 134344 6 data_out[5]
port 154 nsew signal output
rlabel metal3 s 0 11088 400 11144 6 data_out[60]
port 155 nsew signal output
rlabel metal3 s 0 8848 400 8904 6 data_out[61]
port 156 nsew signal output
rlabel metal3 s 0 6608 400 6664 6 data_out[62]
port 157 nsew signal output
rlabel metal3 s 0 4368 400 4424 6 data_out[63]
port 158 nsew signal output
rlabel metal3 s 0 132048 400 132104 6 data_out[6]
port 159 nsew signal output
rlabel metal3 s 0 129808 400 129864 6 data_out[7]
port 160 nsew signal output
rlabel metal3 s 0 127568 400 127624 6 data_out[8]
port 161 nsew signal output
rlabel metal3 s 0 125328 400 125384 6 data_out[9]
port 162 nsew signal output
rlabel metal2 s 6832 0 6888 400 6 stb
port 163 nsew signal input
rlabel metal4 s 2224 1538 2384 148206 6 vdd
port 164 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 148206 6 vdd
port 164 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 148206 6 vdd
port 164 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 148206 6 vdd
port 164 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 148206 6 vdd
port 164 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 148206 6 vdd
port 164 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 148206 6 vdd
port 164 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 148206 6 vdd
port 164 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 148206 6 vdd
port 164 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 148206 6 vdd
port 164 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 148206 6 vss
port 165 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 148206 6 vss
port 165 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 148206 6 vss
port 165 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 148206 6 vss
port 165 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 148206 6 vss
port 165 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 148206 6 vss
port 165 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 148206 6 vss
port 165 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 148206 6 vss
port 165 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 148206 6 vss
port 165 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 148206 6 vss
port 165 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 150000 150000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 33126100
string GDS_FILE /home/thomas/Documents/Projects/tilerisc/openlane/gpu_core/runs/23_12_08_22_57/results/signoff/gpu_core.magic.gds
string GDS_START 492804
<< end >>

