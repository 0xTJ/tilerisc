magic
tech gf180mcuD
magscale 1 5
timestamp 1702302053
<< obsm1 >>
rect 672 855 279328 174078
<< metal2 >>
rect 5040 0 5096 400
rect 5936 0 5992 400
rect 6832 0 6888 400
rect 7728 0 7784 400
rect 8624 0 8680 400
rect 9520 0 9576 400
rect 10416 0 10472 400
rect 11312 0 11368 400
rect 12208 0 12264 400
rect 13104 0 13160 400
rect 14000 0 14056 400
rect 14896 0 14952 400
rect 15792 0 15848 400
rect 16688 0 16744 400
rect 17584 0 17640 400
rect 18480 0 18536 400
rect 19376 0 19432 400
rect 20272 0 20328 400
rect 21168 0 21224 400
rect 22064 0 22120 400
rect 22960 0 23016 400
rect 23856 0 23912 400
rect 24752 0 24808 400
rect 25648 0 25704 400
rect 26544 0 26600 400
rect 27440 0 27496 400
rect 28336 0 28392 400
rect 29232 0 29288 400
rect 30128 0 30184 400
rect 31024 0 31080 400
rect 31920 0 31976 400
rect 32816 0 32872 400
rect 33712 0 33768 400
rect 34608 0 34664 400
rect 35504 0 35560 400
rect 36400 0 36456 400
rect 37296 0 37352 400
rect 38192 0 38248 400
rect 39088 0 39144 400
rect 39984 0 40040 400
rect 40880 0 40936 400
rect 41776 0 41832 400
rect 42672 0 42728 400
rect 43568 0 43624 400
rect 44464 0 44520 400
rect 45360 0 45416 400
rect 46256 0 46312 400
rect 47152 0 47208 400
rect 48048 0 48104 400
rect 48944 0 49000 400
rect 49840 0 49896 400
rect 50736 0 50792 400
rect 51632 0 51688 400
rect 52528 0 52584 400
rect 53424 0 53480 400
rect 54320 0 54376 400
rect 55216 0 55272 400
rect 56112 0 56168 400
rect 57008 0 57064 400
rect 57904 0 57960 400
rect 58800 0 58856 400
rect 59696 0 59752 400
rect 60592 0 60648 400
rect 61488 0 61544 400
rect 62384 0 62440 400
rect 63280 0 63336 400
rect 64176 0 64232 400
rect 65072 0 65128 400
rect 65968 0 66024 400
rect 66864 0 66920 400
rect 67760 0 67816 400
rect 68656 0 68712 400
rect 69552 0 69608 400
rect 70448 0 70504 400
rect 71344 0 71400 400
rect 72240 0 72296 400
rect 73136 0 73192 400
rect 74032 0 74088 400
rect 74928 0 74984 400
rect 75824 0 75880 400
rect 76720 0 76776 400
rect 77616 0 77672 400
rect 78512 0 78568 400
rect 79408 0 79464 400
rect 80304 0 80360 400
rect 81200 0 81256 400
rect 82096 0 82152 400
rect 82992 0 83048 400
rect 83888 0 83944 400
rect 84784 0 84840 400
rect 85680 0 85736 400
rect 86576 0 86632 400
rect 87472 0 87528 400
rect 88368 0 88424 400
rect 89264 0 89320 400
rect 90160 0 90216 400
rect 91056 0 91112 400
rect 91952 0 92008 400
rect 92848 0 92904 400
rect 93744 0 93800 400
rect 94640 0 94696 400
rect 95536 0 95592 400
rect 96432 0 96488 400
rect 97328 0 97384 400
rect 98224 0 98280 400
rect 99120 0 99176 400
rect 100016 0 100072 400
rect 100912 0 100968 400
rect 101808 0 101864 400
rect 102704 0 102760 400
rect 103600 0 103656 400
rect 104496 0 104552 400
rect 105392 0 105448 400
rect 106288 0 106344 400
rect 107184 0 107240 400
rect 108080 0 108136 400
rect 108976 0 109032 400
rect 109872 0 109928 400
rect 110768 0 110824 400
rect 111664 0 111720 400
rect 112560 0 112616 400
rect 113456 0 113512 400
rect 114352 0 114408 400
rect 115248 0 115304 400
rect 116144 0 116200 400
rect 117040 0 117096 400
rect 117936 0 117992 400
rect 118832 0 118888 400
rect 119728 0 119784 400
rect 120624 0 120680 400
rect 121520 0 121576 400
rect 122416 0 122472 400
rect 123312 0 123368 400
rect 124208 0 124264 400
rect 125104 0 125160 400
rect 126000 0 126056 400
rect 126896 0 126952 400
rect 127792 0 127848 400
rect 128688 0 128744 400
rect 129584 0 129640 400
rect 130480 0 130536 400
rect 131376 0 131432 400
rect 132272 0 132328 400
rect 133168 0 133224 400
rect 134064 0 134120 400
rect 134960 0 135016 400
rect 135856 0 135912 400
rect 136752 0 136808 400
rect 137648 0 137704 400
rect 138544 0 138600 400
rect 139440 0 139496 400
rect 140336 0 140392 400
rect 141232 0 141288 400
rect 142128 0 142184 400
rect 143024 0 143080 400
rect 143920 0 143976 400
rect 144816 0 144872 400
rect 145712 0 145768 400
rect 146608 0 146664 400
rect 147504 0 147560 400
rect 148400 0 148456 400
rect 149296 0 149352 400
rect 150192 0 150248 400
rect 151088 0 151144 400
rect 151984 0 152040 400
rect 152880 0 152936 400
rect 153776 0 153832 400
rect 154672 0 154728 400
rect 155568 0 155624 400
rect 156464 0 156520 400
rect 157360 0 157416 400
rect 158256 0 158312 400
rect 159152 0 159208 400
rect 160048 0 160104 400
rect 160944 0 161000 400
rect 161840 0 161896 400
rect 162736 0 162792 400
rect 163632 0 163688 400
rect 164528 0 164584 400
rect 165424 0 165480 400
rect 166320 0 166376 400
rect 167216 0 167272 400
rect 168112 0 168168 400
rect 169008 0 169064 400
rect 169904 0 169960 400
rect 170800 0 170856 400
rect 171696 0 171752 400
rect 172592 0 172648 400
rect 173488 0 173544 400
rect 174384 0 174440 400
rect 175280 0 175336 400
rect 176176 0 176232 400
rect 177072 0 177128 400
rect 177968 0 178024 400
rect 178864 0 178920 400
rect 179760 0 179816 400
rect 180656 0 180712 400
rect 181552 0 181608 400
rect 182448 0 182504 400
rect 183344 0 183400 400
rect 184240 0 184296 400
rect 185136 0 185192 400
rect 186032 0 186088 400
rect 186928 0 186984 400
rect 187824 0 187880 400
rect 188720 0 188776 400
rect 189616 0 189672 400
rect 190512 0 190568 400
rect 191408 0 191464 400
rect 192304 0 192360 400
rect 193200 0 193256 400
rect 194096 0 194152 400
rect 194992 0 195048 400
rect 195888 0 195944 400
rect 196784 0 196840 400
rect 197680 0 197736 400
rect 198576 0 198632 400
rect 199472 0 199528 400
rect 200368 0 200424 400
rect 201264 0 201320 400
rect 202160 0 202216 400
rect 203056 0 203112 400
rect 203952 0 204008 400
rect 204848 0 204904 400
rect 205744 0 205800 400
rect 206640 0 206696 400
rect 207536 0 207592 400
rect 208432 0 208488 400
rect 209328 0 209384 400
rect 210224 0 210280 400
rect 211120 0 211176 400
rect 212016 0 212072 400
rect 212912 0 212968 400
rect 213808 0 213864 400
rect 214704 0 214760 400
rect 215600 0 215656 400
rect 216496 0 216552 400
rect 217392 0 217448 400
rect 218288 0 218344 400
rect 219184 0 219240 400
rect 220080 0 220136 400
rect 220976 0 221032 400
rect 221872 0 221928 400
rect 222768 0 222824 400
rect 223664 0 223720 400
rect 224560 0 224616 400
rect 225456 0 225512 400
rect 226352 0 226408 400
rect 227248 0 227304 400
rect 228144 0 228200 400
rect 229040 0 229096 400
rect 229936 0 229992 400
rect 230832 0 230888 400
rect 231728 0 231784 400
rect 232624 0 232680 400
rect 233520 0 233576 400
rect 234416 0 234472 400
rect 235312 0 235368 400
rect 236208 0 236264 400
rect 237104 0 237160 400
rect 238000 0 238056 400
rect 238896 0 238952 400
rect 239792 0 239848 400
rect 240688 0 240744 400
rect 241584 0 241640 400
rect 242480 0 242536 400
rect 243376 0 243432 400
rect 244272 0 244328 400
rect 245168 0 245224 400
rect 246064 0 246120 400
rect 246960 0 247016 400
rect 247856 0 247912 400
rect 248752 0 248808 400
rect 249648 0 249704 400
rect 250544 0 250600 400
rect 251440 0 251496 400
rect 252336 0 252392 400
rect 253232 0 253288 400
rect 254128 0 254184 400
rect 255024 0 255080 400
rect 255920 0 255976 400
rect 256816 0 256872 400
rect 257712 0 257768 400
rect 258608 0 258664 400
rect 259504 0 259560 400
rect 260400 0 260456 400
rect 261296 0 261352 400
rect 262192 0 262248 400
rect 263088 0 263144 400
rect 263984 0 264040 400
rect 264880 0 264936 400
rect 265776 0 265832 400
rect 266672 0 266728 400
rect 267568 0 267624 400
rect 268464 0 268520 400
rect 269360 0 269416 400
rect 270256 0 270312 400
rect 271152 0 271208 400
rect 272048 0 272104 400
rect 272944 0 273000 400
rect 273840 0 273896 400
rect 274736 0 274792 400
<< obsm2 >>
rect 854 430 279146 174067
rect 854 233 5010 430
rect 5126 233 5906 430
rect 6022 233 6802 430
rect 6918 233 7698 430
rect 7814 233 8594 430
rect 8710 233 9490 430
rect 9606 233 10386 430
rect 10502 233 11282 430
rect 11398 233 12178 430
rect 12294 233 13074 430
rect 13190 233 13970 430
rect 14086 233 14866 430
rect 14982 233 15762 430
rect 15878 233 16658 430
rect 16774 233 17554 430
rect 17670 233 18450 430
rect 18566 233 19346 430
rect 19462 233 20242 430
rect 20358 233 21138 430
rect 21254 233 22034 430
rect 22150 233 22930 430
rect 23046 233 23826 430
rect 23942 233 24722 430
rect 24838 233 25618 430
rect 25734 233 26514 430
rect 26630 233 27410 430
rect 27526 233 28306 430
rect 28422 233 29202 430
rect 29318 233 30098 430
rect 30214 233 30994 430
rect 31110 233 31890 430
rect 32006 233 32786 430
rect 32902 233 33682 430
rect 33798 233 34578 430
rect 34694 233 35474 430
rect 35590 233 36370 430
rect 36486 233 37266 430
rect 37382 233 38162 430
rect 38278 233 39058 430
rect 39174 233 39954 430
rect 40070 233 40850 430
rect 40966 233 41746 430
rect 41862 233 42642 430
rect 42758 233 43538 430
rect 43654 233 44434 430
rect 44550 233 45330 430
rect 45446 233 46226 430
rect 46342 233 47122 430
rect 47238 233 48018 430
rect 48134 233 48914 430
rect 49030 233 49810 430
rect 49926 233 50706 430
rect 50822 233 51602 430
rect 51718 233 52498 430
rect 52614 233 53394 430
rect 53510 233 54290 430
rect 54406 233 55186 430
rect 55302 233 56082 430
rect 56198 233 56978 430
rect 57094 233 57874 430
rect 57990 233 58770 430
rect 58886 233 59666 430
rect 59782 233 60562 430
rect 60678 233 61458 430
rect 61574 233 62354 430
rect 62470 233 63250 430
rect 63366 233 64146 430
rect 64262 233 65042 430
rect 65158 233 65938 430
rect 66054 233 66834 430
rect 66950 233 67730 430
rect 67846 233 68626 430
rect 68742 233 69522 430
rect 69638 233 70418 430
rect 70534 233 71314 430
rect 71430 233 72210 430
rect 72326 233 73106 430
rect 73222 233 74002 430
rect 74118 233 74898 430
rect 75014 233 75794 430
rect 75910 233 76690 430
rect 76806 233 77586 430
rect 77702 233 78482 430
rect 78598 233 79378 430
rect 79494 233 80274 430
rect 80390 233 81170 430
rect 81286 233 82066 430
rect 82182 233 82962 430
rect 83078 233 83858 430
rect 83974 233 84754 430
rect 84870 233 85650 430
rect 85766 233 86546 430
rect 86662 233 87442 430
rect 87558 233 88338 430
rect 88454 233 89234 430
rect 89350 233 90130 430
rect 90246 233 91026 430
rect 91142 233 91922 430
rect 92038 233 92818 430
rect 92934 233 93714 430
rect 93830 233 94610 430
rect 94726 233 95506 430
rect 95622 233 96402 430
rect 96518 233 97298 430
rect 97414 233 98194 430
rect 98310 233 99090 430
rect 99206 233 99986 430
rect 100102 233 100882 430
rect 100998 233 101778 430
rect 101894 233 102674 430
rect 102790 233 103570 430
rect 103686 233 104466 430
rect 104582 233 105362 430
rect 105478 233 106258 430
rect 106374 233 107154 430
rect 107270 233 108050 430
rect 108166 233 108946 430
rect 109062 233 109842 430
rect 109958 233 110738 430
rect 110854 233 111634 430
rect 111750 233 112530 430
rect 112646 233 113426 430
rect 113542 233 114322 430
rect 114438 233 115218 430
rect 115334 233 116114 430
rect 116230 233 117010 430
rect 117126 233 117906 430
rect 118022 233 118802 430
rect 118918 233 119698 430
rect 119814 233 120594 430
rect 120710 233 121490 430
rect 121606 233 122386 430
rect 122502 233 123282 430
rect 123398 233 124178 430
rect 124294 233 125074 430
rect 125190 233 125970 430
rect 126086 233 126866 430
rect 126982 233 127762 430
rect 127878 233 128658 430
rect 128774 233 129554 430
rect 129670 233 130450 430
rect 130566 233 131346 430
rect 131462 233 132242 430
rect 132358 233 133138 430
rect 133254 233 134034 430
rect 134150 233 134930 430
rect 135046 233 135826 430
rect 135942 233 136722 430
rect 136838 233 137618 430
rect 137734 233 138514 430
rect 138630 233 139410 430
rect 139526 233 140306 430
rect 140422 233 141202 430
rect 141318 233 142098 430
rect 142214 233 142994 430
rect 143110 233 143890 430
rect 144006 233 144786 430
rect 144902 233 145682 430
rect 145798 233 146578 430
rect 146694 233 147474 430
rect 147590 233 148370 430
rect 148486 233 149266 430
rect 149382 233 150162 430
rect 150278 233 151058 430
rect 151174 233 151954 430
rect 152070 233 152850 430
rect 152966 233 153746 430
rect 153862 233 154642 430
rect 154758 233 155538 430
rect 155654 233 156434 430
rect 156550 233 157330 430
rect 157446 233 158226 430
rect 158342 233 159122 430
rect 159238 233 160018 430
rect 160134 233 160914 430
rect 161030 233 161810 430
rect 161926 233 162706 430
rect 162822 233 163602 430
rect 163718 233 164498 430
rect 164614 233 165394 430
rect 165510 233 166290 430
rect 166406 233 167186 430
rect 167302 233 168082 430
rect 168198 233 168978 430
rect 169094 233 169874 430
rect 169990 233 170770 430
rect 170886 233 171666 430
rect 171782 233 172562 430
rect 172678 233 173458 430
rect 173574 233 174354 430
rect 174470 233 175250 430
rect 175366 233 176146 430
rect 176262 233 177042 430
rect 177158 233 177938 430
rect 178054 233 178834 430
rect 178950 233 179730 430
rect 179846 233 180626 430
rect 180742 233 181522 430
rect 181638 233 182418 430
rect 182534 233 183314 430
rect 183430 233 184210 430
rect 184326 233 185106 430
rect 185222 233 186002 430
rect 186118 233 186898 430
rect 187014 233 187794 430
rect 187910 233 188690 430
rect 188806 233 189586 430
rect 189702 233 190482 430
rect 190598 233 191378 430
rect 191494 233 192274 430
rect 192390 233 193170 430
rect 193286 233 194066 430
rect 194182 233 194962 430
rect 195078 233 195858 430
rect 195974 233 196754 430
rect 196870 233 197650 430
rect 197766 233 198546 430
rect 198662 233 199442 430
rect 199558 233 200338 430
rect 200454 233 201234 430
rect 201350 233 202130 430
rect 202246 233 203026 430
rect 203142 233 203922 430
rect 204038 233 204818 430
rect 204934 233 205714 430
rect 205830 233 206610 430
rect 206726 233 207506 430
rect 207622 233 208402 430
rect 208518 233 209298 430
rect 209414 233 210194 430
rect 210310 233 211090 430
rect 211206 233 211986 430
rect 212102 233 212882 430
rect 212998 233 213778 430
rect 213894 233 214674 430
rect 214790 233 215570 430
rect 215686 233 216466 430
rect 216582 233 217362 430
rect 217478 233 218258 430
rect 218374 233 219154 430
rect 219270 233 220050 430
rect 220166 233 220946 430
rect 221062 233 221842 430
rect 221958 233 222738 430
rect 222854 233 223634 430
rect 223750 233 224530 430
rect 224646 233 225426 430
rect 225542 233 226322 430
rect 226438 233 227218 430
rect 227334 233 228114 430
rect 228230 233 229010 430
rect 229126 233 229906 430
rect 230022 233 230802 430
rect 230918 233 231698 430
rect 231814 233 232594 430
rect 232710 233 233490 430
rect 233606 233 234386 430
rect 234502 233 235282 430
rect 235398 233 236178 430
rect 236294 233 237074 430
rect 237190 233 237970 430
rect 238086 233 238866 430
rect 238982 233 239762 430
rect 239878 233 240658 430
rect 240774 233 241554 430
rect 241670 233 242450 430
rect 242566 233 243346 430
rect 243462 233 244242 430
rect 244358 233 245138 430
rect 245254 233 246034 430
rect 246150 233 246930 430
rect 247046 233 247826 430
rect 247942 233 248722 430
rect 248838 233 249618 430
rect 249734 233 250514 430
rect 250630 233 251410 430
rect 251526 233 252306 430
rect 252422 233 253202 430
rect 253318 233 254098 430
rect 254214 233 254994 430
rect 255110 233 255890 430
rect 256006 233 256786 430
rect 256902 233 257682 430
rect 257798 233 258578 430
rect 258694 233 259474 430
rect 259590 233 260370 430
rect 260486 233 261266 430
rect 261382 233 262162 430
rect 262278 233 263058 430
rect 263174 233 263954 430
rect 264070 233 264850 430
rect 264966 233 265746 430
rect 265862 233 266642 430
rect 266758 233 267538 430
rect 267654 233 268434 430
rect 268550 233 269330 430
rect 269446 233 270226 430
rect 270342 233 271122 430
rect 271238 233 272018 430
rect 272134 233 272914 430
rect 273030 233 273810 430
rect 273926 233 274706 430
rect 274822 233 279146 430
<< metal3 >>
rect 0 171696 400 171752
rect 279600 171696 280000 171752
rect 0 164416 400 164472
rect 279600 164416 280000 164472
rect 0 157136 400 157192
rect 279600 157136 280000 157192
rect 0 149856 400 149912
rect 279600 149856 280000 149912
rect 0 142576 400 142632
rect 279600 142576 280000 142632
rect 0 135296 400 135352
rect 279600 135296 280000 135352
rect 0 128016 400 128072
rect 279600 128016 280000 128072
rect 0 120736 400 120792
rect 279600 120736 280000 120792
rect 0 113456 400 113512
rect 279600 113456 280000 113512
rect 0 106176 400 106232
rect 279600 106176 280000 106232
rect 0 98896 400 98952
rect 279600 98896 280000 98952
rect 0 91616 400 91672
rect 279600 91616 280000 91672
rect 0 84336 400 84392
rect 279600 84336 280000 84392
rect 0 77056 400 77112
rect 279600 77056 280000 77112
rect 0 69776 400 69832
rect 279600 69776 280000 69832
rect 0 62496 400 62552
rect 279600 62496 280000 62552
rect 0 55216 400 55272
rect 279600 55216 280000 55272
rect 0 47936 400 47992
rect 279600 47936 280000 47992
rect 0 40656 400 40712
rect 279600 40656 280000 40712
rect 0 33376 400 33432
rect 279600 33376 280000 33432
rect 0 26096 400 26152
rect 279600 26096 280000 26152
rect 0 18816 400 18872
rect 279600 18816 280000 18872
rect 0 11536 400 11592
rect 279600 11536 280000 11592
rect 0 4256 400 4312
rect 279600 4256 280000 4312
<< obsm3 >>
rect 400 171782 279650 174062
rect 430 171666 279570 171782
rect 400 164502 279650 171666
rect 430 164386 279570 164502
rect 400 157222 279650 164386
rect 430 157106 279570 157222
rect 400 149942 279650 157106
rect 430 149826 279570 149942
rect 400 142662 279650 149826
rect 430 142546 279570 142662
rect 400 135382 279650 142546
rect 430 135266 279570 135382
rect 400 128102 279650 135266
rect 430 127986 279570 128102
rect 400 120822 279650 127986
rect 430 120706 279570 120822
rect 400 113542 279650 120706
rect 430 113426 279570 113542
rect 400 106262 279650 113426
rect 430 106146 279570 106262
rect 400 98982 279650 106146
rect 430 98866 279570 98982
rect 400 91702 279650 98866
rect 430 91586 279570 91702
rect 400 84422 279650 91586
rect 430 84306 279570 84422
rect 400 77142 279650 84306
rect 430 77026 279570 77142
rect 400 69862 279650 77026
rect 430 69746 279570 69862
rect 400 62582 279650 69746
rect 430 62466 279570 62582
rect 400 55302 279650 62466
rect 430 55186 279570 55302
rect 400 48022 279650 55186
rect 430 47906 279570 48022
rect 400 40742 279650 47906
rect 430 40626 279570 40742
rect 400 33462 279650 40626
rect 430 33346 279570 33462
rect 400 26182 279650 33346
rect 430 26066 279570 26182
rect 400 18902 279650 26066
rect 430 18786 279570 18902
rect 400 11622 279650 18786
rect 430 11506 279570 11622
rect 400 4342 279650 11506
rect 430 4226 279570 4342
rect 400 238 279650 4226
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< obsm4 >>
rect 8134 1508 9874 67247
rect 10094 1508 17554 67247
rect 17774 1508 25234 67247
rect 25454 1508 32914 67247
rect 33134 1508 40594 67247
rect 40814 1508 48274 67247
rect 48494 1508 55954 67247
rect 56174 1508 63634 67247
rect 63854 1508 71314 67247
rect 71534 1508 78994 67247
rect 79214 1508 86674 67247
rect 86894 1508 94354 67247
rect 94574 1508 102034 67247
rect 102254 1508 109714 67247
rect 109934 1508 117394 67247
rect 117614 1508 125074 67247
rect 125294 1508 132754 67247
rect 132974 1508 140434 67247
rect 140654 1508 148114 67247
rect 148334 1508 155794 67247
rect 156014 1508 163474 67247
rect 163694 1508 171154 67247
rect 171374 1508 178834 67247
rect 179054 1508 186514 67247
rect 186734 1508 194194 67247
rect 194414 1508 201874 67247
rect 202094 1508 204106 67247
rect 8134 345 204106 1508
<< labels >>
rlabel metal3 s 279600 4256 280000 4312 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 128016 400 128072 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 106176 400 106232 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 84336 400 84392 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 62496 400 62552 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 40656 400 40712 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 18816 400 18872 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 279600 26096 280000 26152 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 279600 47936 280000 47992 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 279600 69776 280000 69832 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 279600 91616 280000 91672 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 279600 113456 280000 113512 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 279600 135296 280000 135352 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 279600 157136 280000 157192 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 171696 400 171752 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 149856 400 149912 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 279600 18816 280000 18872 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 113456 400 113512 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 91616 400 91672 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 69776 400 69832 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 47936 400 47992 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 26096 400 26152 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 4256 400 4312 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 279600 40656 280000 40712 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 279600 62496 280000 62552 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 279600 84336 280000 84392 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 279600 106176 280000 106232 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 279600 128016 280000 128072 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 279600 149856 280000 149912 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 279600 171696 280000 171752 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 157136 400 157192 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 135296 400 135352 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 279600 11536 280000 11592 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 120736 400 120792 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 98896 400 98952 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 77056 400 77112 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 55216 400 55272 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 33376 400 33432 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 11536 400 11592 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 279600 33376 280000 33432 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 279600 55216 280000 55272 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 279600 77056 280000 77112 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 279600 98896 280000 98952 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 279600 120736 280000 120792 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 279600 142576 280000 142632 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 279600 164416 280000 164472 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 164416 400 164472 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 142576 400 142632 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 272048 0 272104 400 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 272944 0 273000 400 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 273840 0 273896 400 6 irq[2]
port 51 nsew signal output
rlabel metal2 s 100016 0 100072 400 6 la_data_in[0]
port 52 nsew signal input
rlabel metal2 s 126896 0 126952 400 6 la_data_in[10]
port 53 nsew signal input
rlabel metal2 s 129584 0 129640 400 6 la_data_in[11]
port 54 nsew signal input
rlabel metal2 s 132272 0 132328 400 6 la_data_in[12]
port 55 nsew signal input
rlabel metal2 s 134960 0 135016 400 6 la_data_in[13]
port 56 nsew signal input
rlabel metal2 s 137648 0 137704 400 6 la_data_in[14]
port 57 nsew signal input
rlabel metal2 s 140336 0 140392 400 6 la_data_in[15]
port 58 nsew signal input
rlabel metal2 s 143024 0 143080 400 6 la_data_in[16]
port 59 nsew signal input
rlabel metal2 s 145712 0 145768 400 6 la_data_in[17]
port 60 nsew signal input
rlabel metal2 s 148400 0 148456 400 6 la_data_in[18]
port 61 nsew signal input
rlabel metal2 s 151088 0 151144 400 6 la_data_in[19]
port 62 nsew signal input
rlabel metal2 s 102704 0 102760 400 6 la_data_in[1]
port 63 nsew signal input
rlabel metal2 s 153776 0 153832 400 6 la_data_in[20]
port 64 nsew signal input
rlabel metal2 s 156464 0 156520 400 6 la_data_in[21]
port 65 nsew signal input
rlabel metal2 s 159152 0 159208 400 6 la_data_in[22]
port 66 nsew signal input
rlabel metal2 s 161840 0 161896 400 6 la_data_in[23]
port 67 nsew signal input
rlabel metal2 s 164528 0 164584 400 6 la_data_in[24]
port 68 nsew signal input
rlabel metal2 s 167216 0 167272 400 6 la_data_in[25]
port 69 nsew signal input
rlabel metal2 s 169904 0 169960 400 6 la_data_in[26]
port 70 nsew signal input
rlabel metal2 s 172592 0 172648 400 6 la_data_in[27]
port 71 nsew signal input
rlabel metal2 s 175280 0 175336 400 6 la_data_in[28]
port 72 nsew signal input
rlabel metal2 s 177968 0 178024 400 6 la_data_in[29]
port 73 nsew signal input
rlabel metal2 s 105392 0 105448 400 6 la_data_in[2]
port 74 nsew signal input
rlabel metal2 s 180656 0 180712 400 6 la_data_in[30]
port 75 nsew signal input
rlabel metal2 s 183344 0 183400 400 6 la_data_in[31]
port 76 nsew signal input
rlabel metal2 s 186032 0 186088 400 6 la_data_in[32]
port 77 nsew signal input
rlabel metal2 s 188720 0 188776 400 6 la_data_in[33]
port 78 nsew signal input
rlabel metal2 s 191408 0 191464 400 6 la_data_in[34]
port 79 nsew signal input
rlabel metal2 s 194096 0 194152 400 6 la_data_in[35]
port 80 nsew signal input
rlabel metal2 s 196784 0 196840 400 6 la_data_in[36]
port 81 nsew signal input
rlabel metal2 s 199472 0 199528 400 6 la_data_in[37]
port 82 nsew signal input
rlabel metal2 s 202160 0 202216 400 6 la_data_in[38]
port 83 nsew signal input
rlabel metal2 s 204848 0 204904 400 6 la_data_in[39]
port 84 nsew signal input
rlabel metal2 s 108080 0 108136 400 6 la_data_in[3]
port 85 nsew signal input
rlabel metal2 s 207536 0 207592 400 6 la_data_in[40]
port 86 nsew signal input
rlabel metal2 s 210224 0 210280 400 6 la_data_in[41]
port 87 nsew signal input
rlabel metal2 s 212912 0 212968 400 6 la_data_in[42]
port 88 nsew signal input
rlabel metal2 s 215600 0 215656 400 6 la_data_in[43]
port 89 nsew signal input
rlabel metal2 s 218288 0 218344 400 6 la_data_in[44]
port 90 nsew signal input
rlabel metal2 s 220976 0 221032 400 6 la_data_in[45]
port 91 nsew signal input
rlabel metal2 s 223664 0 223720 400 6 la_data_in[46]
port 92 nsew signal input
rlabel metal2 s 226352 0 226408 400 6 la_data_in[47]
port 93 nsew signal input
rlabel metal2 s 229040 0 229096 400 6 la_data_in[48]
port 94 nsew signal input
rlabel metal2 s 231728 0 231784 400 6 la_data_in[49]
port 95 nsew signal input
rlabel metal2 s 110768 0 110824 400 6 la_data_in[4]
port 96 nsew signal input
rlabel metal2 s 234416 0 234472 400 6 la_data_in[50]
port 97 nsew signal input
rlabel metal2 s 237104 0 237160 400 6 la_data_in[51]
port 98 nsew signal input
rlabel metal2 s 239792 0 239848 400 6 la_data_in[52]
port 99 nsew signal input
rlabel metal2 s 242480 0 242536 400 6 la_data_in[53]
port 100 nsew signal input
rlabel metal2 s 245168 0 245224 400 6 la_data_in[54]
port 101 nsew signal input
rlabel metal2 s 247856 0 247912 400 6 la_data_in[55]
port 102 nsew signal input
rlabel metal2 s 250544 0 250600 400 6 la_data_in[56]
port 103 nsew signal input
rlabel metal2 s 253232 0 253288 400 6 la_data_in[57]
port 104 nsew signal input
rlabel metal2 s 255920 0 255976 400 6 la_data_in[58]
port 105 nsew signal input
rlabel metal2 s 258608 0 258664 400 6 la_data_in[59]
port 106 nsew signal input
rlabel metal2 s 113456 0 113512 400 6 la_data_in[5]
port 107 nsew signal input
rlabel metal2 s 261296 0 261352 400 6 la_data_in[60]
port 108 nsew signal input
rlabel metal2 s 263984 0 264040 400 6 la_data_in[61]
port 109 nsew signal input
rlabel metal2 s 266672 0 266728 400 6 la_data_in[62]
port 110 nsew signal input
rlabel metal2 s 269360 0 269416 400 6 la_data_in[63]
port 111 nsew signal input
rlabel metal2 s 116144 0 116200 400 6 la_data_in[6]
port 112 nsew signal input
rlabel metal2 s 118832 0 118888 400 6 la_data_in[7]
port 113 nsew signal input
rlabel metal2 s 121520 0 121576 400 6 la_data_in[8]
port 114 nsew signal input
rlabel metal2 s 124208 0 124264 400 6 la_data_in[9]
port 115 nsew signal input
rlabel metal2 s 100912 0 100968 400 6 la_data_out[0]
port 116 nsew signal output
rlabel metal2 s 127792 0 127848 400 6 la_data_out[10]
port 117 nsew signal output
rlabel metal2 s 130480 0 130536 400 6 la_data_out[11]
port 118 nsew signal output
rlabel metal2 s 133168 0 133224 400 6 la_data_out[12]
port 119 nsew signal output
rlabel metal2 s 135856 0 135912 400 6 la_data_out[13]
port 120 nsew signal output
rlabel metal2 s 138544 0 138600 400 6 la_data_out[14]
port 121 nsew signal output
rlabel metal2 s 141232 0 141288 400 6 la_data_out[15]
port 122 nsew signal output
rlabel metal2 s 143920 0 143976 400 6 la_data_out[16]
port 123 nsew signal output
rlabel metal2 s 146608 0 146664 400 6 la_data_out[17]
port 124 nsew signal output
rlabel metal2 s 149296 0 149352 400 6 la_data_out[18]
port 125 nsew signal output
rlabel metal2 s 151984 0 152040 400 6 la_data_out[19]
port 126 nsew signal output
rlabel metal2 s 103600 0 103656 400 6 la_data_out[1]
port 127 nsew signal output
rlabel metal2 s 154672 0 154728 400 6 la_data_out[20]
port 128 nsew signal output
rlabel metal2 s 157360 0 157416 400 6 la_data_out[21]
port 129 nsew signal output
rlabel metal2 s 160048 0 160104 400 6 la_data_out[22]
port 130 nsew signal output
rlabel metal2 s 162736 0 162792 400 6 la_data_out[23]
port 131 nsew signal output
rlabel metal2 s 165424 0 165480 400 6 la_data_out[24]
port 132 nsew signal output
rlabel metal2 s 168112 0 168168 400 6 la_data_out[25]
port 133 nsew signal output
rlabel metal2 s 170800 0 170856 400 6 la_data_out[26]
port 134 nsew signal output
rlabel metal2 s 173488 0 173544 400 6 la_data_out[27]
port 135 nsew signal output
rlabel metal2 s 176176 0 176232 400 6 la_data_out[28]
port 136 nsew signal output
rlabel metal2 s 178864 0 178920 400 6 la_data_out[29]
port 137 nsew signal output
rlabel metal2 s 106288 0 106344 400 6 la_data_out[2]
port 138 nsew signal output
rlabel metal2 s 181552 0 181608 400 6 la_data_out[30]
port 139 nsew signal output
rlabel metal2 s 184240 0 184296 400 6 la_data_out[31]
port 140 nsew signal output
rlabel metal2 s 186928 0 186984 400 6 la_data_out[32]
port 141 nsew signal output
rlabel metal2 s 189616 0 189672 400 6 la_data_out[33]
port 142 nsew signal output
rlabel metal2 s 192304 0 192360 400 6 la_data_out[34]
port 143 nsew signal output
rlabel metal2 s 194992 0 195048 400 6 la_data_out[35]
port 144 nsew signal output
rlabel metal2 s 197680 0 197736 400 6 la_data_out[36]
port 145 nsew signal output
rlabel metal2 s 200368 0 200424 400 6 la_data_out[37]
port 146 nsew signal output
rlabel metal2 s 203056 0 203112 400 6 la_data_out[38]
port 147 nsew signal output
rlabel metal2 s 205744 0 205800 400 6 la_data_out[39]
port 148 nsew signal output
rlabel metal2 s 108976 0 109032 400 6 la_data_out[3]
port 149 nsew signal output
rlabel metal2 s 208432 0 208488 400 6 la_data_out[40]
port 150 nsew signal output
rlabel metal2 s 211120 0 211176 400 6 la_data_out[41]
port 151 nsew signal output
rlabel metal2 s 213808 0 213864 400 6 la_data_out[42]
port 152 nsew signal output
rlabel metal2 s 216496 0 216552 400 6 la_data_out[43]
port 153 nsew signal output
rlabel metal2 s 219184 0 219240 400 6 la_data_out[44]
port 154 nsew signal output
rlabel metal2 s 221872 0 221928 400 6 la_data_out[45]
port 155 nsew signal output
rlabel metal2 s 224560 0 224616 400 6 la_data_out[46]
port 156 nsew signal output
rlabel metal2 s 227248 0 227304 400 6 la_data_out[47]
port 157 nsew signal output
rlabel metal2 s 229936 0 229992 400 6 la_data_out[48]
port 158 nsew signal output
rlabel metal2 s 232624 0 232680 400 6 la_data_out[49]
port 159 nsew signal output
rlabel metal2 s 111664 0 111720 400 6 la_data_out[4]
port 160 nsew signal output
rlabel metal2 s 235312 0 235368 400 6 la_data_out[50]
port 161 nsew signal output
rlabel metal2 s 238000 0 238056 400 6 la_data_out[51]
port 162 nsew signal output
rlabel metal2 s 240688 0 240744 400 6 la_data_out[52]
port 163 nsew signal output
rlabel metal2 s 243376 0 243432 400 6 la_data_out[53]
port 164 nsew signal output
rlabel metal2 s 246064 0 246120 400 6 la_data_out[54]
port 165 nsew signal output
rlabel metal2 s 248752 0 248808 400 6 la_data_out[55]
port 166 nsew signal output
rlabel metal2 s 251440 0 251496 400 6 la_data_out[56]
port 167 nsew signal output
rlabel metal2 s 254128 0 254184 400 6 la_data_out[57]
port 168 nsew signal output
rlabel metal2 s 256816 0 256872 400 6 la_data_out[58]
port 169 nsew signal output
rlabel metal2 s 259504 0 259560 400 6 la_data_out[59]
port 170 nsew signal output
rlabel metal2 s 114352 0 114408 400 6 la_data_out[5]
port 171 nsew signal output
rlabel metal2 s 262192 0 262248 400 6 la_data_out[60]
port 172 nsew signal output
rlabel metal2 s 264880 0 264936 400 6 la_data_out[61]
port 173 nsew signal output
rlabel metal2 s 267568 0 267624 400 6 la_data_out[62]
port 174 nsew signal output
rlabel metal2 s 270256 0 270312 400 6 la_data_out[63]
port 175 nsew signal output
rlabel metal2 s 117040 0 117096 400 6 la_data_out[6]
port 176 nsew signal output
rlabel metal2 s 119728 0 119784 400 6 la_data_out[7]
port 177 nsew signal output
rlabel metal2 s 122416 0 122472 400 6 la_data_out[8]
port 178 nsew signal output
rlabel metal2 s 125104 0 125160 400 6 la_data_out[9]
port 179 nsew signal output
rlabel metal2 s 101808 0 101864 400 6 la_oenb[0]
port 180 nsew signal input
rlabel metal2 s 128688 0 128744 400 6 la_oenb[10]
port 181 nsew signal input
rlabel metal2 s 131376 0 131432 400 6 la_oenb[11]
port 182 nsew signal input
rlabel metal2 s 134064 0 134120 400 6 la_oenb[12]
port 183 nsew signal input
rlabel metal2 s 136752 0 136808 400 6 la_oenb[13]
port 184 nsew signal input
rlabel metal2 s 139440 0 139496 400 6 la_oenb[14]
port 185 nsew signal input
rlabel metal2 s 142128 0 142184 400 6 la_oenb[15]
port 186 nsew signal input
rlabel metal2 s 144816 0 144872 400 6 la_oenb[16]
port 187 nsew signal input
rlabel metal2 s 147504 0 147560 400 6 la_oenb[17]
port 188 nsew signal input
rlabel metal2 s 150192 0 150248 400 6 la_oenb[18]
port 189 nsew signal input
rlabel metal2 s 152880 0 152936 400 6 la_oenb[19]
port 190 nsew signal input
rlabel metal2 s 104496 0 104552 400 6 la_oenb[1]
port 191 nsew signal input
rlabel metal2 s 155568 0 155624 400 6 la_oenb[20]
port 192 nsew signal input
rlabel metal2 s 158256 0 158312 400 6 la_oenb[21]
port 193 nsew signal input
rlabel metal2 s 160944 0 161000 400 6 la_oenb[22]
port 194 nsew signal input
rlabel metal2 s 163632 0 163688 400 6 la_oenb[23]
port 195 nsew signal input
rlabel metal2 s 166320 0 166376 400 6 la_oenb[24]
port 196 nsew signal input
rlabel metal2 s 169008 0 169064 400 6 la_oenb[25]
port 197 nsew signal input
rlabel metal2 s 171696 0 171752 400 6 la_oenb[26]
port 198 nsew signal input
rlabel metal2 s 174384 0 174440 400 6 la_oenb[27]
port 199 nsew signal input
rlabel metal2 s 177072 0 177128 400 6 la_oenb[28]
port 200 nsew signal input
rlabel metal2 s 179760 0 179816 400 6 la_oenb[29]
port 201 nsew signal input
rlabel metal2 s 107184 0 107240 400 6 la_oenb[2]
port 202 nsew signal input
rlabel metal2 s 182448 0 182504 400 6 la_oenb[30]
port 203 nsew signal input
rlabel metal2 s 185136 0 185192 400 6 la_oenb[31]
port 204 nsew signal input
rlabel metal2 s 187824 0 187880 400 6 la_oenb[32]
port 205 nsew signal input
rlabel metal2 s 190512 0 190568 400 6 la_oenb[33]
port 206 nsew signal input
rlabel metal2 s 193200 0 193256 400 6 la_oenb[34]
port 207 nsew signal input
rlabel metal2 s 195888 0 195944 400 6 la_oenb[35]
port 208 nsew signal input
rlabel metal2 s 198576 0 198632 400 6 la_oenb[36]
port 209 nsew signal input
rlabel metal2 s 201264 0 201320 400 6 la_oenb[37]
port 210 nsew signal input
rlabel metal2 s 203952 0 204008 400 6 la_oenb[38]
port 211 nsew signal input
rlabel metal2 s 206640 0 206696 400 6 la_oenb[39]
port 212 nsew signal input
rlabel metal2 s 109872 0 109928 400 6 la_oenb[3]
port 213 nsew signal input
rlabel metal2 s 209328 0 209384 400 6 la_oenb[40]
port 214 nsew signal input
rlabel metal2 s 212016 0 212072 400 6 la_oenb[41]
port 215 nsew signal input
rlabel metal2 s 214704 0 214760 400 6 la_oenb[42]
port 216 nsew signal input
rlabel metal2 s 217392 0 217448 400 6 la_oenb[43]
port 217 nsew signal input
rlabel metal2 s 220080 0 220136 400 6 la_oenb[44]
port 218 nsew signal input
rlabel metal2 s 222768 0 222824 400 6 la_oenb[45]
port 219 nsew signal input
rlabel metal2 s 225456 0 225512 400 6 la_oenb[46]
port 220 nsew signal input
rlabel metal2 s 228144 0 228200 400 6 la_oenb[47]
port 221 nsew signal input
rlabel metal2 s 230832 0 230888 400 6 la_oenb[48]
port 222 nsew signal input
rlabel metal2 s 233520 0 233576 400 6 la_oenb[49]
port 223 nsew signal input
rlabel metal2 s 112560 0 112616 400 6 la_oenb[4]
port 224 nsew signal input
rlabel metal2 s 236208 0 236264 400 6 la_oenb[50]
port 225 nsew signal input
rlabel metal2 s 238896 0 238952 400 6 la_oenb[51]
port 226 nsew signal input
rlabel metal2 s 241584 0 241640 400 6 la_oenb[52]
port 227 nsew signal input
rlabel metal2 s 244272 0 244328 400 6 la_oenb[53]
port 228 nsew signal input
rlabel metal2 s 246960 0 247016 400 6 la_oenb[54]
port 229 nsew signal input
rlabel metal2 s 249648 0 249704 400 6 la_oenb[55]
port 230 nsew signal input
rlabel metal2 s 252336 0 252392 400 6 la_oenb[56]
port 231 nsew signal input
rlabel metal2 s 255024 0 255080 400 6 la_oenb[57]
port 232 nsew signal input
rlabel metal2 s 257712 0 257768 400 6 la_oenb[58]
port 233 nsew signal input
rlabel metal2 s 260400 0 260456 400 6 la_oenb[59]
port 234 nsew signal input
rlabel metal2 s 115248 0 115304 400 6 la_oenb[5]
port 235 nsew signal input
rlabel metal2 s 263088 0 263144 400 6 la_oenb[60]
port 236 nsew signal input
rlabel metal2 s 265776 0 265832 400 6 la_oenb[61]
port 237 nsew signal input
rlabel metal2 s 268464 0 268520 400 6 la_oenb[62]
port 238 nsew signal input
rlabel metal2 s 271152 0 271208 400 6 la_oenb[63]
port 239 nsew signal input
rlabel metal2 s 117936 0 117992 400 6 la_oenb[6]
port 240 nsew signal input
rlabel metal2 s 120624 0 120680 400 6 la_oenb[7]
port 241 nsew signal input
rlabel metal2 s 123312 0 123368 400 6 la_oenb[8]
port 242 nsew signal input
rlabel metal2 s 126000 0 126056 400 6 la_oenb[9]
port 243 nsew signal input
rlabel metal2 s 274736 0 274792 400 6 user_clock2
port 244 nsew signal input
rlabel metal4 s 2224 1538 2384 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vdd
port 245 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vss
port 246 nsew ground bidirectional
rlabel metal2 s 5040 0 5096 400 6 wb_clk_i
port 247 nsew signal input
rlabel metal2 s 5936 0 5992 400 6 wb_rst_i
port 248 nsew signal input
rlabel metal2 s 6832 0 6888 400 6 wbs_ack_o
port 249 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 wbs_adr_i[0]
port 250 nsew signal input
rlabel metal2 s 40880 0 40936 400 6 wbs_adr_i[10]
port 251 nsew signal input
rlabel metal2 s 43568 0 43624 400 6 wbs_adr_i[11]
port 252 nsew signal input
rlabel metal2 s 46256 0 46312 400 6 wbs_adr_i[12]
port 253 nsew signal input
rlabel metal2 s 48944 0 49000 400 6 wbs_adr_i[13]
port 254 nsew signal input
rlabel metal2 s 51632 0 51688 400 6 wbs_adr_i[14]
port 255 nsew signal input
rlabel metal2 s 54320 0 54376 400 6 wbs_adr_i[15]
port 256 nsew signal input
rlabel metal2 s 57008 0 57064 400 6 wbs_adr_i[16]
port 257 nsew signal input
rlabel metal2 s 59696 0 59752 400 6 wbs_adr_i[17]
port 258 nsew signal input
rlabel metal2 s 62384 0 62440 400 6 wbs_adr_i[18]
port 259 nsew signal input
rlabel metal2 s 65072 0 65128 400 6 wbs_adr_i[19]
port 260 nsew signal input
rlabel metal2 s 14000 0 14056 400 6 wbs_adr_i[1]
port 261 nsew signal input
rlabel metal2 s 67760 0 67816 400 6 wbs_adr_i[20]
port 262 nsew signal input
rlabel metal2 s 70448 0 70504 400 6 wbs_adr_i[21]
port 263 nsew signal input
rlabel metal2 s 73136 0 73192 400 6 wbs_adr_i[22]
port 264 nsew signal input
rlabel metal2 s 75824 0 75880 400 6 wbs_adr_i[23]
port 265 nsew signal input
rlabel metal2 s 78512 0 78568 400 6 wbs_adr_i[24]
port 266 nsew signal input
rlabel metal2 s 81200 0 81256 400 6 wbs_adr_i[25]
port 267 nsew signal input
rlabel metal2 s 83888 0 83944 400 6 wbs_adr_i[26]
port 268 nsew signal input
rlabel metal2 s 86576 0 86632 400 6 wbs_adr_i[27]
port 269 nsew signal input
rlabel metal2 s 89264 0 89320 400 6 wbs_adr_i[28]
port 270 nsew signal input
rlabel metal2 s 91952 0 92008 400 6 wbs_adr_i[29]
port 271 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 wbs_adr_i[2]
port 272 nsew signal input
rlabel metal2 s 94640 0 94696 400 6 wbs_adr_i[30]
port 273 nsew signal input
rlabel metal2 s 97328 0 97384 400 6 wbs_adr_i[31]
port 274 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 wbs_adr_i[3]
port 275 nsew signal input
rlabel metal2 s 24752 0 24808 400 6 wbs_adr_i[4]
port 276 nsew signal input
rlabel metal2 s 27440 0 27496 400 6 wbs_adr_i[5]
port 277 nsew signal input
rlabel metal2 s 30128 0 30184 400 6 wbs_adr_i[6]
port 278 nsew signal input
rlabel metal2 s 32816 0 32872 400 6 wbs_adr_i[7]
port 279 nsew signal input
rlabel metal2 s 35504 0 35560 400 6 wbs_adr_i[8]
port 280 nsew signal input
rlabel metal2 s 38192 0 38248 400 6 wbs_adr_i[9]
port 281 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 wbs_cyc_i
port 282 nsew signal input
rlabel metal2 s 11312 0 11368 400 6 wbs_dat_i[0]
port 283 nsew signal input
rlabel metal2 s 41776 0 41832 400 6 wbs_dat_i[10]
port 284 nsew signal input
rlabel metal2 s 44464 0 44520 400 6 wbs_dat_i[11]
port 285 nsew signal input
rlabel metal2 s 47152 0 47208 400 6 wbs_dat_i[12]
port 286 nsew signal input
rlabel metal2 s 49840 0 49896 400 6 wbs_dat_i[13]
port 287 nsew signal input
rlabel metal2 s 52528 0 52584 400 6 wbs_dat_i[14]
port 288 nsew signal input
rlabel metal2 s 55216 0 55272 400 6 wbs_dat_i[15]
port 289 nsew signal input
rlabel metal2 s 57904 0 57960 400 6 wbs_dat_i[16]
port 290 nsew signal input
rlabel metal2 s 60592 0 60648 400 6 wbs_dat_i[17]
port 291 nsew signal input
rlabel metal2 s 63280 0 63336 400 6 wbs_dat_i[18]
port 292 nsew signal input
rlabel metal2 s 65968 0 66024 400 6 wbs_dat_i[19]
port 293 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 wbs_dat_i[1]
port 294 nsew signal input
rlabel metal2 s 68656 0 68712 400 6 wbs_dat_i[20]
port 295 nsew signal input
rlabel metal2 s 71344 0 71400 400 6 wbs_dat_i[21]
port 296 nsew signal input
rlabel metal2 s 74032 0 74088 400 6 wbs_dat_i[22]
port 297 nsew signal input
rlabel metal2 s 76720 0 76776 400 6 wbs_dat_i[23]
port 298 nsew signal input
rlabel metal2 s 79408 0 79464 400 6 wbs_dat_i[24]
port 299 nsew signal input
rlabel metal2 s 82096 0 82152 400 6 wbs_dat_i[25]
port 300 nsew signal input
rlabel metal2 s 84784 0 84840 400 6 wbs_dat_i[26]
port 301 nsew signal input
rlabel metal2 s 87472 0 87528 400 6 wbs_dat_i[27]
port 302 nsew signal input
rlabel metal2 s 90160 0 90216 400 6 wbs_dat_i[28]
port 303 nsew signal input
rlabel metal2 s 92848 0 92904 400 6 wbs_dat_i[29]
port 304 nsew signal input
rlabel metal2 s 18480 0 18536 400 6 wbs_dat_i[2]
port 305 nsew signal input
rlabel metal2 s 95536 0 95592 400 6 wbs_dat_i[30]
port 306 nsew signal input
rlabel metal2 s 98224 0 98280 400 6 wbs_dat_i[31]
port 307 nsew signal input
rlabel metal2 s 22064 0 22120 400 6 wbs_dat_i[3]
port 308 nsew signal input
rlabel metal2 s 25648 0 25704 400 6 wbs_dat_i[4]
port 309 nsew signal input
rlabel metal2 s 28336 0 28392 400 6 wbs_dat_i[5]
port 310 nsew signal input
rlabel metal2 s 31024 0 31080 400 6 wbs_dat_i[6]
port 311 nsew signal input
rlabel metal2 s 33712 0 33768 400 6 wbs_dat_i[7]
port 312 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 wbs_dat_i[8]
port 313 nsew signal input
rlabel metal2 s 39088 0 39144 400 6 wbs_dat_i[9]
port 314 nsew signal input
rlabel metal2 s 12208 0 12264 400 6 wbs_dat_o[0]
port 315 nsew signal output
rlabel metal2 s 42672 0 42728 400 6 wbs_dat_o[10]
port 316 nsew signal output
rlabel metal2 s 45360 0 45416 400 6 wbs_dat_o[11]
port 317 nsew signal output
rlabel metal2 s 48048 0 48104 400 6 wbs_dat_o[12]
port 318 nsew signal output
rlabel metal2 s 50736 0 50792 400 6 wbs_dat_o[13]
port 319 nsew signal output
rlabel metal2 s 53424 0 53480 400 6 wbs_dat_o[14]
port 320 nsew signal output
rlabel metal2 s 56112 0 56168 400 6 wbs_dat_o[15]
port 321 nsew signal output
rlabel metal2 s 58800 0 58856 400 6 wbs_dat_o[16]
port 322 nsew signal output
rlabel metal2 s 61488 0 61544 400 6 wbs_dat_o[17]
port 323 nsew signal output
rlabel metal2 s 64176 0 64232 400 6 wbs_dat_o[18]
port 324 nsew signal output
rlabel metal2 s 66864 0 66920 400 6 wbs_dat_o[19]
port 325 nsew signal output
rlabel metal2 s 15792 0 15848 400 6 wbs_dat_o[1]
port 326 nsew signal output
rlabel metal2 s 69552 0 69608 400 6 wbs_dat_o[20]
port 327 nsew signal output
rlabel metal2 s 72240 0 72296 400 6 wbs_dat_o[21]
port 328 nsew signal output
rlabel metal2 s 74928 0 74984 400 6 wbs_dat_o[22]
port 329 nsew signal output
rlabel metal2 s 77616 0 77672 400 6 wbs_dat_o[23]
port 330 nsew signal output
rlabel metal2 s 80304 0 80360 400 6 wbs_dat_o[24]
port 331 nsew signal output
rlabel metal2 s 82992 0 83048 400 6 wbs_dat_o[25]
port 332 nsew signal output
rlabel metal2 s 85680 0 85736 400 6 wbs_dat_o[26]
port 333 nsew signal output
rlabel metal2 s 88368 0 88424 400 6 wbs_dat_o[27]
port 334 nsew signal output
rlabel metal2 s 91056 0 91112 400 6 wbs_dat_o[28]
port 335 nsew signal output
rlabel metal2 s 93744 0 93800 400 6 wbs_dat_o[29]
port 336 nsew signal output
rlabel metal2 s 19376 0 19432 400 6 wbs_dat_o[2]
port 337 nsew signal output
rlabel metal2 s 96432 0 96488 400 6 wbs_dat_o[30]
port 338 nsew signal output
rlabel metal2 s 99120 0 99176 400 6 wbs_dat_o[31]
port 339 nsew signal output
rlabel metal2 s 22960 0 23016 400 6 wbs_dat_o[3]
port 340 nsew signal output
rlabel metal2 s 26544 0 26600 400 6 wbs_dat_o[4]
port 341 nsew signal output
rlabel metal2 s 29232 0 29288 400 6 wbs_dat_o[5]
port 342 nsew signal output
rlabel metal2 s 31920 0 31976 400 6 wbs_dat_o[6]
port 343 nsew signal output
rlabel metal2 s 34608 0 34664 400 6 wbs_dat_o[7]
port 344 nsew signal output
rlabel metal2 s 37296 0 37352 400 6 wbs_dat_o[8]
port 345 nsew signal output
rlabel metal2 s 39984 0 40040 400 6 wbs_dat_o[9]
port 346 nsew signal output
rlabel metal2 s 13104 0 13160 400 6 wbs_sel_i[0]
port 347 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 wbs_sel_i[1]
port 348 nsew signal input
rlabel metal2 s 20272 0 20328 400 6 wbs_sel_i[2]
port 349 nsew signal input
rlabel metal2 s 23856 0 23912 400 6 wbs_sel_i[3]
port 350 nsew signal input
rlabel metal2 s 8624 0 8680 400 6 wbs_stb_i
port 351 nsew signal input
rlabel metal2 s 9520 0 9576 400 6 wbs_we_i
port 352 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 42159254
string GDS_FILE /home/thomas/Documents/Projects/tilerisc/openlane/tjrpu/runs/23_12_11_07_45/results/signoff/tjrpu.magic.gds
string GDS_START 519380
<< end >>

