VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tinyrv
  CLASS BLOCK ;
  FOREIGN tinyrv ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 15.680 0.000 16.240 4.000 ;
    END
  END clk
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END inst[0]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 4.000 ;
    END
  END inst[10]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 0.000 137.200 4.000 ;
    END
  END inst[11]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 0.000 147.280 4.000 ;
    END
  END inst[12]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 0.000 157.360 4.000 ;
    END
  END inst[13]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END inst[14]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 0.000 177.520 4.000 ;
    END
  END inst[15]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 4.000 ;
    END
  END inst[16]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 0.000 197.680 4.000 ;
    END
  END inst[17]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 0.000 207.760 4.000 ;
    END
  END inst[18]
  PIN inst[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 0.000 217.840 4.000 ;
    END
  END inst[19]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 0.000 36.400 4.000 ;
    END
  END inst[1]
  PIN inst[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 0.000 227.920 4.000 ;
    END
  END inst[20]
  PIN inst[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 0.000 238.000 4.000 ;
    END
  END inst[21]
  PIN inst[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 0.000 248.080 4.000 ;
    END
  END inst[22]
  PIN inst[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 0.000 258.160 4.000 ;
    END
  END inst[23]
  PIN inst[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 0.000 268.240 4.000 ;
    END
  END inst[24]
  PIN inst[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 0.000 278.320 4.000 ;
    END
  END inst[25]
  PIN inst[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 0.000 288.400 4.000 ;
    END
  END inst[26]
  PIN inst[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 0.000 298.480 4.000 ;
    END
  END inst[27]
  PIN inst[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 0.000 308.560 4.000 ;
    END
  END inst[28]
  PIN inst[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 318.080 0.000 318.640 4.000 ;
    END
  END inst[29]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 4.000 ;
    END
  END inst[2]
  PIN inst[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 0.000 328.720 4.000 ;
    END
  END inst[30]
  PIN inst[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 0.000 338.800 4.000 ;
    END
  END inst[31]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 4.000 ;
    END
  END inst[3]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 4.000 ;
    END
  END inst[4]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 0.000 76.720 4.000 ;
    END
  END inst[5]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 4.000 ;
    END
  END inst[6]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 0.000 96.880 4.000 ;
    END
  END inst[7]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 4.000 ;
    END
  END inst[8]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 4.000 ;
    END
  END inst[9]
  PIN mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 969.920 996.000 970.480 1000.000 ;
    END
  END mem_addr[0]
  PIN mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 880.320 996.000 880.880 1000.000 ;
    END
  END mem_addr[10]
  PIN mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 871.360 996.000 871.920 1000.000 ;
    END
  END mem_addr[11]
  PIN mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 996.000 862.960 1000.000 ;
    END
  END mem_addr[12]
  PIN mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 853.440 996.000 854.000 1000.000 ;
    END
  END mem_addr[13]
  PIN mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 844.480 996.000 845.040 1000.000 ;
    END
  END mem_addr[14]
  PIN mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 835.520 996.000 836.080 1000.000 ;
    END
  END mem_addr[15]
  PIN mem_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 826.560 996.000 827.120 1000.000 ;
    END
  END mem_addr[16]
  PIN mem_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 817.600 996.000 818.160 1000.000 ;
    END
  END mem_addr[17]
  PIN mem_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 808.640 996.000 809.200 1000.000 ;
    END
  END mem_addr[18]
  PIN mem_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 996.000 800.240 1000.000 ;
    END
  END mem_addr[19]
  PIN mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 960.960 996.000 961.520 1000.000 ;
    END
  END mem_addr[1]
  PIN mem_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 790.720 996.000 791.280 1000.000 ;
    END
  END mem_addr[20]
  PIN mem_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 781.760 996.000 782.320 1000.000 ;
    END
  END mem_addr[21]
  PIN mem_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 996.000 773.360 1000.000 ;
    END
  END mem_addr[22]
  PIN mem_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 763.840 996.000 764.400 1000.000 ;
    END
  END mem_addr[23]
  PIN mem_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 754.880 996.000 755.440 1000.000 ;
    END
  END mem_addr[24]
  PIN mem_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 996.000 746.480 1000.000 ;
    END
  END mem_addr[25]
  PIN mem_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 736.960 996.000 737.520 1000.000 ;
    END
  END mem_addr[26]
  PIN mem_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 728.000 996.000 728.560 1000.000 ;
    END
  END mem_addr[27]
  PIN mem_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 996.000 719.600 1000.000 ;
    END
  END mem_addr[28]
  PIN mem_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 710.080 996.000 710.640 1000.000 ;
    END
  END mem_addr[29]
  PIN mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 952.000 996.000 952.560 1000.000 ;
    END
  END mem_addr[2]
  PIN mem_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 701.120 996.000 701.680 1000.000 ;
    END
  END mem_addr[30]
  PIN mem_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 996.000 692.720 1000.000 ;
    END
  END mem_addr[31]
  PIN mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 943.040 996.000 943.600 1000.000 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 934.080 996.000 934.640 1000.000 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 925.120 996.000 925.680 1000.000 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 916.160 996.000 916.720 1000.000 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 996.000 907.760 1000.000 ;
    END
  END mem_addr[7]
  PIN mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 898.240 996.000 898.800 1000.000 ;
    END
  END mem_addr[8]
  PIN mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 889.280 996.000 889.840 1000.000 ;
    END
  END mem_addr[9]
  PIN mem_ld_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 996.000 638.960 1000.000 ;
    END
  END mem_ld_dat[0]
  PIN mem_ld_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 996.000 549.360 1000.000 ;
    END
  END mem_ld_dat[10]
  PIN mem_ld_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 996.000 540.400 1000.000 ;
    END
  END mem_ld_dat[11]
  PIN mem_ld_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 996.000 531.440 1000.000 ;
    END
  END mem_ld_dat[12]
  PIN mem_ld_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 521.920 996.000 522.480 1000.000 ;
    END
  END mem_ld_dat[13]
  PIN mem_ld_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 512.960 996.000 513.520 1000.000 ;
    END
  END mem_ld_dat[14]
  PIN mem_ld_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 996.000 504.560 1000.000 ;
    END
  END mem_ld_dat[15]
  PIN mem_ld_dat[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 495.040 996.000 495.600 1000.000 ;
    END
  END mem_ld_dat[16]
  PIN mem_ld_dat[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 486.080 996.000 486.640 1000.000 ;
    END
  END mem_ld_dat[17]
  PIN mem_ld_dat[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 996.000 477.680 1000.000 ;
    END
  END mem_ld_dat[18]
  PIN mem_ld_dat[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 468.160 996.000 468.720 1000.000 ;
    END
  END mem_ld_dat[19]
  PIN mem_ld_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 629.440 996.000 630.000 1000.000 ;
    END
  END mem_ld_dat[1]
  PIN mem_ld_dat[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 996.000 459.760 1000.000 ;
    END
  END mem_ld_dat[20]
  PIN mem_ld_dat[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 996.000 450.800 1000.000 ;
    END
  END mem_ld_dat[21]
  PIN mem_ld_dat[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 996.000 441.840 1000.000 ;
    END
  END mem_ld_dat[22]
  PIN mem_ld_dat[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 996.000 432.880 1000.000 ;
    END
  END mem_ld_dat[23]
  PIN mem_ld_dat[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 996.000 423.920 1000.000 ;
    END
  END mem_ld_dat[24]
  PIN mem_ld_dat[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 996.000 414.960 1000.000 ;
    END
  END mem_ld_dat[25]
  PIN mem_ld_dat[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 405.440 996.000 406.000 1000.000 ;
    END
  END mem_ld_dat[26]
  PIN mem_ld_dat[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 996.000 397.040 1000.000 ;
    END
  END mem_ld_dat[27]
  PIN mem_ld_dat[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 996.000 388.080 1000.000 ;
    END
  END mem_ld_dat[28]
  PIN mem_ld_dat[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 996.000 379.120 1000.000 ;
    END
  END mem_ld_dat[29]
  PIN mem_ld_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 620.480 996.000 621.040 1000.000 ;
    END
  END mem_ld_dat[2]
  PIN mem_ld_dat[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 996.000 370.160 1000.000 ;
    END
  END mem_ld_dat[30]
  PIN mem_ld_dat[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 996.000 361.200 1000.000 ;
    END
  END mem_ld_dat[31]
  PIN mem_ld_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 996.000 612.080 1000.000 ;
    END
  END mem_ld_dat[3]
  PIN mem_ld_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 602.560 996.000 603.120 1000.000 ;
    END
  END mem_ld_dat[4]
  PIN mem_ld_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 593.600 996.000 594.160 1000.000 ;
    END
  END mem_ld_dat[5]
  PIN mem_ld_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 996.000 585.200 1000.000 ;
    END
  END mem_ld_dat[6]
  PIN mem_ld_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 996.000 576.240 1000.000 ;
    END
  END mem_ld_dat[7]
  PIN mem_ld_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 566.720 996.000 567.280 1000.000 ;
    END
  END mem_ld_dat[8]
  PIN mem_ld_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 996.000 558.320 1000.000 ;
    END
  END mem_ld_dat[9]
  PIN mem_ld_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 683.200 996.000 683.760 1000.000 ;
    END
  END mem_ld_en
  PIN mem_ld_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 674.240 996.000 674.800 1000.000 ;
    END
  END mem_ld_mask[0]
  PIN mem_ld_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 996.000 665.840 1000.000 ;
    END
  END mem_ld_mask[1]
  PIN mem_ld_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 656.320 996.000 656.880 1000.000 ;
    END
  END mem_ld_mask[2]
  PIN mem_ld_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 647.360 996.000 647.920 1000.000 ;
    END
  END mem_ld_mask[3]
  PIN mem_st_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 996.000 307.440 1000.000 ;
    END
  END mem_st_dat[0]
  PIN mem_st_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 996.000 217.840 1000.000 ;
    END
  END mem_st_dat[10]
  PIN mem_st_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 996.000 208.880 1000.000 ;
    END
  END mem_st_dat[11]
  PIN mem_st_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 996.000 199.920 1000.000 ;
    END
  END mem_st_dat[12]
  PIN mem_st_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 996.000 190.960 1000.000 ;
    END
  END mem_st_dat[13]
  PIN mem_st_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 996.000 182.000 1000.000 ;
    END
  END mem_st_dat[14]
  PIN mem_st_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 996.000 173.040 1000.000 ;
    END
  END mem_st_dat[15]
  PIN mem_st_dat[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 996.000 164.080 1000.000 ;
    END
  END mem_st_dat[16]
  PIN mem_st_dat[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 996.000 155.120 1000.000 ;
    END
  END mem_st_dat[17]
  PIN mem_st_dat[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 996.000 146.160 1000.000 ;
    END
  END mem_st_dat[18]
  PIN mem_st_dat[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 996.000 137.200 1000.000 ;
    END
  END mem_st_dat[19]
  PIN mem_st_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 996.000 298.480 1000.000 ;
    END
  END mem_st_dat[1]
  PIN mem_st_dat[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 996.000 128.240 1000.000 ;
    END
  END mem_st_dat[20]
  PIN mem_st_dat[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 996.000 119.280 1000.000 ;
    END
  END mem_st_dat[21]
  PIN mem_st_dat[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 996.000 110.320 1000.000 ;
    END
  END mem_st_dat[22]
  PIN mem_st_dat[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 996.000 101.360 1000.000 ;
    END
  END mem_st_dat[23]
  PIN mem_st_dat[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 996.000 92.400 1000.000 ;
    END
  END mem_st_dat[24]
  PIN mem_st_dat[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 996.000 83.440 1000.000 ;
    END
  END mem_st_dat[25]
  PIN mem_st_dat[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 996.000 74.480 1000.000 ;
    END
  END mem_st_dat[26]
  PIN mem_st_dat[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 996.000 65.520 1000.000 ;
    END
  END mem_st_dat[27]
  PIN mem_st_dat[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 996.000 56.560 1000.000 ;
    END
  END mem_st_dat[28]
  PIN mem_st_dat[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 996.000 47.600 1000.000 ;
    END
  END mem_st_dat[29]
  PIN mem_st_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 996.000 289.520 1000.000 ;
    END
  END mem_st_dat[2]
  PIN mem_st_dat[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 996.000 38.640 1000.000 ;
    END
  END mem_st_dat[30]
  PIN mem_st_dat[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 996.000 29.680 1000.000 ;
    END
  END mem_st_dat[31]
  PIN mem_st_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 996.000 280.560 1000.000 ;
    END
  END mem_st_dat[3]
  PIN mem_st_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 996.000 271.600 1000.000 ;
    END
  END mem_st_dat[4]
  PIN mem_st_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 996.000 262.640 1000.000 ;
    END
  END mem_st_dat[5]
  PIN mem_st_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 996.000 253.680 1000.000 ;
    END
  END mem_st_dat[6]
  PIN mem_st_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 996.000 244.720 1000.000 ;
    END
  END mem_st_dat[7]
  PIN mem_st_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 996.000 235.760 1000.000 ;
    END
  END mem_st_dat[8]
  PIN mem_st_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 996.000 226.800 1000.000 ;
    END
  END mem_st_dat[9]
  PIN mem_st_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 996.000 352.240 1000.000 ;
    END
  END mem_st_en
  PIN mem_st_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 996.000 343.280 1000.000 ;
    END
  END mem_st_mask[0]
  PIN mem_st_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 996.000 334.320 1000.000 ;
    END
  END mem_st_mask[1]
  PIN mem_st_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 996.000 325.360 1000.000 ;
    END
  END mem_st_mask[2]
  PIN mem_st_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 996.000 316.400 1000.000 ;
    END
  END mem_st_mask[3]
  PIN pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 0.000 348.880 4.000 ;
    END
  END pc[0]
  PIN pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 0.000 449.680 4.000 ;
    END
  END pc[10]
  PIN pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 0.000 459.760 4.000 ;
    END
  END pc[11]
  PIN pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 0.000 469.840 4.000 ;
    END
  END pc[12]
  PIN pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 479.360 0.000 479.920 4.000 ;
    END
  END pc[13]
  PIN pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 489.440 0.000 490.000 4.000 ;
    END
  END pc[14]
  PIN pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 0.000 500.080 4.000 ;
    END
  END pc[15]
  PIN pc[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 509.600 0.000 510.160 4.000 ;
    END
  END pc[16]
  PIN pc[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 519.680 0.000 520.240 4.000 ;
    END
  END pc[17]
  PIN pc[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 0.000 530.320 4.000 ;
    END
  END pc[18]
  PIN pc[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 0.000 540.400 4.000 ;
    END
  END pc[19]
  PIN pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 358.400 0.000 358.960 4.000 ;
    END
  END pc[1]
  PIN pc[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 549.920 0.000 550.480 4.000 ;
    END
  END pc[20]
  PIN pc[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 560.000 0.000 560.560 4.000 ;
    END
  END pc[21]
  PIN pc[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 570.080 0.000 570.640 4.000 ;
    END
  END pc[22]
  PIN pc[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 0.000 580.720 4.000 ;
    END
  END pc[23]
  PIN pc[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 0.000 590.800 4.000 ;
    END
  END pc[24]
  PIN pc[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 600.320 0.000 600.880 4.000 ;
    END
  END pc[25]
  PIN pc[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 610.400 0.000 610.960 4.000 ;
    END
  END pc[26]
  PIN pc[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 620.480 0.000 621.040 4.000 ;
    END
  END pc[27]
  PIN pc[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 630.560 0.000 631.120 4.000 ;
    END
  END pc[28]
  PIN pc[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 640.640 0.000 641.200 4.000 ;
    END
  END pc[29]
  PIN pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 368.480 0.000 369.040 4.000 ;
    END
  END pc[2]
  PIN pc[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 650.720 0.000 651.280 4.000 ;
    END
  END pc[30]
  PIN pc[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 660.800 0.000 661.360 4.000 ;
    END
  END pc[31]
  PIN pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 0.000 379.120 4.000 ;
    END
  END pc[3]
  PIN pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 388.640 0.000 389.200 4.000 ;
    END
  END pc[4]
  PIN pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 398.720 0.000 399.280 4.000 ;
    END
  END pc[5]
  PIN pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 0.000 409.360 4.000 ;
    END
  END pc[6]
  PIN pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 0.000 419.440 4.000 ;
    END
  END pc[7]
  PIN pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 428.960 0.000 429.520 4.000 ;
    END
  END pc[8]
  PIN pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 439.040 0.000 439.600 4.000 ;
    END
  END pc[9]
  PIN pc_next[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 670.880 0.000 671.440 4.000 ;
    END
  END pc_next[0]
  PIN pc_next[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 771.680 0.000 772.240 4.000 ;
    END
  END pc_next[10]
  PIN pc_next[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 781.760 0.000 782.320 4.000 ;
    END
  END pc_next[11]
  PIN pc_next[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 791.840 0.000 792.400 4.000 ;
    END
  END pc_next[12]
  PIN pc_next[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 801.920 0.000 802.480 4.000 ;
    END
  END pc_next[13]
  PIN pc_next[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 812.000 0.000 812.560 4.000 ;
    END
  END pc_next[14]
  PIN pc_next[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 822.080 0.000 822.640 4.000 ;
    END
  END pc_next[15]
  PIN pc_next[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 832.160 0.000 832.720 4.000 ;
    END
  END pc_next[16]
  PIN pc_next[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 842.240 0.000 842.800 4.000 ;
    END
  END pc_next[17]
  PIN pc_next[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 852.320 0.000 852.880 4.000 ;
    END
  END pc_next[18]
  PIN pc_next[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 0.000 862.960 4.000 ;
    END
  END pc_next[19]
  PIN pc_next[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 680.960 0.000 681.520 4.000 ;
    END
  END pc_next[1]
  PIN pc_next[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 872.480 0.000 873.040 4.000 ;
    END
  END pc_next[20]
  PIN pc_next[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 882.560 0.000 883.120 4.000 ;
    END
  END pc_next[21]
  PIN pc_next[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 892.640 0.000 893.200 4.000 ;
    END
  END pc_next[22]
  PIN pc_next[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 902.720 0.000 903.280 4.000 ;
    END
  END pc_next[23]
  PIN pc_next[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 912.800 0.000 913.360 4.000 ;
    END
  END pc_next[24]
  PIN pc_next[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 922.880 0.000 923.440 4.000 ;
    END
  END pc_next[25]
  PIN pc_next[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 932.960 0.000 933.520 4.000 ;
    END
  END pc_next[26]
  PIN pc_next[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 943.040 0.000 943.600 4.000 ;
    END
  END pc_next[27]
  PIN pc_next[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 953.120 0.000 953.680 4.000 ;
    END
  END pc_next[28]
  PIN pc_next[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 963.200 0.000 963.760 4.000 ;
    END
  END pc_next[29]
  PIN pc_next[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 691.040 0.000 691.600 4.000 ;
    END
  END pc_next[2]
  PIN pc_next[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 973.280 0.000 973.840 4.000 ;
    END
  END pc_next[30]
  PIN pc_next[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 983.360 0.000 983.920 4.000 ;
    END
  END pc_next[31]
  PIN pc_next[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 701.120 0.000 701.680 4.000 ;
    END
  END pc_next[3]
  PIN pc_next[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 711.200 0.000 711.760 4.000 ;
    END
  END pc_next[4]
  PIN pc_next[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 721.280 0.000 721.840 4.000 ;
    END
  END pc_next[5]
  PIN pc_next[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 731.360 0.000 731.920 4.000 ;
    END
  END pc_next[6]
  PIN pc_next[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 741.440 0.000 742.000 4.000 ;
    END
  END pc_next[7]
  PIN pc_next[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 751.520 0.000 752.080 4.000 ;
    END
  END pc_next[8]
  PIN pc_next[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 761.600 0.000 762.160 4.000 ;
    END
  END pc_next[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 984.220 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 984.220 ;
    END
  END vss
  OBS
      LAYER Nwell ;
        RECT 6.290 981.885 993.310 984.350 ;
        RECT 6.290 981.760 391.980 981.885 ;
      LAYER Pwell ;
        RECT 6.290 978.240 993.310 981.760 ;
      LAYER Nwell ;
        RECT 6.290 978.115 294.945 978.240 ;
        RECT 6.290 974.045 993.310 978.115 ;
        RECT 6.290 973.920 348.145 974.045 ;
      LAYER Pwell ;
        RECT 6.290 970.400 993.310 973.920 ;
      LAYER Nwell ;
        RECT 6.290 970.275 230.545 970.400 ;
        RECT 6.290 966.205 993.310 970.275 ;
        RECT 6.290 966.080 171.745 966.205 ;
      LAYER Pwell ;
        RECT 6.290 962.560 993.310 966.080 ;
      LAYER Nwell ;
        RECT 6.290 962.435 338.625 962.560 ;
        RECT 6.290 958.365 993.310 962.435 ;
        RECT 6.290 958.240 196.945 958.365 ;
      LAYER Pwell ;
        RECT 6.290 954.720 993.310 958.240 ;
      LAYER Nwell ;
        RECT 6.290 954.595 227.185 954.720 ;
        RECT 6.290 950.525 993.310 954.595 ;
        RECT 6.290 950.400 281.505 950.525 ;
      LAYER Pwell ;
        RECT 6.290 946.880 993.310 950.400 ;
      LAYER Nwell ;
        RECT 6.290 946.755 155.720 946.880 ;
        RECT 6.290 942.685 993.310 946.755 ;
        RECT 6.290 942.560 166.705 942.685 ;
      LAYER Pwell ;
        RECT 6.290 939.040 993.310 942.560 ;
      LAYER Nwell ;
        RECT 6.290 938.915 152.145 939.040 ;
        RECT 6.290 934.845 993.310 938.915 ;
        RECT 6.290 934.720 198.065 934.845 ;
      LAYER Pwell ;
        RECT 6.290 931.200 993.310 934.720 ;
      LAYER Nwell ;
        RECT 6.290 931.075 221.585 931.200 ;
        RECT 6.290 927.005 993.310 931.075 ;
        RECT 6.290 926.880 359.345 927.005 ;
      LAYER Pwell ;
        RECT 6.290 923.360 993.310 926.880 ;
      LAYER Nwell ;
        RECT 6.290 923.235 137.585 923.360 ;
        RECT 6.290 919.165 993.310 923.235 ;
        RECT 6.290 919.040 328.545 919.165 ;
      LAYER Pwell ;
        RECT 6.290 915.520 993.310 919.040 ;
      LAYER Nwell ;
        RECT 6.290 915.395 135.905 915.520 ;
        RECT 6.290 911.325 993.310 915.395 ;
        RECT 6.290 911.200 274.225 911.325 ;
      LAYER Pwell ;
        RECT 6.290 907.680 993.310 911.200 ;
      LAYER Nwell ;
        RECT 6.290 907.555 218.785 907.680 ;
        RECT 6.290 903.485 993.310 907.555 ;
        RECT 6.290 903.360 119.105 903.485 ;
      LAYER Pwell ;
        RECT 6.290 899.840 993.310 903.360 ;
      LAYER Nwell ;
        RECT 6.290 899.715 191.345 899.840 ;
        RECT 6.290 895.645 993.310 899.715 ;
        RECT 6.290 895.520 123.025 895.645 ;
      LAYER Pwell ;
        RECT 6.290 892.000 993.310 895.520 ;
      LAYER Nwell ;
        RECT 6.290 891.875 248.465 892.000 ;
        RECT 6.290 887.805 993.310 891.875 ;
        RECT 6.290 887.680 435.720 887.805 ;
      LAYER Pwell ;
        RECT 6.290 884.160 993.310 887.680 ;
      LAYER Nwell ;
        RECT 6.290 884.035 218.785 884.160 ;
        RECT 6.290 879.965 993.310 884.035 ;
        RECT 6.290 879.840 327.985 879.965 ;
      LAYER Pwell ;
        RECT 6.290 876.320 993.310 879.840 ;
      LAYER Nwell ;
        RECT 6.290 876.195 112.945 876.320 ;
        RECT 6.290 872.125 993.310 876.195 ;
        RECT 6.290 872.000 110.705 872.125 ;
      LAYER Pwell ;
        RECT 6.290 868.480 993.310 872.000 ;
      LAYER Nwell ;
        RECT 6.290 868.355 450.625 868.480 ;
        RECT 6.290 864.285 993.310 868.355 ;
        RECT 6.290 864.160 482.545 864.285 ;
      LAYER Pwell ;
        RECT 6.290 860.640 993.310 864.160 ;
      LAYER Nwell ;
        RECT 6.290 860.515 185.745 860.640 ;
        RECT 6.290 856.445 993.310 860.515 ;
        RECT 6.290 856.320 210.600 856.445 ;
      LAYER Pwell ;
        RECT 6.290 852.800 993.310 856.320 ;
      LAYER Nwell ;
        RECT 6.290 852.675 91.105 852.800 ;
        RECT 6.290 848.605 993.310 852.675 ;
        RECT 6.290 848.480 112.385 848.605 ;
      LAYER Pwell ;
        RECT 6.290 844.960 993.310 848.480 ;
      LAYER Nwell ;
        RECT 6.290 844.835 144.305 844.960 ;
        RECT 6.290 840.765 993.310 844.835 ;
        RECT 6.290 840.640 83.825 840.765 ;
      LAYER Pwell ;
        RECT 6.290 837.120 993.310 840.640 ;
      LAYER Nwell ;
        RECT 6.290 836.995 60.865 837.120 ;
        RECT 6.290 832.925 993.310 836.995 ;
        RECT 6.290 832.800 54.145 832.925 ;
      LAYER Pwell ;
        RECT 6.290 829.280 993.310 832.800 ;
      LAYER Nwell ;
        RECT 6.290 829.155 374.465 829.280 ;
        RECT 6.290 825.085 993.310 829.155 ;
        RECT 6.290 824.960 79.345 825.085 ;
      LAYER Pwell ;
        RECT 6.290 821.440 993.310 824.960 ;
      LAYER Nwell ;
        RECT 6.290 821.315 110.705 821.440 ;
        RECT 6.290 817.245 993.310 821.315 ;
        RECT 6.290 817.120 110.705 817.245 ;
      LAYER Pwell ;
        RECT 6.290 813.600 993.310 817.120 ;
      LAYER Nwell ;
        RECT 6.290 813.475 51.905 813.600 ;
        RECT 6.290 809.405 993.310 813.475 ;
        RECT 6.290 809.280 45.745 809.405 ;
      LAYER Pwell ;
        RECT 6.290 805.760 993.310 809.280 ;
      LAYER Nwell ;
        RECT 6.290 805.635 22.785 805.760 ;
        RECT 6.290 801.565 993.310 805.635 ;
        RECT 6.290 801.440 139.305 801.565 ;
      LAYER Pwell ;
        RECT 6.290 797.920 993.310 801.440 ;
      LAYER Nwell ;
        RECT 6.290 797.795 24.465 797.920 ;
        RECT 6.290 793.725 993.310 797.795 ;
        RECT 6.290 793.600 14.945 793.725 ;
      LAYER Pwell ;
        RECT 6.290 790.080 993.310 793.600 ;
      LAYER Nwell ;
        RECT 6.290 789.955 104.545 790.080 ;
        RECT 6.290 785.885 993.310 789.955 ;
        RECT 6.290 785.760 134.915 785.885 ;
      LAYER Pwell ;
        RECT 6.290 782.240 993.310 785.760 ;
      LAYER Nwell ;
        RECT 6.290 782.115 100.840 782.240 ;
        RECT 6.290 778.045 993.310 782.115 ;
        RECT 6.290 777.920 134.915 778.045 ;
      LAYER Pwell ;
        RECT 6.290 774.400 993.310 777.920 ;
      LAYER Nwell ;
        RECT 6.290 774.275 18.305 774.400 ;
        RECT 6.290 770.205 993.310 774.275 ;
        RECT 6.290 770.080 14.945 770.205 ;
      LAYER Pwell ;
        RECT 6.290 766.560 993.310 770.080 ;
      LAYER Nwell ;
        RECT 6.290 766.435 340.305 766.560 ;
        RECT 6.290 762.365 993.310 766.435 ;
        RECT 6.290 762.240 170.625 762.365 ;
      LAYER Pwell ;
        RECT 6.290 758.720 993.310 762.240 ;
      LAYER Nwell ;
        RECT 6.290 758.595 109.585 758.720 ;
        RECT 6.290 754.525 993.310 758.595 ;
        RECT 6.290 754.400 87.745 754.525 ;
      LAYER Pwell ;
        RECT 6.290 750.880 993.310 754.400 ;
      LAYER Nwell ;
        RECT 6.290 750.755 16.065 750.880 ;
        RECT 6.290 746.685 993.310 750.755 ;
        RECT 6.290 746.560 47.425 746.685 ;
      LAYER Pwell ;
        RECT 6.290 743.040 993.310 746.560 ;
      LAYER Nwell ;
        RECT 6.290 742.915 16.065 743.040 ;
        RECT 6.290 738.845 993.310 742.915 ;
        RECT 6.290 738.720 189.105 738.845 ;
      LAYER Pwell ;
        RECT 6.290 735.200 993.310 738.720 ;
      LAYER Nwell ;
        RECT 6.290 735.075 103.985 735.200 ;
        RECT 6.290 731.005 993.310 735.075 ;
        RECT 6.290 730.880 718.635 731.005 ;
      LAYER Pwell ;
        RECT 6.290 727.360 993.310 730.880 ;
      LAYER Nwell ;
        RECT 6.290 727.235 298.965 727.360 ;
        RECT 6.290 723.165 993.310 727.235 ;
        RECT 6.290 723.040 14.945 723.165 ;
      LAYER Pwell ;
        RECT 6.290 719.520 993.310 723.040 ;
      LAYER Nwell ;
        RECT 6.290 719.395 17.185 719.520 ;
        RECT 6.290 715.325 993.310 719.395 ;
        RECT 6.290 715.200 117.985 715.325 ;
      LAYER Pwell ;
        RECT 6.290 711.680 993.310 715.200 ;
      LAYER Nwell ;
        RECT 6.290 711.555 305.675 711.680 ;
        RECT 6.290 707.485 993.310 711.555 ;
        RECT 6.290 707.360 312.405 707.485 ;
      LAYER Pwell ;
        RECT 6.290 703.840 993.310 707.360 ;
      LAYER Nwell ;
        RECT 6.290 703.715 106.785 703.840 ;
        RECT 6.290 699.645 993.310 703.715 ;
        RECT 6.290 699.520 54.145 699.645 ;
      LAYER Pwell ;
        RECT 6.290 696.000 993.310 699.520 ;
      LAYER Nwell ;
        RECT 6.290 695.875 18.865 696.000 ;
        RECT 6.290 691.805 993.310 695.875 ;
        RECT 6.290 691.680 14.945 691.805 ;
      LAYER Pwell ;
        RECT 6.290 688.160 993.310 691.680 ;
      LAYER Nwell ;
        RECT 6.290 688.035 226.850 688.160 ;
        RECT 6.290 683.965 993.310 688.035 ;
        RECT 6.290 683.840 84.040 683.965 ;
      LAYER Pwell ;
        RECT 6.290 680.320 993.310 683.840 ;
      LAYER Nwell ;
        RECT 6.290 680.195 16.065 680.320 ;
        RECT 6.290 676.125 993.310 680.195 ;
        RECT 6.290 676.000 197.160 676.125 ;
      LAYER Pwell ;
        RECT 6.290 672.480 993.310 676.000 ;
      LAYER Nwell ;
        RECT 6.290 672.355 51.905 672.480 ;
        RECT 6.290 668.285 993.310 672.355 ;
        RECT 6.290 668.160 46.305 668.285 ;
      LAYER Pwell ;
        RECT 6.290 664.640 993.310 668.160 ;
      LAYER Nwell ;
        RECT 6.290 664.515 19.425 664.640 ;
        RECT 6.290 660.445 993.310 664.515 ;
        RECT 6.290 660.320 202.545 660.445 ;
      LAYER Pwell ;
        RECT 6.290 656.800 993.310 660.320 ;
      LAYER Nwell ;
        RECT 6.290 656.675 21.665 656.800 ;
        RECT 6.290 652.605 993.310 656.675 ;
        RECT 6.290 652.480 14.945 652.605 ;
      LAYER Pwell ;
        RECT 6.290 648.960 993.310 652.480 ;
      LAYER Nwell ;
        RECT 6.290 648.835 547.830 648.960 ;
        RECT 6.290 644.765 993.310 648.835 ;
        RECT 6.290 644.640 189.105 644.765 ;
      LAYER Pwell ;
        RECT 6.290 641.120 993.310 644.640 ;
      LAYER Nwell ;
        RECT 6.290 640.995 107.905 641.120 ;
        RECT 6.290 636.925 993.310 640.995 ;
        RECT 6.290 636.800 49.105 636.925 ;
      LAYER Pwell ;
        RECT 6.290 633.280 993.310 636.800 ;
      LAYER Nwell ;
        RECT 6.290 633.155 24.465 633.280 ;
        RECT 6.290 629.085 993.310 633.155 ;
        RECT 6.290 628.960 14.945 629.085 ;
      LAYER Pwell ;
        RECT 6.290 625.440 993.310 628.960 ;
      LAYER Nwell ;
        RECT 6.290 625.315 187.985 625.440 ;
        RECT 6.290 621.245 993.310 625.315 ;
        RECT 6.290 621.120 171.185 621.245 ;
      LAYER Pwell ;
        RECT 6.290 617.600 993.310 621.120 ;
      LAYER Nwell ;
        RECT 6.290 617.475 97.265 617.600 ;
        RECT 6.290 613.405 993.310 617.475 ;
        RECT 6.290 613.280 43.505 613.405 ;
      LAYER Pwell ;
        RECT 6.290 609.760 993.310 613.280 ;
      LAYER Nwell ;
        RECT 6.290 609.635 16.625 609.760 ;
        RECT 6.290 605.565 993.310 609.635 ;
        RECT 6.290 605.440 14.945 605.565 ;
      LAYER Pwell ;
        RECT 6.290 601.920 993.310 605.440 ;
      LAYER Nwell ;
        RECT 6.290 601.795 19.985 601.920 ;
        RECT 6.290 597.725 993.310 601.795 ;
        RECT 6.290 597.600 113.685 597.725 ;
      LAYER Pwell ;
        RECT 6.290 594.080 993.310 597.600 ;
      LAYER Nwell ;
        RECT 6.290 593.955 61.425 594.080 ;
        RECT 6.290 589.885 993.310 593.955 ;
        RECT 6.290 589.760 189.105 589.885 ;
      LAYER Pwell ;
        RECT 6.290 586.240 993.310 589.760 ;
      LAYER Nwell ;
        RECT 6.290 586.115 152.145 586.240 ;
        RECT 6.290 582.045 993.310 586.115 ;
        RECT 6.290 581.920 91.105 582.045 ;
      LAYER Pwell ;
        RECT 6.290 578.400 993.310 581.920 ;
      LAYER Nwell ;
        RECT 6.290 578.275 51.905 578.400 ;
        RECT 6.290 574.205 993.310 578.275 ;
        RECT 6.290 574.080 14.385 574.205 ;
      LAYER Pwell ;
        RECT 6.290 570.560 993.310 574.080 ;
      LAYER Nwell ;
        RECT 6.290 570.435 14.945 570.560 ;
        RECT 6.290 566.365 993.310 570.435 ;
        RECT 6.290 566.240 39.025 566.365 ;
      LAYER Pwell ;
        RECT 6.290 562.720 993.310 566.240 ;
      LAYER Nwell ;
        RECT 6.290 562.595 152.145 562.720 ;
        RECT 6.290 558.525 993.310 562.595 ;
        RECT 6.290 558.400 54.145 558.525 ;
      LAYER Pwell ;
        RECT 6.290 554.880 993.310 558.400 ;
      LAYER Nwell ;
        RECT 6.290 554.755 62.545 554.880 ;
        RECT 6.290 550.685 993.310 554.755 ;
        RECT 6.290 550.560 236.145 550.685 ;
      LAYER Pwell ;
        RECT 6.290 547.040 993.310 550.560 ;
      LAYER Nwell ;
        RECT 6.290 546.915 16.625 547.040 ;
        RECT 6.290 542.845 993.310 546.915 ;
        RECT 6.290 542.720 14.945 542.845 ;
      LAYER Pwell ;
        RECT 6.290 539.200 993.310 542.720 ;
      LAYER Nwell ;
        RECT 6.290 539.075 183.160 539.200 ;
        RECT 6.290 535.005 993.310 539.075 ;
        RECT 6.290 534.880 196.945 535.005 ;
      LAYER Pwell ;
        RECT 6.290 531.360 993.310 534.880 ;
      LAYER Nwell ;
        RECT 6.290 531.235 51.905 531.360 ;
        RECT 6.290 527.165 993.310 531.235 ;
        RECT 6.290 527.040 72.625 527.165 ;
      LAYER Pwell ;
        RECT 6.290 523.520 993.310 527.040 ;
      LAYER Nwell ;
        RECT 6.290 523.395 18.305 523.520 ;
        RECT 6.290 519.325 993.310 523.395 ;
        RECT 6.290 519.200 32.865 519.325 ;
      LAYER Pwell ;
        RECT 6.290 515.680 993.310 519.200 ;
      LAYER Nwell ;
        RECT 6.290 515.555 14.945 515.680 ;
        RECT 6.290 511.485 993.310 515.555 ;
        RECT 6.290 511.360 618.110 511.485 ;
      LAYER Pwell ;
        RECT 6.290 507.840 993.310 511.360 ;
      LAYER Nwell ;
        RECT 6.290 507.715 103.425 507.840 ;
        RECT 6.290 503.645 993.310 507.715 ;
        RECT 6.290 503.520 240.065 503.645 ;
      LAYER Pwell ;
        RECT 6.290 500.000 993.310 503.520 ;
      LAYER Nwell ;
        RECT 6.290 499.875 53.585 500.000 ;
        RECT 6.290 495.805 993.310 499.875 ;
        RECT 6.290 495.680 51.905 495.805 ;
      LAYER Pwell ;
        RECT 6.290 492.160 993.310 495.680 ;
      LAYER Nwell ;
        RECT 6.290 492.035 26.705 492.160 ;
        RECT 6.290 487.965 993.310 492.035 ;
        RECT 6.290 487.840 14.385 487.965 ;
      LAYER Pwell ;
        RECT 6.290 484.320 993.310 487.840 ;
      LAYER Nwell ;
        RECT 6.290 484.195 23.345 484.320 ;
        RECT 6.290 480.125 993.310 484.195 ;
        RECT 6.290 480.000 230.545 480.125 ;
      LAYER Pwell ;
        RECT 6.290 476.480 993.310 480.000 ;
      LAYER Nwell ;
        RECT 6.290 476.355 54.145 476.480 ;
        RECT 6.290 472.285 993.310 476.355 ;
        RECT 6.290 472.160 51.345 472.285 ;
      LAYER Pwell ;
        RECT 6.290 468.640 993.310 472.160 ;
      LAYER Nwell ;
        RECT 6.290 468.515 212.065 468.640 ;
        RECT 6.290 464.445 993.310 468.515 ;
        RECT 6.290 464.320 32.305 464.445 ;
      LAYER Pwell ;
        RECT 6.290 460.800 993.310 464.320 ;
      LAYER Nwell ;
        RECT 6.290 460.675 67.585 460.800 ;
        RECT 6.290 456.605 993.310 460.675 ;
        RECT 6.290 456.480 125.825 456.605 ;
      LAYER Pwell ;
        RECT 6.290 452.960 993.310 456.480 ;
      LAYER Nwell ;
        RECT 6.290 452.835 110.705 452.960 ;
        RECT 6.290 448.765 993.310 452.835 ;
        RECT 6.290 448.640 52.465 448.765 ;
      LAYER Pwell ;
        RECT 6.290 445.120 993.310 448.640 ;
      LAYER Nwell ;
        RECT 6.290 444.995 182.600 445.120 ;
        RECT 6.290 440.925 993.310 444.995 ;
        RECT 6.290 440.800 44.625 440.925 ;
      LAYER Pwell ;
        RECT 6.290 437.280 993.310 440.800 ;
      LAYER Nwell ;
        RECT 6.290 437.155 169.505 437.280 ;
        RECT 6.290 433.085 993.310 437.155 ;
        RECT 6.290 432.960 90.760 433.085 ;
      LAYER Pwell ;
        RECT 6.290 429.440 993.310 432.960 ;
      LAYER Nwell ;
        RECT 6.290 429.315 53.585 429.440 ;
        RECT 6.290 425.245 993.310 429.315 ;
        RECT 6.290 425.120 111.265 425.245 ;
      LAYER Pwell ;
        RECT 6.290 421.600 993.310 425.120 ;
      LAYER Nwell ;
        RECT 6.290 421.475 141.505 421.600 ;
        RECT 6.290 417.405 993.310 421.475 ;
        RECT 6.290 417.280 132.545 417.405 ;
      LAYER Pwell ;
        RECT 6.290 413.760 993.310 417.280 ;
      LAYER Nwell ;
        RECT 6.290 413.635 70.385 413.760 ;
        RECT 6.290 409.565 993.310 413.635 ;
        RECT 6.290 409.440 82.145 409.565 ;
      LAYER Pwell ;
        RECT 6.290 405.920 993.310 409.440 ;
      LAYER Nwell ;
        RECT 6.290 405.795 101.185 405.920 ;
        RECT 6.290 401.725 993.310 405.795 ;
        RECT 6.290 401.600 78.785 401.725 ;
      LAYER Pwell ;
        RECT 6.290 398.080 993.310 401.600 ;
      LAYER Nwell ;
        RECT 6.290 397.955 174.760 398.080 ;
        RECT 6.290 393.885 993.310 397.955 ;
        RECT 6.290 393.760 93.345 393.885 ;
      LAYER Pwell ;
        RECT 6.290 390.240 993.310 393.760 ;
      LAYER Nwell ;
        RECT 6.290 390.115 141.505 390.240 ;
        RECT 6.290 386.045 993.310 390.115 ;
        RECT 6.290 385.920 93.345 386.045 ;
      LAYER Pwell ;
        RECT 6.290 382.400 993.310 385.920 ;
      LAYER Nwell ;
        RECT 6.290 382.275 140.385 382.400 ;
        RECT 6.290 378.205 993.310 382.275 ;
        RECT 6.290 378.080 198.625 378.205 ;
      LAYER Pwell ;
        RECT 6.290 374.560 993.310 378.080 ;
      LAYER Nwell ;
        RECT 6.290 374.435 169.505 374.560 ;
        RECT 6.290 370.365 993.310 374.435 ;
        RECT 6.290 370.240 164.465 370.365 ;
      LAYER Pwell ;
        RECT 6.290 366.720 993.310 370.240 ;
      LAYER Nwell ;
        RECT 6.290 366.595 106.225 366.720 ;
        RECT 6.290 362.525 993.310 366.595 ;
        RECT 6.290 362.400 79.905 362.525 ;
      LAYER Pwell ;
        RECT 6.290 358.880 993.310 362.400 ;
      LAYER Nwell ;
        RECT 6.290 358.755 105.105 358.880 ;
        RECT 6.290 354.685 993.310 358.755 ;
        RECT 6.290 354.560 81.025 354.685 ;
      LAYER Pwell ;
        RECT 6.290 351.040 993.310 354.560 ;
      LAYER Nwell ;
        RECT 6.290 350.915 152.145 351.040 ;
        RECT 6.290 346.845 993.310 350.915 ;
        RECT 6.290 346.720 165.800 346.845 ;
      LAYER Pwell ;
        RECT 6.290 343.200 993.310 346.720 ;
      LAYER Nwell ;
        RECT 6.290 343.075 264.705 343.200 ;
        RECT 6.290 339.005 993.310 343.075 ;
        RECT 6.290 338.880 93.345 339.005 ;
      LAYER Pwell ;
        RECT 6.290 335.360 993.310 338.880 ;
      LAYER Nwell ;
        RECT 6.290 335.235 91.105 335.360 ;
        RECT 6.290 331.165 993.310 335.235 ;
        RECT 6.290 331.040 217.285 331.165 ;
      LAYER Pwell ;
        RECT 6.290 327.520 993.310 331.040 ;
      LAYER Nwell ;
        RECT 6.290 327.395 73.745 327.520 ;
        RECT 6.290 323.325 993.310 327.395 ;
        RECT 6.290 323.200 117.985 323.325 ;
      LAYER Pwell ;
        RECT 6.290 319.680 993.310 323.200 ;
      LAYER Nwell ;
        RECT 6.290 319.555 79.000 319.680 ;
        RECT 6.290 315.485 993.310 319.555 ;
        RECT 6.290 315.360 157.185 315.485 ;
      LAYER Pwell ;
        RECT 6.290 311.840 993.310 315.360 ;
      LAYER Nwell ;
        RECT 6.290 311.715 315.285 311.840 ;
        RECT 6.290 307.645 993.310 311.715 ;
        RECT 6.290 307.520 121.345 307.645 ;
      LAYER Pwell ;
        RECT 6.290 304.000 993.310 307.520 ;
      LAYER Nwell ;
        RECT 6.290 303.875 106.225 304.000 ;
        RECT 6.290 299.805 993.310 303.875 ;
        RECT 6.290 299.680 86.625 299.805 ;
      LAYER Pwell ;
        RECT 6.290 296.160 993.310 299.680 ;
      LAYER Nwell ;
        RECT 6.290 296.035 218.935 296.160 ;
        RECT 6.290 291.965 993.310 296.035 ;
        RECT 6.290 291.840 784.710 291.965 ;
      LAYER Pwell ;
        RECT 6.290 288.320 993.310 291.840 ;
      LAYER Nwell ;
        RECT 6.290 288.195 73.745 288.320 ;
        RECT 6.290 284.125 993.310 288.195 ;
        RECT 6.290 284.000 150.645 284.125 ;
      LAYER Pwell ;
        RECT 6.290 280.480 993.310 284.000 ;
      LAYER Nwell ;
        RECT 6.290 280.355 73.745 280.480 ;
        RECT 6.290 276.285 993.310 280.355 ;
        RECT 6.290 276.160 202.165 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 993.310 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 72.065 272.640 ;
        RECT 6.290 268.445 993.310 272.515 ;
        RECT 6.290 268.320 202.725 268.445 ;
      LAYER Pwell ;
        RECT 6.290 264.800 993.310 268.320 ;
      LAYER Nwell ;
        RECT 6.290 264.675 340.305 264.800 ;
        RECT 6.290 260.605 993.310 264.675 ;
        RECT 6.290 260.480 194.360 260.605 ;
      LAYER Pwell ;
        RECT 6.290 256.960 993.310 260.480 ;
      LAYER Nwell ;
        RECT 6.290 256.835 65.345 256.960 ;
        RECT 6.290 252.765 993.310 256.835 ;
        RECT 6.290 252.640 200.485 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 993.310 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 217.665 249.120 ;
        RECT 6.290 244.925 993.310 248.995 ;
        RECT 6.290 244.800 131.425 244.925 ;
      LAYER Pwell ;
        RECT 6.290 241.280 993.310 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 58.625 241.280 ;
        RECT 6.290 237.085 993.310 241.155 ;
        RECT 6.290 236.960 54.145 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 993.310 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 131.985 233.440 ;
        RECT 6.290 229.245 993.310 233.315 ;
        RECT 6.290 229.120 189.105 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 993.310 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 101.185 225.600 ;
        RECT 6.290 221.405 993.310 225.475 ;
        RECT 6.290 221.280 71.505 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 993.310 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 98.945 217.760 ;
        RECT 6.290 213.565 993.310 217.635 ;
        RECT 6.290 213.440 71.505 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 993.310 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 100.065 209.920 ;
        RECT 6.290 205.725 993.310 209.795 ;
        RECT 6.290 205.600 279.825 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 993.310 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 422.840 202.080 ;
        RECT 6.290 197.885 993.310 201.955 ;
        RECT 6.290 197.760 195.825 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 993.310 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 191.345 194.240 ;
        RECT 6.290 190.045 993.310 194.115 ;
        RECT 6.290 189.920 77.105 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 993.310 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 141.160 186.400 ;
        RECT 6.290 182.205 993.310 186.275 ;
        RECT 6.290 182.080 250.145 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 993.310 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 67.585 178.560 ;
        RECT 6.290 174.365 993.310 178.435 ;
        RECT 6.290 174.240 174.165 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 993.310 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 63.105 170.720 ;
        RECT 6.290 166.525 993.310 170.595 ;
        RECT 6.290 166.400 196.945 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 993.310 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 64.225 162.880 ;
        RECT 6.290 158.685 993.310 162.755 ;
        RECT 6.290 158.560 162.965 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 993.310 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 91.105 155.040 ;
        RECT 6.290 150.845 993.310 154.915 ;
        RECT 6.290 150.720 83.265 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 993.310 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 137.800 147.200 ;
        RECT 6.290 143.005 993.310 147.075 ;
        RECT 6.290 142.880 328.200 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 993.310 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 70.945 139.360 ;
        RECT 6.290 135.165 993.310 139.235 ;
        RECT 6.290 135.040 160.725 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 993.310 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 73.185 131.520 ;
        RECT 6.290 127.325 993.310 131.395 ;
        RECT 6.290 127.200 110.705 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 993.310 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 269.745 123.680 ;
        RECT 6.290 119.485 993.310 123.555 ;
        RECT 6.290 119.360 132.545 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 993.310 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 215.985 115.840 ;
        RECT 6.290 111.645 993.310 115.715 ;
        RECT 6.290 111.520 78.225 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 993.310 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 208.705 108.000 ;
        RECT 6.290 103.805 993.310 107.875 ;
        RECT 6.290 103.680 78.785 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 993.310 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 110.705 100.160 ;
        RECT 6.290 95.965 993.310 100.035 ;
        RECT 6.290 95.840 124.145 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 993.310 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 106.225 92.320 ;
        RECT 6.290 88.125 993.310 92.195 ;
        RECT 6.290 88.000 133.880 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 993.310 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 144.865 84.480 ;
        RECT 6.290 80.285 993.310 84.355 ;
        RECT 6.290 80.160 157.745 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 993.310 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 193.800 76.640 ;
        RECT 6.290 72.445 993.310 76.515 ;
        RECT 6.290 72.320 247.905 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 993.310 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 177.345 68.800 ;
        RECT 6.290 64.605 993.310 68.675 ;
        RECT 6.290 64.480 267.505 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 993.310 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 215.985 60.960 ;
        RECT 6.290 56.765 993.310 60.835 ;
        RECT 6.290 56.640 171.745 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 993.310 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 302.785 53.120 ;
        RECT 6.290 48.925 993.310 52.995 ;
        RECT 6.290 48.800 289.345 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 993.310 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 184.625 45.280 ;
        RECT 6.290 41.085 993.310 45.155 ;
        RECT 6.290 40.960 189.105 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 993.310 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 258.545 37.440 ;
        RECT 6.290 33.245 993.310 37.315 ;
        RECT 6.290 33.120 210.945 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 993.310 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 257.425 29.600 ;
        RECT 6.290 25.405 993.310 29.475 ;
        RECT 6.290 25.280 195.825 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 993.310 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 212.625 21.760 ;
        RECT 6.290 17.565 993.310 21.635 ;
        RECT 6.290 17.440 665.320 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 993.310 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 992.880 984.220 ;
      LAYER Metal2 ;
        RECT 7.980 995.700 28.820 996.660 ;
        RECT 29.980 995.700 37.780 996.660 ;
        RECT 38.940 995.700 46.740 996.660 ;
        RECT 47.900 995.700 55.700 996.660 ;
        RECT 56.860 995.700 64.660 996.660 ;
        RECT 65.820 995.700 73.620 996.660 ;
        RECT 74.780 995.700 82.580 996.660 ;
        RECT 83.740 995.700 91.540 996.660 ;
        RECT 92.700 995.700 100.500 996.660 ;
        RECT 101.660 995.700 109.460 996.660 ;
        RECT 110.620 995.700 118.420 996.660 ;
        RECT 119.580 995.700 127.380 996.660 ;
        RECT 128.540 995.700 136.340 996.660 ;
        RECT 137.500 995.700 145.300 996.660 ;
        RECT 146.460 995.700 154.260 996.660 ;
        RECT 155.420 995.700 163.220 996.660 ;
        RECT 164.380 995.700 172.180 996.660 ;
        RECT 173.340 995.700 181.140 996.660 ;
        RECT 182.300 995.700 190.100 996.660 ;
        RECT 191.260 995.700 199.060 996.660 ;
        RECT 200.220 995.700 208.020 996.660 ;
        RECT 209.180 995.700 216.980 996.660 ;
        RECT 218.140 995.700 225.940 996.660 ;
        RECT 227.100 995.700 234.900 996.660 ;
        RECT 236.060 995.700 243.860 996.660 ;
        RECT 245.020 995.700 252.820 996.660 ;
        RECT 253.980 995.700 261.780 996.660 ;
        RECT 262.940 995.700 270.740 996.660 ;
        RECT 271.900 995.700 279.700 996.660 ;
        RECT 280.860 995.700 288.660 996.660 ;
        RECT 289.820 995.700 297.620 996.660 ;
        RECT 298.780 995.700 306.580 996.660 ;
        RECT 307.740 995.700 315.540 996.660 ;
        RECT 316.700 995.700 324.500 996.660 ;
        RECT 325.660 995.700 333.460 996.660 ;
        RECT 334.620 995.700 342.420 996.660 ;
        RECT 343.580 995.700 351.380 996.660 ;
        RECT 352.540 995.700 360.340 996.660 ;
        RECT 361.500 995.700 369.300 996.660 ;
        RECT 370.460 995.700 378.260 996.660 ;
        RECT 379.420 995.700 387.220 996.660 ;
        RECT 388.380 995.700 396.180 996.660 ;
        RECT 397.340 995.700 405.140 996.660 ;
        RECT 406.300 995.700 414.100 996.660 ;
        RECT 415.260 995.700 423.060 996.660 ;
        RECT 424.220 995.700 432.020 996.660 ;
        RECT 433.180 995.700 440.980 996.660 ;
        RECT 442.140 995.700 449.940 996.660 ;
        RECT 451.100 995.700 458.900 996.660 ;
        RECT 460.060 995.700 467.860 996.660 ;
        RECT 469.020 995.700 476.820 996.660 ;
        RECT 477.980 995.700 485.780 996.660 ;
        RECT 486.940 995.700 494.740 996.660 ;
        RECT 495.900 995.700 503.700 996.660 ;
        RECT 504.860 995.700 512.660 996.660 ;
        RECT 513.820 995.700 521.620 996.660 ;
        RECT 522.780 995.700 530.580 996.660 ;
        RECT 531.740 995.700 539.540 996.660 ;
        RECT 540.700 995.700 548.500 996.660 ;
        RECT 549.660 995.700 557.460 996.660 ;
        RECT 558.620 995.700 566.420 996.660 ;
        RECT 567.580 995.700 575.380 996.660 ;
        RECT 576.540 995.700 584.340 996.660 ;
        RECT 585.500 995.700 593.300 996.660 ;
        RECT 594.460 995.700 602.260 996.660 ;
        RECT 603.420 995.700 611.220 996.660 ;
        RECT 612.380 995.700 620.180 996.660 ;
        RECT 621.340 995.700 629.140 996.660 ;
        RECT 630.300 995.700 638.100 996.660 ;
        RECT 639.260 995.700 647.060 996.660 ;
        RECT 648.220 995.700 656.020 996.660 ;
        RECT 657.180 995.700 664.980 996.660 ;
        RECT 666.140 995.700 673.940 996.660 ;
        RECT 675.100 995.700 682.900 996.660 ;
        RECT 684.060 995.700 691.860 996.660 ;
        RECT 693.020 995.700 700.820 996.660 ;
        RECT 701.980 995.700 709.780 996.660 ;
        RECT 710.940 995.700 718.740 996.660 ;
        RECT 719.900 995.700 727.700 996.660 ;
        RECT 728.860 995.700 736.660 996.660 ;
        RECT 737.820 995.700 745.620 996.660 ;
        RECT 746.780 995.700 754.580 996.660 ;
        RECT 755.740 995.700 763.540 996.660 ;
        RECT 764.700 995.700 772.500 996.660 ;
        RECT 773.660 995.700 781.460 996.660 ;
        RECT 782.620 995.700 790.420 996.660 ;
        RECT 791.580 995.700 799.380 996.660 ;
        RECT 800.540 995.700 808.340 996.660 ;
        RECT 809.500 995.700 817.300 996.660 ;
        RECT 818.460 995.700 826.260 996.660 ;
        RECT 827.420 995.700 835.220 996.660 ;
        RECT 836.380 995.700 844.180 996.660 ;
        RECT 845.340 995.700 853.140 996.660 ;
        RECT 854.300 995.700 862.100 996.660 ;
        RECT 863.260 995.700 871.060 996.660 ;
        RECT 872.220 995.700 880.020 996.660 ;
        RECT 881.180 995.700 888.980 996.660 ;
        RECT 890.140 995.700 897.940 996.660 ;
        RECT 899.100 995.700 906.900 996.660 ;
        RECT 908.060 995.700 915.860 996.660 ;
        RECT 917.020 995.700 924.820 996.660 ;
        RECT 925.980 995.700 933.780 996.660 ;
        RECT 934.940 995.700 942.740 996.660 ;
        RECT 943.900 995.700 951.700 996.660 ;
        RECT 952.860 995.700 960.660 996.660 ;
        RECT 961.820 995.700 969.620 996.660 ;
        RECT 970.780 995.700 992.180 996.660 ;
        RECT 7.980 4.300 992.180 995.700 ;
        RECT 7.980 2.330 15.380 4.300 ;
        RECT 16.540 2.330 25.460 4.300 ;
        RECT 26.620 2.330 35.540 4.300 ;
        RECT 36.700 2.330 45.620 4.300 ;
        RECT 46.780 2.330 55.700 4.300 ;
        RECT 56.860 2.330 65.780 4.300 ;
        RECT 66.940 2.330 75.860 4.300 ;
        RECT 77.020 2.330 85.940 4.300 ;
        RECT 87.100 2.330 96.020 4.300 ;
        RECT 97.180 2.330 106.100 4.300 ;
        RECT 107.260 2.330 116.180 4.300 ;
        RECT 117.340 2.330 126.260 4.300 ;
        RECT 127.420 2.330 136.340 4.300 ;
        RECT 137.500 2.330 146.420 4.300 ;
        RECT 147.580 2.330 156.500 4.300 ;
        RECT 157.660 2.330 166.580 4.300 ;
        RECT 167.740 2.330 176.660 4.300 ;
        RECT 177.820 2.330 186.740 4.300 ;
        RECT 187.900 2.330 196.820 4.300 ;
        RECT 197.980 2.330 206.900 4.300 ;
        RECT 208.060 2.330 216.980 4.300 ;
        RECT 218.140 2.330 227.060 4.300 ;
        RECT 228.220 2.330 237.140 4.300 ;
        RECT 238.300 2.330 247.220 4.300 ;
        RECT 248.380 2.330 257.300 4.300 ;
        RECT 258.460 2.330 267.380 4.300 ;
        RECT 268.540 2.330 277.460 4.300 ;
        RECT 278.620 2.330 287.540 4.300 ;
        RECT 288.700 2.330 297.620 4.300 ;
        RECT 298.780 2.330 307.700 4.300 ;
        RECT 308.860 2.330 317.780 4.300 ;
        RECT 318.940 2.330 327.860 4.300 ;
        RECT 329.020 2.330 337.940 4.300 ;
        RECT 339.100 2.330 348.020 4.300 ;
        RECT 349.180 2.330 358.100 4.300 ;
        RECT 359.260 2.330 368.180 4.300 ;
        RECT 369.340 2.330 378.260 4.300 ;
        RECT 379.420 2.330 388.340 4.300 ;
        RECT 389.500 2.330 398.420 4.300 ;
        RECT 399.580 2.330 408.500 4.300 ;
        RECT 409.660 2.330 418.580 4.300 ;
        RECT 419.740 2.330 428.660 4.300 ;
        RECT 429.820 2.330 438.740 4.300 ;
        RECT 439.900 2.330 448.820 4.300 ;
        RECT 449.980 2.330 458.900 4.300 ;
        RECT 460.060 2.330 468.980 4.300 ;
        RECT 470.140 2.330 479.060 4.300 ;
        RECT 480.220 2.330 489.140 4.300 ;
        RECT 490.300 2.330 499.220 4.300 ;
        RECT 500.380 2.330 509.300 4.300 ;
        RECT 510.460 2.330 519.380 4.300 ;
        RECT 520.540 2.330 529.460 4.300 ;
        RECT 530.620 2.330 539.540 4.300 ;
        RECT 540.700 2.330 549.620 4.300 ;
        RECT 550.780 2.330 559.700 4.300 ;
        RECT 560.860 2.330 569.780 4.300 ;
        RECT 570.940 2.330 579.860 4.300 ;
        RECT 581.020 2.330 589.940 4.300 ;
        RECT 591.100 2.330 600.020 4.300 ;
        RECT 601.180 2.330 610.100 4.300 ;
        RECT 611.260 2.330 620.180 4.300 ;
        RECT 621.340 2.330 630.260 4.300 ;
        RECT 631.420 2.330 640.340 4.300 ;
        RECT 641.500 2.330 650.420 4.300 ;
        RECT 651.580 2.330 660.500 4.300 ;
        RECT 661.660 2.330 670.580 4.300 ;
        RECT 671.740 2.330 680.660 4.300 ;
        RECT 681.820 2.330 690.740 4.300 ;
        RECT 691.900 2.330 700.820 4.300 ;
        RECT 701.980 2.330 710.900 4.300 ;
        RECT 712.060 2.330 720.980 4.300 ;
        RECT 722.140 2.330 731.060 4.300 ;
        RECT 732.220 2.330 741.140 4.300 ;
        RECT 742.300 2.330 751.220 4.300 ;
        RECT 752.380 2.330 761.300 4.300 ;
        RECT 762.460 2.330 771.380 4.300 ;
        RECT 772.540 2.330 781.460 4.300 ;
        RECT 782.620 2.330 791.540 4.300 ;
        RECT 792.700 2.330 801.620 4.300 ;
        RECT 802.780 2.330 811.700 4.300 ;
        RECT 812.860 2.330 821.780 4.300 ;
        RECT 822.940 2.330 831.860 4.300 ;
        RECT 833.020 2.330 841.940 4.300 ;
        RECT 843.100 2.330 852.020 4.300 ;
        RECT 853.180 2.330 862.100 4.300 ;
        RECT 863.260 2.330 872.180 4.300 ;
        RECT 873.340 2.330 882.260 4.300 ;
        RECT 883.420 2.330 892.340 4.300 ;
        RECT 893.500 2.330 902.420 4.300 ;
        RECT 903.580 2.330 912.500 4.300 ;
        RECT 913.660 2.330 922.580 4.300 ;
        RECT 923.740 2.330 932.660 4.300 ;
        RECT 933.820 2.330 942.740 4.300 ;
        RECT 943.900 2.330 952.820 4.300 ;
        RECT 953.980 2.330 962.900 4.300 ;
        RECT 964.060 2.330 972.980 4.300 ;
        RECT 974.140 2.330 983.060 4.300 ;
        RECT 984.220 2.330 992.180 4.300 ;
      LAYER Metal3 ;
        RECT 7.930 2.380 992.230 994.980 ;
      LAYER Metal4 ;
        RECT 74.620 15.080 98.740 981.030 ;
        RECT 100.940 15.080 175.540 981.030 ;
        RECT 177.740 15.080 252.340 981.030 ;
        RECT 254.540 15.080 329.140 981.030 ;
        RECT 331.340 15.080 405.940 981.030 ;
        RECT 408.140 15.080 482.740 981.030 ;
        RECT 484.940 15.080 559.540 981.030 ;
        RECT 561.740 15.080 636.340 981.030 ;
        RECT 638.540 15.080 713.140 981.030 ;
        RECT 715.340 15.080 789.940 981.030 ;
        RECT 792.140 15.080 866.740 981.030 ;
        RECT 868.940 15.080 943.540 981.030 ;
        RECT 945.740 15.080 955.220 981.030 ;
        RECT 74.620 2.890 955.220 15.080 ;
  END
END tinyrv
END LIBRARY

